magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -307 -6982 307 6982
<< psubdiff >>
rect -271 6912 -175 6946
rect 175 6912 271 6946
rect -271 6850 -237 6912
rect 237 6850 271 6912
rect -271 -6912 -237 -6850
rect 237 -6912 271 -6850
rect -271 -6946 -175 -6912
rect 175 -6946 271 -6912
<< psubdiffcont >>
rect -175 6912 175 6946
rect -271 -6850 -237 6850
rect 237 -6850 271 6850
rect -175 -6946 175 -6912
<< xpolycontact >>
rect -141 6384 141 6816
rect -141 -6816 141 -6384
<< ppolyres >>
rect -141 -6384 141 6384
<< locali >>
rect -271 6912 -175 6946
rect 175 6912 271 6946
rect -271 6850 -237 6912
rect 237 6850 271 6912
rect -271 -6912 -237 -6850
rect 237 -6912 271 -6850
rect -271 -6946 -175 -6912
rect 175 -6946 271 -6912
<< viali >>
rect -125 6401 125 6798
rect -125 -6798 125 -6401
<< metal1 >>
rect -131 6798 131 6810
rect -131 6401 -125 6798
rect 125 6401 131 6798
rect -131 6389 131 6401
rect -131 -6401 131 -6389
rect -131 -6798 -125 -6401
rect 125 -6798 131 -6401
rect -131 -6810 131 -6798
<< labels >>
rlabel psubdiffcont 0 -6929 0 -6929 0 B
port 1 nsew
rlabel xpolycontact 0 6781 0 6781 0 R1
port 2 nsew
rlabel xpolycontact 0 -6781 0 -6781 0 R2
port 3 nsew
<< properties >>
string FIXED_BBOX -254 -6929 254 6929
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 64.0 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 319.8 val 14.792k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1 mult 1
<< end >>
