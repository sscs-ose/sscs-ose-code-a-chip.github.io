# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  11.35000 BY  4.900000 ;
  PIN DRAIN
    ANTENNADIFFAREA  4.214000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.575000 11.420000 3.855000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  15.049999 ;
    PORT
      LAYER met1 ;
        RECT 1.905000 0.000000 9.585000 0.685000 ;
        RECT 1.905000 4.215000 9.585000 4.900000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  5.056800 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.045000 11.420000 2.325000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  3.010000 ;
    ANTENNAGATEAREA  1.505000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.045000 0.500000 3.855000 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.990000 1.045000 11.285000 3.855000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT  0.205000 0.925000  1.150000 3.975000 ;
      RECT  0.950000 0.485000  1.280000 0.815000 ;
      RECT  0.950000 0.815000  1.150000 0.925000 ;
      RECT  0.950000 3.975000  1.150000 4.085000 ;
      RECT  0.950000 4.085000  1.280000 4.415000 ;
      RECT  1.760000 0.925000  1.930000 3.975000 ;
      RECT  1.925000 0.000000  9.565000 0.685000 ;
      RECT  1.925000 4.215000  9.565000 4.900000 ;
      RECT  2.540000 0.925000  2.710000 3.975000 ;
      RECT  3.320000 0.925000  3.490000 3.975000 ;
      RECT  4.100000 0.925000  4.270000 3.975000 ;
      RECT  4.880000 0.925000  5.050000 3.975000 ;
      RECT  5.660000 0.925000  5.830000 3.975000 ;
      RECT  6.440000 0.925000  6.610000 3.975000 ;
      RECT  7.220000 0.925000  7.390000 3.975000 ;
      RECT  8.000000 0.925000  8.170000 3.975000 ;
      RECT  8.780000 0.925000  8.950000 3.975000 ;
      RECT  9.560000 0.925000  9.730000 3.975000 ;
      RECT 10.210000 0.485000 10.540000 0.815000 ;
      RECT 10.210000 4.085000 10.540000 4.415000 ;
      RECT 10.340000 0.815000 10.540000 0.925000 ;
      RECT 10.340000 0.925000 11.285000 3.975000 ;
      RECT 10.340000 3.975000 10.540000 4.085000 ;
    LAYER mcon ;
      RECT  0.300000 1.105000  0.470000 1.275000 ;
      RECT  0.300000 1.465000  0.470000 1.635000 ;
      RECT  0.300000 1.825000  0.470000 1.995000 ;
      RECT  0.300000 2.185000  0.470000 2.355000 ;
      RECT  0.300000 2.545000  0.470000 2.715000 ;
      RECT  0.300000 2.905000  0.470000 3.075000 ;
      RECT  0.300000 3.265000  0.470000 3.435000 ;
      RECT  0.300000 3.625000  0.470000 3.795000 ;
      RECT  1.760000 1.105000  1.930000 1.275000 ;
      RECT  1.760000 1.465000  1.930000 1.635000 ;
      RECT  1.760000 1.825000  1.930000 1.995000 ;
      RECT  1.760000 2.185000  1.930000 2.355000 ;
      RECT  1.760000 2.545000  1.930000 2.715000 ;
      RECT  1.760000 2.905000  1.930000 3.075000 ;
      RECT  1.760000 3.265000  1.930000 3.435000 ;
      RECT  1.760000 3.625000  1.930000 3.795000 ;
      RECT  2.060000 0.095000  9.430000 0.625000 ;
      RECT  2.060000 4.275000  9.430000 4.805000 ;
      RECT  2.540000 1.105000  2.710000 1.275000 ;
      RECT  2.540000 1.465000  2.710000 1.635000 ;
      RECT  2.540000 1.825000  2.710000 1.995000 ;
      RECT  2.540000 2.185000  2.710000 2.355000 ;
      RECT  2.540000 2.545000  2.710000 2.715000 ;
      RECT  2.540000 2.905000  2.710000 3.075000 ;
      RECT  2.540000 3.265000  2.710000 3.435000 ;
      RECT  2.540000 3.625000  2.710000 3.795000 ;
      RECT  3.320000 1.105000  3.490000 1.275000 ;
      RECT  3.320000 1.465000  3.490000 1.635000 ;
      RECT  3.320000 1.825000  3.490000 1.995000 ;
      RECT  3.320000 2.185000  3.490000 2.355000 ;
      RECT  3.320000 2.545000  3.490000 2.715000 ;
      RECT  3.320000 2.905000  3.490000 3.075000 ;
      RECT  3.320000 3.265000  3.490000 3.435000 ;
      RECT  3.320000 3.625000  3.490000 3.795000 ;
      RECT  4.100000 1.105000  4.270000 1.275000 ;
      RECT  4.100000 1.465000  4.270000 1.635000 ;
      RECT  4.100000 1.825000  4.270000 1.995000 ;
      RECT  4.100000 2.185000  4.270000 2.355000 ;
      RECT  4.100000 2.545000  4.270000 2.715000 ;
      RECT  4.100000 2.905000  4.270000 3.075000 ;
      RECT  4.100000 3.265000  4.270000 3.435000 ;
      RECT  4.100000 3.625000  4.270000 3.795000 ;
      RECT  4.880000 1.105000  5.050000 1.275000 ;
      RECT  4.880000 1.465000  5.050000 1.635000 ;
      RECT  4.880000 1.825000  5.050000 1.995000 ;
      RECT  4.880000 2.185000  5.050000 2.355000 ;
      RECT  4.880000 2.545000  5.050000 2.715000 ;
      RECT  4.880000 2.905000  5.050000 3.075000 ;
      RECT  4.880000 3.265000  5.050000 3.435000 ;
      RECT  4.880000 3.625000  5.050000 3.795000 ;
      RECT  5.660000 1.105000  5.830000 1.275000 ;
      RECT  5.660000 1.465000  5.830000 1.635000 ;
      RECT  5.660000 1.825000  5.830000 1.995000 ;
      RECT  5.660000 2.185000  5.830000 2.355000 ;
      RECT  5.660000 2.545000  5.830000 2.715000 ;
      RECT  5.660000 2.905000  5.830000 3.075000 ;
      RECT  5.660000 3.265000  5.830000 3.435000 ;
      RECT  5.660000 3.625000  5.830000 3.795000 ;
      RECT  6.440000 1.105000  6.610000 1.275000 ;
      RECT  6.440000 1.465000  6.610000 1.635000 ;
      RECT  6.440000 1.825000  6.610000 1.995000 ;
      RECT  6.440000 2.185000  6.610000 2.355000 ;
      RECT  6.440000 2.545000  6.610000 2.715000 ;
      RECT  6.440000 2.905000  6.610000 3.075000 ;
      RECT  6.440000 3.265000  6.610000 3.435000 ;
      RECT  6.440000 3.625000  6.610000 3.795000 ;
      RECT  7.220000 1.105000  7.390000 1.275000 ;
      RECT  7.220000 1.465000  7.390000 1.635000 ;
      RECT  7.220000 1.825000  7.390000 1.995000 ;
      RECT  7.220000 2.185000  7.390000 2.355000 ;
      RECT  7.220000 2.545000  7.390000 2.715000 ;
      RECT  7.220000 2.905000  7.390000 3.075000 ;
      RECT  7.220000 3.265000  7.390000 3.435000 ;
      RECT  7.220000 3.625000  7.390000 3.795000 ;
      RECT  8.000000 1.105000  8.170000 1.275000 ;
      RECT  8.000000 1.465000  8.170000 1.635000 ;
      RECT  8.000000 1.825000  8.170000 1.995000 ;
      RECT  8.000000 2.185000  8.170000 2.355000 ;
      RECT  8.000000 2.545000  8.170000 2.715000 ;
      RECT  8.000000 2.905000  8.170000 3.075000 ;
      RECT  8.000000 3.265000  8.170000 3.435000 ;
      RECT  8.000000 3.625000  8.170000 3.795000 ;
      RECT  8.780000 1.105000  8.950000 1.275000 ;
      RECT  8.780000 1.465000  8.950000 1.635000 ;
      RECT  8.780000 1.825000  8.950000 1.995000 ;
      RECT  8.780000 2.185000  8.950000 2.355000 ;
      RECT  8.780000 2.545000  8.950000 2.715000 ;
      RECT  8.780000 2.905000  8.950000 3.075000 ;
      RECT  8.780000 3.265000  8.950000 3.435000 ;
      RECT  8.780000 3.625000  8.950000 3.795000 ;
      RECT  9.560000 1.105000  9.730000 1.275000 ;
      RECT  9.560000 1.465000  9.730000 1.635000 ;
      RECT  9.560000 1.825000  9.730000 1.995000 ;
      RECT  9.560000 2.185000  9.730000 2.355000 ;
      RECT  9.560000 2.545000  9.730000 2.715000 ;
      RECT  9.560000 2.905000  9.730000 3.075000 ;
      RECT  9.560000 3.265000  9.730000 3.435000 ;
      RECT  9.560000 3.625000  9.730000 3.795000 ;
      RECT 11.020000 1.105000 11.190000 1.275000 ;
      RECT 11.020000 1.465000 11.190000 1.635000 ;
      RECT 11.020000 1.825000 11.190000 1.995000 ;
      RECT 11.020000 2.185000 11.190000 2.355000 ;
      RECT 11.020000 2.545000 11.190000 2.715000 ;
      RECT 11.020000 2.905000 11.190000 3.075000 ;
      RECT 11.020000 3.265000 11.190000 3.435000 ;
      RECT 11.020000 3.625000 11.190000 3.795000 ;
    LAYER met1 ;
      RECT 1.715000 1.045000 1.975000 3.855000 ;
      RECT 2.495000 1.045000 2.755000 3.855000 ;
      RECT 3.275000 1.045000 3.535000 3.855000 ;
      RECT 4.055000 1.045000 4.315000 3.855000 ;
      RECT 4.835000 1.045000 5.095000 3.855000 ;
      RECT 5.615000 1.045000 5.875000 3.855000 ;
      RECT 6.395000 1.045000 6.655000 3.855000 ;
      RECT 7.175000 1.045000 7.435000 3.855000 ;
      RECT 7.955000 1.045000 8.215000 3.855000 ;
      RECT 8.735000 1.045000 8.995000 3.855000 ;
      RECT 9.515000 1.045000 9.775000 3.855000 ;
    LAYER via ;
      RECT 1.715000 1.075000 1.975000 1.335000 ;
      RECT 1.715000 1.395000 1.975000 1.655000 ;
      RECT 1.715000 1.715000 1.975000 1.975000 ;
      RECT 1.715000 2.035000 1.975000 2.295000 ;
      RECT 2.495000 2.605000 2.755000 2.865000 ;
      RECT 2.495000 2.925000 2.755000 3.185000 ;
      RECT 2.495000 3.245000 2.755000 3.505000 ;
      RECT 2.495000 3.565000 2.755000 3.825000 ;
      RECT 3.275000 1.075000 3.535000 1.335000 ;
      RECT 3.275000 1.395000 3.535000 1.655000 ;
      RECT 3.275000 1.715000 3.535000 1.975000 ;
      RECT 3.275000 2.035000 3.535000 2.295000 ;
      RECT 4.055000 2.605000 4.315000 2.865000 ;
      RECT 4.055000 2.925000 4.315000 3.185000 ;
      RECT 4.055000 3.245000 4.315000 3.505000 ;
      RECT 4.055000 3.565000 4.315000 3.825000 ;
      RECT 4.835000 1.075000 5.095000 1.335000 ;
      RECT 4.835000 1.395000 5.095000 1.655000 ;
      RECT 4.835000 1.715000 5.095000 1.975000 ;
      RECT 4.835000 2.035000 5.095000 2.295000 ;
      RECT 5.615000 2.605000 5.875000 2.865000 ;
      RECT 5.615000 2.925000 5.875000 3.185000 ;
      RECT 5.615000 3.245000 5.875000 3.505000 ;
      RECT 5.615000 3.565000 5.875000 3.825000 ;
      RECT 6.395000 1.075000 6.655000 1.335000 ;
      RECT 6.395000 1.395000 6.655000 1.655000 ;
      RECT 6.395000 1.715000 6.655000 1.975000 ;
      RECT 6.395000 2.035000 6.655000 2.295000 ;
      RECT 7.175000 2.605000 7.435000 2.865000 ;
      RECT 7.175000 2.925000 7.435000 3.185000 ;
      RECT 7.175000 3.245000 7.435000 3.505000 ;
      RECT 7.175000 3.565000 7.435000 3.825000 ;
      RECT 7.955000 1.075000 8.215000 1.335000 ;
      RECT 7.955000 1.395000 8.215000 1.655000 ;
      RECT 7.955000 1.715000 8.215000 1.975000 ;
      RECT 7.955000 2.035000 8.215000 2.295000 ;
      RECT 8.735000 2.605000 8.995000 2.865000 ;
      RECT 8.735000 2.925000 8.995000 3.185000 ;
      RECT 8.735000 3.245000 8.995000 3.505000 ;
      RECT 8.735000 3.565000 8.995000 3.825000 ;
      RECT 9.515000 1.075000 9.775000 1.335000 ;
      RECT 9.515000 1.395000 9.775000 1.655000 ;
      RECT 9.515000 1.715000 9.775000 1.975000 ;
      RECT 9.515000 2.035000 9.775000 2.295000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50
END LIBRARY
