# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF02W1p65L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF02W1p65L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  1.140000 BY  2.760000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.462000 ;
    PORT
      LAYER met2 ;
        RECT 0.620000 1.120000 0.880000 1.760000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.495000 ;
    PORT
      LAYER met1 ;
        RECT 0.425000 2.005000 1.075000 2.295000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 1.295000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  1.785000 ;
        RECT 1.065000 -0.145000 1.295000  1.785000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.390000 1.865000 0.440000 1.945000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.255000 0.405000 1.785000 ;
      RECT 0.415000 1.985000 1.085000 2.315000 ;
      RECT 0.665000 0.255000 0.835000 1.785000 ;
      RECT 1.095000 0.255000 1.265000 1.785000 ;
    LAYER mcon ;
      RECT 0.235000 0.395000 0.405000 0.565000 ;
      RECT 0.235000 0.755000 0.405000 0.925000 ;
      RECT 0.235000 1.115000 0.405000 1.285000 ;
      RECT 0.235000 1.475000 0.405000 1.645000 ;
      RECT 0.485000 2.065000 0.655000 2.235000 ;
      RECT 0.665000 0.395000 0.835000 0.565000 ;
      RECT 0.665000 0.755000 0.835000 0.925000 ;
      RECT 0.665000 1.115000 0.835000 1.285000 ;
      RECT 0.665000 1.475000 0.835000 1.645000 ;
      RECT 0.845000 2.065000 1.015000 2.235000 ;
      RECT 1.095000 0.395000 1.265000 0.565000 ;
      RECT 1.095000 0.755000 1.265000 0.925000 ;
      RECT 1.095000 1.115000 1.265000 1.285000 ;
      RECT 1.095000 1.475000 1.265000 1.645000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 1.785000 ;
    LAYER via ;
      RECT 0.620000 1.150000 0.880000 1.410000 ;
      RECT 0.620000 1.470000 0.880000 1.730000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF02W1p65L0p15
END LIBRARY
