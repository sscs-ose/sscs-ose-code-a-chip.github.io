.param w1_2=30.15
.param w3_4=4.82
.param w5_6=181.25
.param w7_8=29.00
.param w9_10=60.3
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=65u
.param iref_post_layout=65u
