* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+ sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult = 0.94
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult = 1.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult = 0.7
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult = 0.93222
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult = 0.94436
+ sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff = 1.7325e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff = -3.2175e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff = 1.7325e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0 = -0.0038637
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0 = 0.0001511
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0 = -39322.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0 = 0.051917
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0 = 0.055075
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0 = 2.5385e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0 = -3.7667e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0 = 0.10067
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0 = 6.9005e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0 = -0.295
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1 = 7.0812e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1 = -0.29348
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1 = -0.0040259
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1 = 0.00027138
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1 = -36371.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1 = 0.060494
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1 = 2.9833e-13
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1 = 0.076479
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1 = -3.4315e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1 = 0.10562
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2 = 0.090588
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2 = 7.4877e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2 = -0.28595
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2 = -0.0035475
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2 = -2.9036e-5
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2 = 0.061555
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2 = 6.8019e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2 = -35489.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2 = 0.073805
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2 = -3.2017e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3 = 0.10485
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3 = 7.0535e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3 = -0.29455
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3 = -0.0039581
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3 = 0.00037927
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3 = 0.055516
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3 = 7.5609e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3 = -41289.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3 = 0.074445
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3 = -3.2769e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4 = 0.095773
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4 = 7.1146e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4 = -0.29519
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4 = -0.0035685
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4 = -9.8839e-5
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4 = 0.052857
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4 = -3.5551e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4 = -32637.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4 = 0.07767
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4 = -3.8565e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5 = 0.095491
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5 = 7.2833e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5 = -0.29455
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5 = -0.0042313
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5 = 0.00026379
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5 = 0.0542
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5 = 3.0966e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5 = -31131.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5 = 0.07709
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5 = -2.4624e-19
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6 = -3.0234e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6 = 0.10418
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6 = 7.1978e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6 = -0.295
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6 = -0.0038572
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6 = 7.053e-5
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6 = 0.055107
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6 = 2.686e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6 = -32971.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6 = 0.14893
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7 = -3.572e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7 = 0.14303
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7 = 7.5709e-9
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7 = -0.295
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7 = -0.0040301
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7 = 0.00017124
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7 = 0.05296
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7 = -8.4538e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7 = -29165.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7 = 0.35112
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7 = 0.0
.include "sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"
