* SKY130 Spice File.
.param sky130_fd_bs_flash__special_sonosfet_original__tox_slope=5e-3
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_slope=0.026
