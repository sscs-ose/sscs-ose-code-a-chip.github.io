* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.model sky130_fd_pr__diode_pd2nw_05v5_lvt d
+ level = 3.0
+ tlevc = 1.0
+ area = 1.0e+12
* Junction Capacitance Parameters
+ cj = '0.00076823*1e-12*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult' $ Units: farad/meter^2
+ mj = 0.3362
+ pb = 0.6587 $ Units: volt
+ cjsw = '9.152e-011*1e-6*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult' $ Units: farad/meter
+ mjsw = 0.2659
+ php = 0.7418 $ Units: volt
+ cta = 0.0012407 $ Units: 1/coulomb
+ ctp = 0.00037357 $ Units: 1/coulomb
+ tpb = 0.001671 $ Units: volt/coulomb
+ tphp = 0.001246 $ Units: volt/coulomb
* Diode IV Parameters
+ js = 2.1483e-017 $ Units: amper/meter^2
+ jsw = 1.447e-16 $ Units: amper/meter
+ n = 1.3632
+ rs = 600 $ Units: ohm (ohm/meter^2 if area defined)
+ ik = '4.76e-008/1e-12' $ Units: amper/meter^2
+ ikr = '0/1e-12' $ Units: amper/meter^2
+ vb = 12.69 $ Units: volt
+ ibv = 0.00106 $ Units: amper
+ trs = 0 $ Units: 1/coulomb
+ eg = 1.05 $ Units: electron-volt
+ xti = 5.2
+ tref = 30 $ Units: coulomb
* Default Parameters
+ tcv = 0 $ Units: 1/coulomb
+ gap1 = 0.000473 $ Units: electron-volt/coulomb
+ gap2 = 1110.0
+ ttt1 = 0 $ Units: 1/coulomb
+ ttt2 = 0 $ Units: 1/coulomb^2
+ tm1 = 0 $ Units: 1/coulomb
+ tm2 = 0 $ Units: 1/coulomb^2
+ lm = 0 $ Units: meter
+ lp = 0 $ Units: meter
+ wm = 0 $ Units: meter
+ wp = 0 $ Units: meter
+ xm = 0 $ Units: meter
+ xoi = 10000.0
+ xom = 10000 $ Units: angstrom
+ xp = 0 $ Units: meter
+ xw = 0 $ Units: meter
