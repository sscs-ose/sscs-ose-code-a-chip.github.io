MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 38.83 BY 21.59 ;
  PIN IREF
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.03 13.7 8.31 18.22 ;
    END
  END IREF
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.46 6.56 8.74 12.76 ;
      LAYER M2 ;
        RECT 29.5 8.26 36.72 8.54 ;
      LAYER M3 ;
        RECT 8.46 7.375 8.74 7.745 ;
      LAYER M2 ;
        RECT 8.6 7.42 27.09 7.7 ;
      LAYER M1 ;
        RECT 26.965 7.56 27.215 8.4 ;
      LAYER M2 ;
        RECT 27.09 8.26 29.67 8.54 ;
    END
  END OUT
  OBS 
  LAYER M3 ;
        RECT 8.03 6.14 8.31 12.34 ;
  LAYER M2 ;
        RECT 6.28 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 23.91 6.16 31.13 6.44 ;
  LAYER M3 ;
        RECT 8.03 12.18 8.31 12.6 ;
  LAYER M4 ;
        RECT 7.74 12.2 8.17 13 ;
  LAYER M3 ;
        RECT 7.6 12.6 7.88 14.28 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 8.03 5.88 8.31 6.3 ;
  LAYER M2 ;
        RECT 8.17 5.74 17.2 6.02 ;
  LAYER M1 ;
        RECT 17.075 5.88 17.325 6.3 ;
  LAYER M2 ;
        RECT 17.2 6.16 24.08 6.44 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M3 ;
        RECT 7.6 12.415 7.88 12.785 ;
  LAYER M4 ;
        RECT 7.575 12.2 7.905 13 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M3 ;
        RECT 7.6 12.415 7.88 12.785 ;
  LAYER M4 ;
        RECT 7.575 12.2 7.905 13 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M1 ;
        RECT 17.075 5.795 17.325 5.965 ;
  LAYER M2 ;
        RECT 17.03 5.74 17.37 6.02 ;
  LAYER M1 ;
        RECT 17.075 6.215 17.325 6.385 ;
  LAYER M2 ;
        RECT 17.03 6.16 17.37 6.44 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M2 ;
        RECT 8.01 5.74 8.33 6.02 ;
  LAYER M3 ;
        RECT 8.03 5.72 8.31 6.04 ;
  LAYER M3 ;
        RECT 7.6 12.415 7.88 12.785 ;
  LAYER M4 ;
        RECT 7.575 12.2 7.905 13 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M1 ;
        RECT 17.075 5.795 17.325 5.965 ;
  LAYER M2 ;
        RECT 17.03 5.74 17.37 6.02 ;
  LAYER M1 ;
        RECT 17.075 6.215 17.325 6.385 ;
  LAYER M2 ;
        RECT 17.03 6.16 17.37 6.44 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M2 ;
        RECT 8.01 5.74 8.33 6.02 ;
  LAYER M3 ;
        RECT 8.03 5.72 8.31 6.04 ;
  LAYER M3 ;
        RECT 7.6 12.415 7.88 12.785 ;
  LAYER M4 ;
        RECT 7.575 12.2 7.905 13 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M2 ;
        RECT 24.34 7 30.7 7.28 ;
  LAYER M3 ;
        RECT 32.11 7.82 32.39 12.34 ;
  LAYER M2 ;
        RECT 30.53 7 32.25 7.28 ;
  LAYER M3 ;
        RECT 32.11 7.14 32.39 7.98 ;
  LAYER M2 ;
        RECT 32.09 7 32.41 7.28 ;
  LAYER M3 ;
        RECT 32.11 6.98 32.39 7.3 ;
  LAYER M2 ;
        RECT 32.09 7 32.41 7.28 ;
  LAYER M3 ;
        RECT 32.11 6.98 32.39 7.3 ;
  LAYER M2 ;
        RECT 25.2 6.58 29.84 6.86 ;
  LAYER M3 ;
        RECT 22.65 7.82 22.93 12.34 ;
  LAYER M2 ;
        RECT 23.65 6.58 25.37 6.86 ;
  LAYER M3 ;
        RECT 23.51 6.72 23.79 7.14 ;
  LAYER M2 ;
        RECT 22.79 7 23.65 7.28 ;
  LAYER M3 ;
        RECT 22.65 7.14 22.93 7.98 ;
  LAYER M2 ;
        RECT 22.63 7 22.95 7.28 ;
  LAYER M3 ;
        RECT 22.65 6.98 22.93 7.3 ;
  LAYER M2 ;
        RECT 23.49 6.58 23.81 6.86 ;
  LAYER M3 ;
        RECT 23.51 6.56 23.79 6.88 ;
  LAYER M2 ;
        RECT 23.49 7 23.81 7.28 ;
  LAYER M3 ;
        RECT 23.51 6.98 23.79 7.3 ;
  LAYER M2 ;
        RECT 22.63 7 22.95 7.28 ;
  LAYER M3 ;
        RECT 22.65 6.98 22.93 7.3 ;
  LAYER M2 ;
        RECT 23.49 6.58 23.81 6.86 ;
  LAYER M3 ;
        RECT 23.51 6.56 23.79 6.88 ;
  LAYER M2 ;
        RECT 23.49 7 23.81 7.28 ;
  LAYER M3 ;
        RECT 23.51 6.98 23.79 7.3 ;
  LAYER M3 ;
        RECT 8.89 2.78 9.17 13.18 ;
  LAYER M2 ;
        RECT 18.32 8.26 25.54 8.54 ;
  LAYER M3 ;
        RECT 8.89 8.215 9.17 8.585 ;
  LAYER M2 ;
        RECT 9.03 8.26 18.49 8.54 ;
  LAYER M2 ;
        RECT 8.87 8.26 9.19 8.54 ;
  LAYER M3 ;
        RECT 8.89 8.24 9.17 8.56 ;
  LAYER M2 ;
        RECT 8.87 8.26 9.19 8.54 ;
  LAYER M3 ;
        RECT 8.89 8.24 9.17 8.56 ;
  LAYER M2 ;
        RECT 24.34 2.8 30.7 3.08 ;
  LAYER M2 ;
        RECT 25.2 2.38 29.84 2.66 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 17.305 ;
  LAYER M1 ;
        RECT 5.465 17.555 5.715 18.565 ;
  LAYER M1 ;
        RECT 5.465 19.655 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.035 13.775 5.285 17.305 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 19.655 6.575 20.665 ;
  LAYER M1 ;
        RECT 6.755 13.775 7.005 17.305 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 17.305 ;
  LAYER M1 ;
        RECT 7.185 17.555 7.435 18.565 ;
  LAYER M1 ;
        RECT 7.185 19.655 7.435 20.665 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 17.305 ;
  LAYER M1 ;
        RECT 8.045 17.555 8.295 18.565 ;
  LAYER M1 ;
        RECT 8.045 19.655 8.295 20.665 ;
  LAYER M1 ;
        RECT 8.475 13.775 8.725 17.305 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 17.305 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 19.655 9.155 20.665 ;
  LAYER M1 ;
        RECT 9.335 13.775 9.585 17.305 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 17.305 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 19.655 10.015 20.665 ;
  LAYER M1 ;
        RECT 10.195 13.775 10.445 17.305 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 17.305 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 19.655 10.875 20.665 ;
  LAYER M1 ;
        RECT 11.055 13.775 11.305 17.305 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 17.305 ;
  LAYER M1 ;
        RECT 11.485 17.555 11.735 18.565 ;
  LAYER M1 ;
        RECT 11.485 19.655 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.915 13.775 12.165 17.305 ;
  LAYER M2 ;
        RECT 5.42 17.92 11.78 18.2 ;
  LAYER M2 ;
        RECT 5.42 13.72 11.78 14 ;
  LAYER M2 ;
        RECT 4.99 14.56 12.21 14.84 ;
  LAYER M2 ;
        RECT 5.42 20.02 11.78 20.3 ;
  LAYER M3 ;
        RECT 8.03 13.7 8.31 18.22 ;
  LAYER M2 ;
        RECT 6.28 14.14 10.92 14.42 ;
  LAYER M3 ;
        RECT 8.89 14.54 9.17 20.32 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 11.425 ;
  LAYER M1 ;
        RECT 28.685 11.675 28.935 12.685 ;
  LAYER M1 ;
        RECT 28.685 13.775 28.935 14.785 ;
  LAYER M1 ;
        RECT 28.255 7.895 28.505 11.425 ;
  LAYER M1 ;
        RECT 29.115 7.895 29.365 11.425 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 11.425 ;
  LAYER M1 ;
        RECT 29.545 11.675 29.795 12.685 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.975 7.895 30.225 11.425 ;
  LAYER M1 ;
        RECT 30.405 7.895 30.655 11.425 ;
  LAYER M1 ;
        RECT 30.405 11.675 30.655 12.685 ;
  LAYER M1 ;
        RECT 30.405 13.775 30.655 14.785 ;
  LAYER M1 ;
        RECT 30.835 7.895 31.085 11.425 ;
  LAYER M1 ;
        RECT 31.265 7.895 31.515 11.425 ;
  LAYER M1 ;
        RECT 31.265 11.675 31.515 12.685 ;
  LAYER M1 ;
        RECT 31.265 13.775 31.515 14.785 ;
  LAYER M1 ;
        RECT 31.695 7.895 31.945 11.425 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 11.425 ;
  LAYER M1 ;
        RECT 32.125 11.675 32.375 12.685 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 14.785 ;
  LAYER M1 ;
        RECT 32.555 7.895 32.805 11.425 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 11.425 ;
  LAYER M1 ;
        RECT 32.985 11.675 33.235 12.685 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 14.785 ;
  LAYER M1 ;
        RECT 33.415 7.895 33.665 11.425 ;
  LAYER M1 ;
        RECT 33.845 7.895 34.095 11.425 ;
  LAYER M1 ;
        RECT 33.845 11.675 34.095 12.685 ;
  LAYER M1 ;
        RECT 33.845 13.775 34.095 14.785 ;
  LAYER M1 ;
        RECT 34.275 7.895 34.525 11.425 ;
  LAYER M1 ;
        RECT 34.705 7.895 34.955 11.425 ;
  LAYER M1 ;
        RECT 34.705 11.675 34.955 12.685 ;
  LAYER M1 ;
        RECT 34.705 13.775 34.955 14.785 ;
  LAYER M1 ;
        RECT 35.135 7.895 35.385 11.425 ;
  LAYER M1 ;
        RECT 35.565 7.895 35.815 11.425 ;
  LAYER M1 ;
        RECT 35.565 11.675 35.815 12.685 ;
  LAYER M1 ;
        RECT 35.565 13.775 35.815 14.785 ;
  LAYER M1 ;
        RECT 35.995 7.895 36.245 11.425 ;
  LAYER M1 ;
        RECT 36.425 7.895 36.675 11.425 ;
  LAYER M1 ;
        RECT 36.425 11.675 36.675 12.685 ;
  LAYER M1 ;
        RECT 36.425 13.775 36.675 14.785 ;
  LAYER M1 ;
        RECT 36.855 7.895 37.105 11.425 ;
  LAYER M2 ;
        RECT 28.64 12.04 36.72 12.32 ;
  LAYER M2 ;
        RECT 28.64 7.84 35.86 8.12 ;
  LAYER M2 ;
        RECT 28.21 8.68 37.15 8.96 ;
  LAYER M2 ;
        RECT 28.64 14.14 36.72 14.42 ;
  LAYER M3 ;
        RECT 32.11 7.82 32.39 12.34 ;
  LAYER M2 ;
        RECT 29.5 8.26 36.72 8.54 ;
  LAYER M3 ;
        RECT 32.97 8.66 33.25 14.44 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 11.425 ;
  LAYER M1 ;
        RECT 26.105 11.675 26.355 12.685 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 11.425 ;
  LAYER M1 ;
        RECT 25.245 11.675 25.495 12.685 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 14.785 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M1 ;
        RECT 24.385 7.895 24.635 11.425 ;
  LAYER M1 ;
        RECT 24.385 11.675 24.635 12.685 ;
  LAYER M1 ;
        RECT 24.385 13.775 24.635 14.785 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 11.425 ;
  LAYER M1 ;
        RECT 23.525 11.675 23.775 12.685 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 14.785 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 22.665 11.675 22.915 12.685 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 14.785 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 14.785 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 11.425 ;
  LAYER M1 ;
        RECT 20.945 11.675 21.195 12.685 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 14.785 ;
  LAYER M1 ;
        RECT 20.515 7.895 20.765 11.425 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M1 ;
        RECT 20.085 11.675 20.335 12.685 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 14.785 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.365 11.675 18.615 12.685 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 14.785 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M2 ;
        RECT 18.32 12.04 26.4 12.32 ;
  LAYER M2 ;
        RECT 19.18 7.84 26.4 8.12 ;
  LAYER M2 ;
        RECT 17.89 8.68 26.83 8.96 ;
  LAYER M2 ;
        RECT 18.32 14.14 26.4 14.42 ;
  LAYER M3 ;
        RECT 22.65 7.82 22.93 12.34 ;
  LAYER M2 ;
        RECT 18.32 8.26 25.54 8.54 ;
  LAYER M3 ;
        RECT 21.79 8.66 22.07 14.44 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 9.575 15.175 13.105 ;
  LAYER M1 ;
        RECT 14.925 8.315 15.175 9.325 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 9.575 12.595 13.105 ;
  LAYER M1 ;
        RECT 12.345 8.315 12.595 9.325 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 9.575 12.165 13.105 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.485 9.575 11.735 13.105 ;
  LAYER M1 ;
        RECT 11.485 8.315 11.735 9.325 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.905 9.575 9.155 13.105 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 9.325 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.045 9.575 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 9.325 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 9.575 7.865 13.105 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.185 9.575 7.435 13.105 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 9.325 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 9.575 7.005 13.105 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 6.325 9.575 6.575 13.105 ;
  LAYER M1 ;
        RECT 6.325 8.315 6.575 9.325 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 9.575 6.145 13.105 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 5.465 9.575 5.715 13.105 ;
  LAYER M1 ;
        RECT 5.465 8.315 5.715 9.325 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.035 9.575 5.285 13.105 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 4.605 9.575 4.855 13.105 ;
  LAYER M1 ;
        RECT 4.605 8.315 4.855 9.325 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 9.575 4.425 13.105 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.745 9.575 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.745 8.315 3.995 9.325 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 9.575 3.565 13.105 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 2.885 9.575 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.885 8.315 3.135 9.325 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 2.455 9.575 2.705 13.105 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.025 9.575 2.275 13.105 ;
  LAYER M1 ;
        RECT 2.025 8.315 2.275 9.325 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 1.595 9.575 1.845 13.105 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 1.165 9.575 1.415 13.105 ;
  LAYER M1 ;
        RECT 1.165 8.315 1.415 9.325 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 9.575 0.985 13.105 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 1.12 8.68 16.08 8.96 ;
  LAYER M2 ;
        RECT 1.98 12.88 16.08 13.16 ;
  LAYER M2 ;
        RECT 1.12 12.46 15.22 12.74 ;
  LAYER M2 ;
        RECT 0.69 12.04 16.51 12.32 ;
  LAYER M2 ;
        RECT 1.12 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 16.08 3.08 ;
  LAYER M2 ;
        RECT 1.98 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 0.69 6.16 16.51 6.44 ;
  LAYER M2 ;
        RECT 1.12 0.7 16.08 0.98 ;
  LAYER M3 ;
        RECT 8.89 2.78 9.17 13.18 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 12.76 ;
  LAYER M3 ;
        RECT 8.03 6.14 8.31 12.34 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M2 ;
        RECT 24.34 0.7 30.7 0.98 ;
  LAYER M2 ;
        RECT 24.34 7 30.7 7.28 ;
  LAYER M2 ;
        RECT 25.2 6.58 29.84 6.86 ;
  LAYER M2 ;
        RECT 24.34 2.8 30.7 3.08 ;
  LAYER M2 ;
        RECT 25.2 2.38 29.84 2.66 ;
  LAYER M2 ;
        RECT 23.91 6.16 31.13 6.44 ;
  END 
END CURRENT_MIRROR_OTA
