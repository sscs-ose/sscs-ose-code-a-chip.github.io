** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/tb_cm_ota_working_v2_extracted_transient.sch
**.subckt tb_cm_ota_working_v2_extracted_transient
V1 avdd_1v8 GND 1.8
C1 out GND 50f m=1
V3 inn GND DC 0.9 AC SIN(0.9 0.1 1Meg)
V4 inp GND 0.9
X1 avdd_1v8 out inp inn iref GND cm_ota
I1 GND iref 24u
**** begin user architecture code

** opencircuitdesign pdks isntsall
.lib /opt/pdk/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.temp 27
.option savecurrents
.save all
.control
	op
	write tb_cm_ota_working_v2_extracted.raw
	tran 0.5ns 10us
	plot v(inn) v(out)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  cm_ota.sym # of pins=6
** sym_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sym
** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sch
.subckt cm_ota VDD VOUT VINP VINN ID VSS

X0 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# VINP m1_2892_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X1 m1_2290_6188# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X2 li_749_5779# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X3 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# VINN li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X4 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# VINN m1_2290_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X5 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# VINP li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X6 li_749_5779# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X7 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# VINN m1_2290_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X8 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# VINP m1_2892_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X9 li_749_5779# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X10 m1_2290_6188# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X11 li_749_5779# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X12 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# VINP li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X13 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# VINP m1_2892_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X14 m1_2892_6188# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X15 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# VINN li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X16 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VINN m1_2290_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X17 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_462# VINN m1_2290_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X18 m1_2892_6188# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X19 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# VINP m1_2892_6188# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X20 li_749_5779# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X21 li_749_5779# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X22 li_749_5779# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X23 li_749_5779# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X24 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# VINN li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X25 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# VINP li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X26 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# VINN li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X27 m1_2290_6188# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X28 m1_2892_6188# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X29 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# VINP li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X30 m1_2892_6188# VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X31 m1_2290_6188# VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X32 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# ID li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X33 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X34 VSS ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X35 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_402_462# ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X36 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_746_462# ID li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X37 VSS ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X38 VSS ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_402_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X39 VSS ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_746_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X40 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_918_462# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X41 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X42 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X43 li_749_5779# ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_918_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X44 ID ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X45 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_230_462# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X46 ID ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_230_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X47 li_749_5779# ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X48 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_1638# m1_2290_6188# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X49 m1_2290_6188# m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_1638# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X50 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_462# m1_2290_6188# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X51 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# m1_2290_6188# m1_2290_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X52 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_462# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X53 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_462# VDD sky130_fd_pr__pfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X54 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_3990# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X55 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X56 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# VDD sky130_fd_pr__pfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X57 VOUT m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X58 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_3990# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X59 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# m1_2290_6188# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X60 m1_2290_6188# m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_3990# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X61 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_2814# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X62 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_3990# m1_2290_6188# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X63 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X64 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# VDD sky130_fd_pr__pfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X65 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_462# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X66 m1_2290_6188# m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X67 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_2814# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X68 VOUT m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_2814# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X69 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X70 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_5166# m1_2290_6188# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X71 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_2814# m1_2290_6188# m1_2290_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X72 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X73 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X74 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X75 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_5166# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X76 m1_2290_6188# m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X77 m1_2290_6188# m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X78 VOUT m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_462# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X79 VOUT m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X80 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_5166# m1_2290_6188# m1_2290_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X81 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# m1_2290_6188# m1_2290_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X82 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_1638# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X83 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X84 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_1638# m1_2290_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X85 VDD m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# VDD sky130_fd_pr__pfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X86 VOUT m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X87 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_462# m1_2290_6188# m1_2290_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X88 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_1638# m1_2892_6188# m2_918_3743# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=1.47 ps=13.3 w=1.05 l=0.15
X89 m1_2892_6188# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_1638# VDD sky130_fd_pr__pfet_01v8 ad=1.47 pd=13.3 as=0.294 ps=2.66 w=1.05 l=0.15
X90 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_462# m1_2892_6188# m2_918_3743# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X91 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_3990# m1_2892_6188# m1_2892_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X92 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_462# VDD sky130_fd_pr__pfet_01v8 ad=8.51 pd=79.2 as=0.294 ps=2.66 w=1.05 l=0.15
X93 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_462# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X94 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_3990# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.294 ps=2.66 w=1.05 l=0.15
X95 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X96 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_3990# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X97 m2_918_3743# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X98 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_3990# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X99 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_2814# m1_2892_6188# m2_918_3743# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X100 m1_2892_6188# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_3990# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X101 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_2814# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.294 ps=2.66 w=1.05 l=0.15
X102 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_3990# m1_2892_6188# m2_918_3743# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X103 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X104 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_2814# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X105 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_462# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X106 m1_2892_6188# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X107 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_2814# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X108 m2_918_3743# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_2814# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X109 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_5166# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.294 ps=2.66 w=1.05 l=0.15
X110 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_5166# m1_2892_6188# m2_918_3743# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X111 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_2814# m1_2892_6188# m1_2892_6188# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X112 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X113 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_5166# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X114 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X115 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_5166# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X116 m1_2892_6188# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X117 m1_2892_6188# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X118 m2_918_3743# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_462# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X119 m2_918_3743# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_5166# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X120 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_5166# m1_2892_6188# m1_2892_6188# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X121 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_1638# m1_2892_6188# m1_2892_6188# VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X122 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_1638# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X123 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.66 as=0 ps=0 w=1.05 l=0.15
X124 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_1638# m1_2892_6188# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X125 VDD m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_1638# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X126 m2_918_3743# m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X127 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_462# m1_2892_6188# m1_2892_6188# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.05 l=0.15
X128 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_1638# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X129 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X130 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X131 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X132 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X133 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X134 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X135 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X136 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X137 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X138 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X139 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X140 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X141 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_1638# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X142 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X143 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X144 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X145 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X146 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_462# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X147 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X148 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X149 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X150 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X151 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X152 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X153 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_3990# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X154 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X155 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X156 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_462# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X157 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X158 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X159 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X160 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X161 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X162 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X163 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X164 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X165 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X166 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X167 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X168 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_2814# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X169 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X170 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X171 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X172 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X173 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X174 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X175 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X176 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X177 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X178 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X179 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X180 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X181 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_2814# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X182 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X183 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X184 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# m2_918_3743# m2_918_3743# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X185 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_2814# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X186 li_749_5779# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# VSS sky130_fd_pr__nfet_01v8 ad=0.278 pd=2.63 as=0.147 ps=1.33 w=1.05 l=0.15
X187 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X188 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# m2_918_3743# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X189 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# m2_918_3743# li_749_5779# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.278 ps=2.63 w=1.05 l=0.15
X190 m2_918_3743# m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
X191 VOUT m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# VSS sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.33 as=0.147 ps=1.33 w=1.05 l=0.15
C0 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# 0.00223f
C1 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_5166# m2_918_3743# 0.00819f
C2 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_918_462# ID 0.00249f
C3 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# m1_2892_6188# 0.00819f
C4 VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# 0.00249f
C5 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# m1_2290_6188# 0.00819f
C6 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# VOUT 0.00819f
C7 li_749_5779# SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# 3.9e-19
C8 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# VDD 9.53e-19
C9 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_1638# 0.0149f
C10 li_749_5779# VINN 0.934f
C11 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_5166# VDD 0.0172f
C12 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# 0.0111f
C13 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# 0.0139f
C14 li_749_5779# VINP 0.825f
C15 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_5166# m1_2290_6188# 0.00249f
C16 VDD SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# 0.00303f
C17 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_402_462# VDD 0.00316f
C18 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_230_462# VDD 0.00324f
C19 VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# 0.0019f
C20 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_5166# 0.0172f
C21 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# VINP 0.0025f
C22 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# m2_918_3743# 5.75e-19
C23 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# 0.0111f
C24 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# m1_2892_6188# 0.00107f
C25 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# m1_2290_6188# 0.011f
C26 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_1638# m2_918_3743# 0.0168f
C27 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# 0.00819f
C28 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# m2_918_3743# 0.0107f
C29 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# 0.00208f
C30 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# VOUT 0.00819f
C31 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# VDD 0.0166f
C32 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# VOUT 0.00819f
C33 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# VINP 0.00249f
C34 VOUT VINP 5.35e-19
C35 ID m1_2892_6188# 1.78e-19
C36 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# li_749_5779# 0.0111f
C37 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# VDD 0.00292f
C38 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# m2_918_3743# 0.00819f
C39 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# VDD 0.00211f
C40 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_1638# m1_2290_6188# 0.0107f
C41 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# 0.00231f
C42 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# m2_918_3743# 0.00249f
C43 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# VOUT 0.00819f
C44 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_1638# m1_2290_6188# 0.00861f
C45 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_1638# VDD 0.0172f
C46 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_1638# VDD 0.0111f
C47 m1_2290_6188# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# 0.00139f
C48 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# m1_2290_6188# 0.011f
C49 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# 0.00175f
C50 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# 0.0111f
C51 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# 0.0117f
C52 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# 0.0128f
C53 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# 0.00208f
C54 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# m2_918_3743# 0.0135f
C55 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# 0.012f
C56 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# VDD 0.00173f
C57 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# 0.0111f
C58 VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# 0.00405f
C59 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# 0.0111f
C60 VDD SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# 0.00245f
C61 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_462# m1_2290_6188# 0.0143f
C62 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# 0.0139f
C63 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_3990# VDD 0.0147f
C64 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_402_462# ID 0.0128f
C65 ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# 0.00532f
C66 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_230_462# ID 0.00971f
C67 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# m2_918_3743# 0.00464f
C68 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# 0.00338f
C69 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# VDD 0.00141f
C70 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# m1_2290_6188# 0.011f
C71 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_1638# m1_2892_6188# 0.00819f
C72 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# m1_2290_6188# 0.00819f
C73 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_5166# m1_2892_6188# 0.00249f
C74 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# 0.0117f
C75 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# VDD 0.00182f
C76 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VDD 9.53e-19
C77 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# 0.0111f
C78 VDD SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# 0.00264f
C79 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# VOUT 0.00819f
C80 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# VINP 0.00127f
C81 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# 0.0111f
C82 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# m2_918_3743# 0.00152f
C83 li_749_5779# VOUT 6.71f
C84 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# m2_918_3743# 0.00249f
C85 m2_918_3743# VINP 5.35e-19
C86 m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# 0.00374f
C87 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# m1_2892_6188# 0.00819f
C88 VINN m1_2290_6188# 0.561f
C89 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_2814# 0.00819f
C90 VDD SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# 0.00254f
C91 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_3990# 0.00819f
C92 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# 0.0116f
C93 VDD VINN 0.11f
C94 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_3990# m2_918_3743# 0.00819f
C95 VINP m1_2290_6188# 0.443f
C96 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# m1_2892_6188# 0.01f
C97 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# 0.00203f
C98 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# m2_918_3743# 0.00401f
C99 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# 0.00155f
C100 VDD VINP 0.21f
C101 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# ID 0.00819f
C102 li_749_5779# SCM_NMOS_5643887_X2_Y1_1725189358_0/a_746_462# 0.0087f
C103 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_3990# VDD 0.0111f
C104 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# 0.0111f
C105 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# VDD 0.00167f
C106 m2_918_3743# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_1638# 0.00819f
C107 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# m2_918_3743# 0.0135f
C108 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# VINP 0.00552f
C109 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# m1_2892_6188# 0.00107f
C110 m1_2892_6188# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# 0.00819f
C111 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# m1_2290_6188# 0.00107f
C112 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# 0.0111f
C113 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_3990# m1_2892_6188# 0.00819f
C114 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# 0.0122f
C115 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# ID 0.00249f
C116 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_1638# 0.0111f
C117 m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# 0.011f
C118 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# VDD 0.00173f
C119 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# 0.0138f
C120 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_2814# m2_918_3743# 0.00819f
C121 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# 0.00819f
C122 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# 0.00819f
C123 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_462# 0.0192f
C124 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# m1_2892_6188# 0.00107f
C125 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# 0.0149f
C126 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_462# 0.0111f
C127 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# 0.00249f
C128 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# 0.0111f
C129 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# VINP 0.00249f
C130 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# m1_2290_6188# 0.00107f
C131 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# 9.53e-19
C132 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# ID 0.0107f
C133 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_2814# VDD 0.0153f
C134 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# 0.00203f
C135 m1_2290_6188# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# 0.00819f
C136 VINN ID 3.92e-19
C137 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# VDD 0.0138f
C138 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_462# li_749_5779# 0.0111f
C139 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# 0.00128f
C140 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# 0.00208f
C141 li_749_5779# m2_918_3743# 6.04f
C142 ID VINP 0.0139f
C143 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# 0.00311f
C144 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_5166# m1_2290_6188# 0.0168f
C145 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_5166# m2_918_3743# 0.00819f
C146 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# 0.0111f
C147 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_2814# VDD 0.0111f
C148 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_5166# 0.0111f
C149 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_5166# 0.0111f
C150 li_749_5779# m1_2290_6188# 2.65f
C151 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# 0.0152f
C152 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_1638# 0.0172f
C153 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_462# 0.00819f
C154 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_2814# m1_2290_6188# 0.0168f
C155 m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# 0.00107f
C156 m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_2814# 0.00249f
C157 li_749_5779# VDD 1.23f
C158 VINN m1_2892_6188# 0.202f
C159 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_2814# 0.0111f
C160 m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_3990# 0.00861f
C161 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_2814# 0.0172f
C162 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_5166# 0.0142f
C163 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_2814# 0.0172f
C164 VINP m1_2892_6188# 0.585f
C165 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_3990# 0.0111f
C166 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# li_749_5779# 0.0132f
C167 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_462# VOUT 0.00819f
C168 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# 9.53e-19
C169 m2_918_3743# VOUT 5.46f
C170 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_3990# m1_2892_6188# 0.00861f
C171 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# 0.0111f
C172 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# li_749_5779# 0.0132f
C173 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_5166# 0.00819f
C174 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# VOUT 0.00819f
C175 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# VOUT 0.00146f
C176 VOUT m1_2290_6188# 4.05f
C177 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_3990# 0.0111f
C178 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# VINN 0.00152f
C179 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# VDD 0.00208f
C180 VDD VOUT 6.28f
C181 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_462# 0.00819f
C182 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_462# m1_2290_6188# 0.0168f
C183 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# m1_2290_6188# 0.00107f
C184 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# m1_2892_6188# 0.011f
C185 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_2814# VOUT 0.00819f
C186 VOUT SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_462# 0.00819f
C187 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_462# 0.0111f
C188 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_918_462# li_749_5779# 0.00819f
C189 m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_1638# 0.00861f
C190 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# 0.012f
C191 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_2814# 0.0111f
C192 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# 0.00107f
C193 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# 0.0132f
C194 m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# 0.00107f
C195 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# m2_918_3743# 0.00819f
C196 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_3990# m1_2290_6188# 0.0107f
C197 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# 0.0158f
C198 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_462# m1_2892_6188# 0.0168f
C199 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_3990# 0.0172f
C200 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# 0.00175f
C201 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# 0.0111f
C202 VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# 0.0018f
C203 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# m1_2290_6188# 0.00107f
C204 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# m1_2892_6188# 0.00819f
C205 VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# 0.00612f
C206 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# li_749_5779# 0.0111f
C207 m1_2290_6188# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# 0.00819f
C208 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# VDD 0.0116f
C209 li_749_5779# ID 0.844f
C210 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# VINP 0.00249f
C211 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# m1_2892_6188# 0.011f
C212 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# VINP 0.00249f
C213 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# 9.53e-19
C214 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# 0.0117f
C215 m1_2892_6188# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# 0.00303f
C216 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_2814# VOUT 0.00819f
C217 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_3990# 0.0172f
C218 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_462# 0.00249f
C219 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_2814# m1_2892_6188# 0.0168f
C220 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# VOUT 0.00819f
C221 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_402_5166# m1_2892_6188# 0.0168f
C222 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# 0.0111f
C223 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# 0.0111f
C224 li_749_5779# m1_2892_6188# 1.6f
C225 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_1638# 0.0172f
C226 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# 0.0101f
C227 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# m2_918_3743# 0.00947f
C228 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_462# m2_918_3743# 0.00861f
C229 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# m1_2290_6188# 0.00819f
C230 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# 0.0132f
C231 VOUT ID 0.00314f
C232 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# VDD 9.53e-19
C233 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_462# m2_918_3743# 0.00819f
C234 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# m1_2892_6188# 0.00819f
C235 VINP DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# 0.00249f
C236 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# m1_2290_6188# 0.00107f
C237 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# 0.00532f
C238 m2_918_3743# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# 0.00186f
C239 m2_918_3743# m1_2290_6188# 0.253f
C240 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_1638# 0.0107f
C241 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_2814# m2_918_3743# 0.00819f
C242 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# VDD 0.0111f
C243 VDD m2_918_3743# 8.17f
C244 m2_918_3743# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_462# 0.00819f
C245 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_462# VINP 0.00249f
C246 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# li_749_5779# 0.0111f
C247 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_462# 0.0172f
C248 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# m1_2290_6188# 0.00819f
C249 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_5166# 0.0148f
C250 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# 0.00819f
C251 ID SCM_NMOS_5643887_X2_Y1_1725189358_0/a_746_462# 0.00861f
C252 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# m1_2892_6188# 0.0121f
C253 VOUT m1_2892_6188# 0.0214f
C254 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# 0.00329f
C255 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_2814# 0.00249f
C256 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# m2_918_3743# 0.0107f
C257 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# 0.0139f
C258 VDD m1_2290_6188# 13.9f
C259 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# 0.00292f
C260 li_749_5779# SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# 0.00819f
C261 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VINN 0.0019f
C262 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# 0.00819f
C263 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_2814# VDD 0.0172f
C264 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# m1_2892_6188# 0.011f
C265 VDD SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_462# 0.0147f
C266 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# m2_918_3743# 0.00819f
C267 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_462# 0.015f
C268 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_462# m1_2290_6188# 0.00249f
C269 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VINP 0.00181f
C270 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_462# 0.0172f
C271 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# VDD 0.00323f
C272 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_3990# m2_918_3743# 0.0168f
C273 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# m1_2290_6188# 0.00195f
C274 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# VDD 0.00331f
C275 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# VDD 9.53e-19
C276 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# 0.0141f
C277 m2_918_3743# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# 5.75e-19
C278 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_1638# 0.0111f
C279 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# m1_2892_6188# 0.00374f
C280 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_2814# 0.00861f
C281 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# 0.0107f
C282 m1_2290_6188# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# 0.00819f
C283 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# li_749_5779# 0.0117f
C284 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_746_1638# li_749_5779# 0.0111f
C285 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_574_5166# VOUT 0.00819f
C286 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# 0.0139f
C287 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_3990# m1_2892_6188# 0.0107f
C288 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# m2_918_3743# 0.00128f
C289 VDD SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# 0.015f
C290 VINN VINP 2.14f
C291 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# 0.0132f
C292 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# 0.00296f
C293 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# 0.00167f
C294 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# m1_2290_6188# 0.00374f
C295 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# m1_2290_6188# 0.00819f
C296 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# 0.0132f
C297 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# m2_918_3743# 0.0128f
C298 m1_2892_6188# SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_1638# 0.0107f
C299 m2_918_3743# ID 0.339f
C300 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# VDD 0.0111f
C301 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# 0.0153f
C302 VDD DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# 0.00208f
C303 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# li_749_5779# 0.0111f
C304 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# VOUT 0.00819f
C305 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# m2_918_3743# 0.00971f
C306 li_749_5779# SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# 5.02e-19
C307 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# 0.00158f
C308 ID m1_2290_6188# 0.0032f
C309 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# VDD 0.00155f
C310 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_462# li_749_5779# 0.0111f
C311 VDD ID 0.356f
C312 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# 0.0111f
C313 VOUT SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# 0.00819f
C314 li_749_5779# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# 0.0133f
C315 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# m1_2892_6188# 0.00374f
C316 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# 0.00608f
C317 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# m2_918_3743# 0.0107f
C318 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# VDD 0.00359f
C319 m2_918_3743# m1_2892_6188# 4.13f
C320 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_462# m1_2892_6188# 0.00249f
C321 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_402_1638# VOUT 0.00819f
C322 m2_918_3743# SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# 0.00249f
C323 li_749_5779# SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# 0.00136f
C324 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# li_749_5779# 0.0111f
C325 m1_2892_6188# m1_2290_6188# 2.32f
C326 li_749_5779# DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# 0.0111f
C327 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# m1_2892_6188# 0.00819f
C328 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# VOUT 0.00819f
C329 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_574_2814# m1_2892_6188# 0.00249f
C330 li_749_5779# SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# 0.0085f
C331 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# VDD 0.00182f
C332 VDD SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# 0.00137f
C333 VDD m1_2892_6188# 13.9f
C334 VINN DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# 0.00472f
C335 VOUT VSS 1.59f
C336 VDD VSS 47.1f
C337 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_462# VSS 0.00208f
C338 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_462# VSS 0.00208f
C339 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_462# VSS 0.00208f
C340 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_462# VSS 0.00573f
C341 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_462# VSS 0.00531f
C342 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_462# VSS 0.00474f
C343 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_1638# VSS 9.53e-19
C344 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_1638# VSS 9.53e-19
C345 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_1638# VSS 9.53e-19
C346 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_1638# VSS 0.00157f
C347 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_1638# VSS 0.00168f
C348 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_1638# VSS 0.00181f
C349 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_2814# VSS 4.71e-19
C350 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_2814# VSS 4.71e-19
C351 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_2814# VSS 4.71e-19
C352 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_2814# VSS 0.00109f
C353 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_2814# VSS 0.0012f
C354 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_2814# VSS 0.00133f
C355 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1434_3990# VSS 0.00208f
C356 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1262_3990# VSS 0.00208f
C357 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_1090_3990# VSS 0.00208f
C358 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_918_3990# VSS 0.00253f
C359 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_574_3990# VSS 0.0027f
C360 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_402_3990# VSS 0.00281f
C361 SCM_NMOS_B_85279373_X2_Y4_1725189359_0/a_230_3990# VSS 0.00293f
C362 m2_918_3743# VSS 17.5f
C363 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_462# VSS 0.00144f
C364 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_462# VSS 0.003f
C365 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_1638# VSS 0.0011f
C366 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_1638# VSS 0.00214f
C367 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_2814# VSS 8.44e-19
C368 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_2814# VSS 0.00149f
C369 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_3990# VSS 0.00144f
C370 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_3990# VSS 0.003f
C371 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_746_5166# VSS 0.0011f
C372 SCM_PMOS_85912433_X1_Y5_1725189360_1/a_230_5166# VSS 0.00214f
C373 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_462# VSS 0.00384f
C374 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_462# VSS 0.00378f
C375 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_1638# VSS 0.00231f
C376 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_1638# VSS 0.00291f
C377 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_2814# VSS 0.00167f
C378 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_2814# VSS 0.00227f
C379 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_3990# VSS 0.00318f
C380 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_3990# VSS 0.00378f
C381 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_746_5166# VSS 0.00231f
C382 SCM_PMOS_85912433_X1_Y5_1725189360_0/a_230_5166# VSS 0.00291f
C383 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1434_462# VSS 0.0139f
C384 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1262_462# VSS 0.0144f
C385 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_1090_462# VSS 0.015f
C386 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_918_462# VSS 0.018f
C387 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_746_462# VSS 0.0111f
C388 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_574_462# VSS 0.0116f
C389 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_402_462# VSS 0.0116f
C390 SCM_NMOS_5643887_X2_Y1_1725189358_0/a_230_462# VSS 0.0116f
C391 ID VSS 5.85f
C392 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_462# VSS 0.00175f
C393 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_462# VSS 0.00311f
C394 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_462# VSS 0.00212f
C395 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_918_462# VSS 0.00174f
C396 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_462# VSS 0.00151f
C397 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_462# VSS 0.00138f
C398 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_462# VSS 0.00124f
C399 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1434_1638# VSS 0.00232f
C400 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1262_1638# VSS 0.00378f
C401 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_1090_1638# VSS 0.00285f
C402 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_746_1638# VSS 0.0022f
C403 m1_2892_6188# VSS 2.89f
C404 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_574_1638# VSS 0.00208f
C405 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_402_1638# VSS 0.00194f
C406 m1_2290_6188# VSS 3.23f
C407 DP_NMOS_B_6171529_X2_Y2_1725189357_0/a_230_1638# VSS 0.0018f
C408 li_749_5779# VSS 7.76f
C409 VINP VSS 3.7f
C410 VINN VSS 4.01f
.ends

.GLOBAL GND
.end
