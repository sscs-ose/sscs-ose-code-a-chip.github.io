MACRO DCL_NMOS_S_54772057_X4_Y24
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_54772057_X4_Y24 0 0 ;
  SIZE 5160 BY 142800 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 260 2720 140020 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 680 3150 142120 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 142465 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 68545 ;
    LAYER M1 ;
      RECT 2025 68795 2275 69805 ;
    LAYER M1 ;
      RECT 2025 70895 2275 74425 ;
    LAYER M1 ;
      RECT 2025 74675 2275 75685 ;
    LAYER M1 ;
      RECT 2025 76775 2275 80305 ;
    LAYER M1 ;
      RECT 2025 80555 2275 81565 ;
    LAYER M1 ;
      RECT 2025 82655 2275 86185 ;
    LAYER M1 ;
      RECT 2025 86435 2275 87445 ;
    LAYER M1 ;
      RECT 2025 88535 2275 92065 ;
    LAYER M1 ;
      RECT 2025 92315 2275 93325 ;
    LAYER M1 ;
      RECT 2025 94415 2275 97945 ;
    LAYER M1 ;
      RECT 2025 98195 2275 99205 ;
    LAYER M1 ;
      RECT 2025 100295 2275 103825 ;
    LAYER M1 ;
      RECT 2025 104075 2275 105085 ;
    LAYER M1 ;
      RECT 2025 106175 2275 109705 ;
    LAYER M1 ;
      RECT 2025 109955 2275 110965 ;
    LAYER M1 ;
      RECT 2025 112055 2275 115585 ;
    LAYER M1 ;
      RECT 2025 115835 2275 116845 ;
    LAYER M1 ;
      RECT 2025 117935 2275 121465 ;
    LAYER M1 ;
      RECT 2025 121715 2275 122725 ;
    LAYER M1 ;
      RECT 2025 123815 2275 127345 ;
    LAYER M1 ;
      RECT 2025 127595 2275 128605 ;
    LAYER M1 ;
      RECT 2025 129695 2275 133225 ;
    LAYER M1 ;
      RECT 2025 133475 2275 134485 ;
    LAYER M1 ;
      RECT 2025 135575 2275 139105 ;
    LAYER M1 ;
      RECT 2025 139355 2275 140365 ;
    LAYER M1 ;
      RECT 2025 141455 2275 142465 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M1 ;
      RECT 2455 65015 2705 68545 ;
    LAYER M1 ;
      RECT 2455 70895 2705 74425 ;
    LAYER M1 ;
      RECT 2455 76775 2705 80305 ;
    LAYER M1 ;
      RECT 2455 82655 2705 86185 ;
    LAYER M1 ;
      RECT 2455 88535 2705 92065 ;
    LAYER M1 ;
      RECT 2455 94415 2705 97945 ;
    LAYER M1 ;
      RECT 2455 100295 2705 103825 ;
    LAYER M1 ;
      RECT 2455 106175 2705 109705 ;
    LAYER M1 ;
      RECT 2455 112055 2705 115585 ;
    LAYER M1 ;
      RECT 2455 117935 2705 121465 ;
    LAYER M1 ;
      RECT 2455 123815 2705 127345 ;
    LAYER M1 ;
      RECT 2455 129695 2705 133225 ;
    LAYER M1 ;
      RECT 2455 135575 2705 139105 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 39145 ;
    LAYER M1 ;
      RECT 2885 39395 3135 40405 ;
    LAYER M1 ;
      RECT 2885 41495 3135 45025 ;
    LAYER M1 ;
      RECT 2885 45275 3135 46285 ;
    LAYER M1 ;
      RECT 2885 47375 3135 50905 ;
    LAYER M1 ;
      RECT 2885 51155 3135 52165 ;
    LAYER M1 ;
      RECT 2885 53255 3135 56785 ;
    LAYER M1 ;
      RECT 2885 57035 3135 58045 ;
    LAYER M1 ;
      RECT 2885 59135 3135 62665 ;
    LAYER M1 ;
      RECT 2885 62915 3135 63925 ;
    LAYER M1 ;
      RECT 2885 65015 3135 68545 ;
    LAYER M1 ;
      RECT 2885 68795 3135 69805 ;
    LAYER M1 ;
      RECT 2885 70895 3135 74425 ;
    LAYER M1 ;
      RECT 2885 74675 3135 75685 ;
    LAYER M1 ;
      RECT 2885 76775 3135 80305 ;
    LAYER M1 ;
      RECT 2885 80555 3135 81565 ;
    LAYER M1 ;
      RECT 2885 82655 3135 86185 ;
    LAYER M1 ;
      RECT 2885 86435 3135 87445 ;
    LAYER M1 ;
      RECT 2885 88535 3135 92065 ;
    LAYER M1 ;
      RECT 2885 92315 3135 93325 ;
    LAYER M1 ;
      RECT 2885 94415 3135 97945 ;
    LAYER M1 ;
      RECT 2885 98195 3135 99205 ;
    LAYER M1 ;
      RECT 2885 100295 3135 103825 ;
    LAYER M1 ;
      RECT 2885 104075 3135 105085 ;
    LAYER M1 ;
      RECT 2885 106175 3135 109705 ;
    LAYER M1 ;
      RECT 2885 109955 3135 110965 ;
    LAYER M1 ;
      RECT 2885 112055 3135 115585 ;
    LAYER M1 ;
      RECT 2885 115835 3135 116845 ;
    LAYER M1 ;
      RECT 2885 117935 3135 121465 ;
    LAYER M1 ;
      RECT 2885 121715 3135 122725 ;
    LAYER M1 ;
      RECT 2885 123815 3135 127345 ;
    LAYER M1 ;
      RECT 2885 127595 3135 128605 ;
    LAYER M1 ;
      RECT 2885 129695 3135 133225 ;
    LAYER M1 ;
      RECT 2885 133475 3135 134485 ;
    LAYER M1 ;
      RECT 2885 135575 3135 139105 ;
    LAYER M1 ;
      RECT 2885 139355 3135 140365 ;
    LAYER M1 ;
      RECT 2885 141455 3135 142465 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3315 47375 3565 50905 ;
    LAYER M1 ;
      RECT 3315 53255 3565 56785 ;
    LAYER M1 ;
      RECT 3315 59135 3565 62665 ;
    LAYER M1 ;
      RECT 3315 65015 3565 68545 ;
    LAYER M1 ;
      RECT 3315 70895 3565 74425 ;
    LAYER M1 ;
      RECT 3315 76775 3565 80305 ;
    LAYER M1 ;
      RECT 3315 82655 3565 86185 ;
    LAYER M1 ;
      RECT 3315 88535 3565 92065 ;
    LAYER M1 ;
      RECT 3315 94415 3565 97945 ;
    LAYER M1 ;
      RECT 3315 100295 3565 103825 ;
    LAYER M1 ;
      RECT 3315 106175 3565 109705 ;
    LAYER M1 ;
      RECT 3315 112055 3565 115585 ;
    LAYER M1 ;
      RECT 3315 117935 3565 121465 ;
    LAYER M1 ;
      RECT 3315 123815 3565 127345 ;
    LAYER M1 ;
      RECT 3315 129695 3565 133225 ;
    LAYER M1 ;
      RECT 3315 135575 3565 139105 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 33265 ;
    LAYER M1 ;
      RECT 3745 33515 3995 34525 ;
    LAYER M1 ;
      RECT 3745 35615 3995 39145 ;
    LAYER M1 ;
      RECT 3745 39395 3995 40405 ;
    LAYER M1 ;
      RECT 3745 41495 3995 45025 ;
    LAYER M1 ;
      RECT 3745 45275 3995 46285 ;
    LAYER M1 ;
      RECT 3745 47375 3995 50905 ;
    LAYER M1 ;
      RECT 3745 51155 3995 52165 ;
    LAYER M1 ;
      RECT 3745 53255 3995 56785 ;
    LAYER M1 ;
      RECT 3745 57035 3995 58045 ;
    LAYER M1 ;
      RECT 3745 59135 3995 62665 ;
    LAYER M1 ;
      RECT 3745 62915 3995 63925 ;
    LAYER M1 ;
      RECT 3745 65015 3995 68545 ;
    LAYER M1 ;
      RECT 3745 68795 3995 69805 ;
    LAYER M1 ;
      RECT 3745 70895 3995 74425 ;
    LAYER M1 ;
      RECT 3745 74675 3995 75685 ;
    LAYER M1 ;
      RECT 3745 76775 3995 80305 ;
    LAYER M1 ;
      RECT 3745 80555 3995 81565 ;
    LAYER M1 ;
      RECT 3745 82655 3995 86185 ;
    LAYER M1 ;
      RECT 3745 86435 3995 87445 ;
    LAYER M1 ;
      RECT 3745 88535 3995 92065 ;
    LAYER M1 ;
      RECT 3745 92315 3995 93325 ;
    LAYER M1 ;
      RECT 3745 94415 3995 97945 ;
    LAYER M1 ;
      RECT 3745 98195 3995 99205 ;
    LAYER M1 ;
      RECT 3745 100295 3995 103825 ;
    LAYER M1 ;
      RECT 3745 104075 3995 105085 ;
    LAYER M1 ;
      RECT 3745 106175 3995 109705 ;
    LAYER M1 ;
      RECT 3745 109955 3995 110965 ;
    LAYER M1 ;
      RECT 3745 112055 3995 115585 ;
    LAYER M1 ;
      RECT 3745 115835 3995 116845 ;
    LAYER M1 ;
      RECT 3745 117935 3995 121465 ;
    LAYER M1 ;
      RECT 3745 121715 3995 122725 ;
    LAYER M1 ;
      RECT 3745 123815 3995 127345 ;
    LAYER M1 ;
      RECT 3745 127595 3995 128605 ;
    LAYER M1 ;
      RECT 3745 129695 3995 133225 ;
    LAYER M1 ;
      RECT 3745 133475 3995 134485 ;
    LAYER M1 ;
      RECT 3745 135575 3995 139105 ;
    LAYER M1 ;
      RECT 3745 139355 3995 140365 ;
    LAYER M1 ;
      RECT 3745 141455 3995 142465 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4175 35615 4425 39145 ;
    LAYER M1 ;
      RECT 4175 41495 4425 45025 ;
    LAYER M1 ;
      RECT 4175 47375 4425 50905 ;
    LAYER M1 ;
      RECT 4175 53255 4425 56785 ;
    LAYER M1 ;
      RECT 4175 59135 4425 62665 ;
    LAYER M1 ;
      RECT 4175 65015 4425 68545 ;
    LAYER M1 ;
      RECT 4175 70895 4425 74425 ;
    LAYER M1 ;
      RECT 4175 76775 4425 80305 ;
    LAYER M1 ;
      RECT 4175 82655 4425 86185 ;
    LAYER M1 ;
      RECT 4175 88535 4425 92065 ;
    LAYER M1 ;
      RECT 4175 94415 4425 97945 ;
    LAYER M1 ;
      RECT 4175 100295 4425 103825 ;
    LAYER M1 ;
      RECT 4175 106175 4425 109705 ;
    LAYER M1 ;
      RECT 4175 112055 4425 115585 ;
    LAYER M1 ;
      RECT 4175 117935 4425 121465 ;
    LAYER M1 ;
      RECT 4175 123815 4425 127345 ;
    LAYER M1 ;
      RECT 4175 129695 4425 133225 ;
    LAYER M1 ;
      RECT 4175 135575 4425 139105 ;
    LAYER M2 ;
      RECT 1120 280 4040 560 ;
    LAYER M2 ;
      RECT 1120 4480 4040 4760 ;
    LAYER M2 ;
      RECT 690 700 4470 980 ;
    LAYER M2 ;
      RECT 1120 6160 4040 6440 ;
    LAYER M2 ;
      RECT 1120 10360 4040 10640 ;
    LAYER M2 ;
      RECT 690 6580 4470 6860 ;
    LAYER M2 ;
      RECT 1120 12040 4040 12320 ;
    LAYER M2 ;
      RECT 1120 16240 4040 16520 ;
    LAYER M2 ;
      RECT 690 12460 4470 12740 ;
    LAYER M2 ;
      RECT 1120 17920 4040 18200 ;
    LAYER M2 ;
      RECT 1120 22120 4040 22400 ;
    LAYER M2 ;
      RECT 690 18340 4470 18620 ;
    LAYER M2 ;
      RECT 1120 23800 4040 24080 ;
    LAYER M2 ;
      RECT 1120 28000 4040 28280 ;
    LAYER M2 ;
      RECT 690 24220 4470 24500 ;
    LAYER M2 ;
      RECT 1120 29680 4040 29960 ;
    LAYER M2 ;
      RECT 1120 33880 4040 34160 ;
    LAYER M2 ;
      RECT 690 30100 4470 30380 ;
    LAYER M2 ;
      RECT 1120 35560 4040 35840 ;
    LAYER M2 ;
      RECT 1120 39760 4040 40040 ;
    LAYER M2 ;
      RECT 690 35980 4470 36260 ;
    LAYER M2 ;
      RECT 1120 41440 4040 41720 ;
    LAYER M2 ;
      RECT 1120 45640 4040 45920 ;
    LAYER M2 ;
      RECT 690 41860 4470 42140 ;
    LAYER M2 ;
      RECT 1120 47320 4040 47600 ;
    LAYER M2 ;
      RECT 1120 51520 4040 51800 ;
    LAYER M2 ;
      RECT 690 47740 4470 48020 ;
    LAYER M2 ;
      RECT 1120 53200 4040 53480 ;
    LAYER M2 ;
      RECT 1120 57400 4040 57680 ;
    LAYER M2 ;
      RECT 690 53620 4470 53900 ;
    LAYER M2 ;
      RECT 1120 59080 4040 59360 ;
    LAYER M2 ;
      RECT 1120 63280 4040 63560 ;
    LAYER M2 ;
      RECT 690 59500 4470 59780 ;
    LAYER M2 ;
      RECT 1120 64960 4040 65240 ;
    LAYER M2 ;
      RECT 1120 69160 4040 69440 ;
    LAYER M2 ;
      RECT 690 65380 4470 65660 ;
    LAYER M2 ;
      RECT 1120 70840 4040 71120 ;
    LAYER M2 ;
      RECT 1120 75040 4040 75320 ;
    LAYER M2 ;
      RECT 690 71260 4470 71540 ;
    LAYER M2 ;
      RECT 1120 76720 4040 77000 ;
    LAYER M2 ;
      RECT 1120 80920 4040 81200 ;
    LAYER M2 ;
      RECT 690 77140 4470 77420 ;
    LAYER M2 ;
      RECT 1120 82600 4040 82880 ;
    LAYER M2 ;
      RECT 1120 86800 4040 87080 ;
    LAYER M2 ;
      RECT 690 83020 4470 83300 ;
    LAYER M2 ;
      RECT 1120 88480 4040 88760 ;
    LAYER M2 ;
      RECT 1120 92680 4040 92960 ;
    LAYER M2 ;
      RECT 690 88900 4470 89180 ;
    LAYER M2 ;
      RECT 1120 94360 4040 94640 ;
    LAYER M2 ;
      RECT 1120 98560 4040 98840 ;
    LAYER M2 ;
      RECT 690 94780 4470 95060 ;
    LAYER M2 ;
      RECT 1120 100240 4040 100520 ;
    LAYER M2 ;
      RECT 1120 104440 4040 104720 ;
    LAYER M2 ;
      RECT 690 100660 4470 100940 ;
    LAYER M2 ;
      RECT 1120 106120 4040 106400 ;
    LAYER M2 ;
      RECT 1120 110320 4040 110600 ;
    LAYER M2 ;
      RECT 690 106540 4470 106820 ;
    LAYER M2 ;
      RECT 1120 112000 4040 112280 ;
    LAYER M2 ;
      RECT 1120 116200 4040 116480 ;
    LAYER M2 ;
      RECT 690 112420 4470 112700 ;
    LAYER M2 ;
      RECT 1120 117880 4040 118160 ;
    LAYER M2 ;
      RECT 1120 122080 4040 122360 ;
    LAYER M2 ;
      RECT 690 118300 4470 118580 ;
    LAYER M2 ;
      RECT 1120 123760 4040 124040 ;
    LAYER M2 ;
      RECT 1120 127960 4040 128240 ;
    LAYER M2 ;
      RECT 690 124180 4470 124460 ;
    LAYER M2 ;
      RECT 1120 129640 4040 129920 ;
    LAYER M2 ;
      RECT 1120 133840 4040 134120 ;
    LAYER M2 ;
      RECT 690 130060 4470 130340 ;
    LAYER M2 ;
      RECT 1120 135520 4040 135800 ;
    LAYER M2 ;
      RECT 1120 139720 4040 140000 ;
    LAYER M2 ;
      RECT 1120 141820 4040 142100 ;
    LAYER M2 ;
      RECT 690 135940 4470 136220 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 35615 3095 35785 ;
    LAYER V1 ;
      RECT 2925 39815 3095 39985 ;
    LAYER V1 ;
      RECT 2925 41495 3095 41665 ;
    LAYER V1 ;
      RECT 2925 45695 3095 45865 ;
    LAYER V1 ;
      RECT 2925 47375 3095 47545 ;
    LAYER V1 ;
      RECT 2925 51575 3095 51745 ;
    LAYER V1 ;
      RECT 2925 53255 3095 53425 ;
    LAYER V1 ;
      RECT 2925 57455 3095 57625 ;
    LAYER V1 ;
      RECT 2925 59135 3095 59305 ;
    LAYER V1 ;
      RECT 2925 63335 3095 63505 ;
    LAYER V1 ;
      RECT 2925 65015 3095 65185 ;
    LAYER V1 ;
      RECT 2925 69215 3095 69385 ;
    LAYER V1 ;
      RECT 2925 70895 3095 71065 ;
    LAYER V1 ;
      RECT 2925 75095 3095 75265 ;
    LAYER V1 ;
      RECT 2925 76775 3095 76945 ;
    LAYER V1 ;
      RECT 2925 80975 3095 81145 ;
    LAYER V1 ;
      RECT 2925 82655 3095 82825 ;
    LAYER V1 ;
      RECT 2925 86855 3095 87025 ;
    LAYER V1 ;
      RECT 2925 88535 3095 88705 ;
    LAYER V1 ;
      RECT 2925 92735 3095 92905 ;
    LAYER V1 ;
      RECT 2925 94415 3095 94585 ;
    LAYER V1 ;
      RECT 2925 98615 3095 98785 ;
    LAYER V1 ;
      RECT 2925 100295 3095 100465 ;
    LAYER V1 ;
      RECT 2925 104495 3095 104665 ;
    LAYER V1 ;
      RECT 2925 106175 3095 106345 ;
    LAYER V1 ;
      RECT 2925 110375 3095 110545 ;
    LAYER V1 ;
      RECT 2925 112055 3095 112225 ;
    LAYER V1 ;
      RECT 2925 116255 3095 116425 ;
    LAYER V1 ;
      RECT 2925 117935 3095 118105 ;
    LAYER V1 ;
      RECT 2925 122135 3095 122305 ;
    LAYER V1 ;
      RECT 2925 123815 3095 123985 ;
    LAYER V1 ;
      RECT 2925 128015 3095 128185 ;
    LAYER V1 ;
      RECT 2925 129695 3095 129865 ;
    LAYER V1 ;
      RECT 2925 133895 3095 134065 ;
    LAYER V1 ;
      RECT 2925 135575 3095 135745 ;
    LAYER V1 ;
      RECT 2925 139775 3095 139945 ;
    LAYER V1 ;
      RECT 2925 141875 3095 142045 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 29735 3955 29905 ;
    LAYER V1 ;
      RECT 3785 33935 3955 34105 ;
    LAYER V1 ;
      RECT 3785 35615 3955 35785 ;
    LAYER V1 ;
      RECT 3785 39815 3955 39985 ;
    LAYER V1 ;
      RECT 3785 41495 3955 41665 ;
    LAYER V1 ;
      RECT 3785 45695 3955 45865 ;
    LAYER V1 ;
      RECT 3785 47375 3955 47545 ;
    LAYER V1 ;
      RECT 3785 51575 3955 51745 ;
    LAYER V1 ;
      RECT 3785 53255 3955 53425 ;
    LAYER V1 ;
      RECT 3785 57455 3955 57625 ;
    LAYER V1 ;
      RECT 3785 59135 3955 59305 ;
    LAYER V1 ;
      RECT 3785 63335 3955 63505 ;
    LAYER V1 ;
      RECT 3785 65015 3955 65185 ;
    LAYER V1 ;
      RECT 3785 69215 3955 69385 ;
    LAYER V1 ;
      RECT 3785 70895 3955 71065 ;
    LAYER V1 ;
      RECT 3785 75095 3955 75265 ;
    LAYER V1 ;
      RECT 3785 76775 3955 76945 ;
    LAYER V1 ;
      RECT 3785 80975 3955 81145 ;
    LAYER V1 ;
      RECT 3785 82655 3955 82825 ;
    LAYER V1 ;
      RECT 3785 86855 3955 87025 ;
    LAYER V1 ;
      RECT 3785 88535 3955 88705 ;
    LAYER V1 ;
      RECT 3785 92735 3955 92905 ;
    LAYER V1 ;
      RECT 3785 94415 3955 94585 ;
    LAYER V1 ;
      RECT 3785 98615 3955 98785 ;
    LAYER V1 ;
      RECT 3785 100295 3955 100465 ;
    LAYER V1 ;
      RECT 3785 104495 3955 104665 ;
    LAYER V1 ;
      RECT 3785 106175 3955 106345 ;
    LAYER V1 ;
      RECT 3785 110375 3955 110545 ;
    LAYER V1 ;
      RECT 3785 112055 3955 112225 ;
    LAYER V1 ;
      RECT 3785 116255 3955 116425 ;
    LAYER V1 ;
      RECT 3785 117935 3955 118105 ;
    LAYER V1 ;
      RECT 3785 122135 3955 122305 ;
    LAYER V1 ;
      RECT 3785 123815 3955 123985 ;
    LAYER V1 ;
      RECT 3785 128015 3955 128185 ;
    LAYER V1 ;
      RECT 3785 129695 3955 129865 ;
    LAYER V1 ;
      RECT 3785 133895 3955 134065 ;
    LAYER V1 ;
      RECT 3785 135575 3955 135745 ;
    LAYER V1 ;
      RECT 3785 139775 3955 139945 ;
    LAYER V1 ;
      RECT 3785 141875 3955 142045 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141875 1375 142045 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59135 2235 59305 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65015 2235 65185 ;
    LAYER V1 ;
      RECT 2065 69215 2235 69385 ;
    LAYER V1 ;
      RECT 2065 70895 2235 71065 ;
    LAYER V1 ;
      RECT 2065 75095 2235 75265 ;
    LAYER V1 ;
      RECT 2065 76775 2235 76945 ;
    LAYER V1 ;
      RECT 2065 80975 2235 81145 ;
    LAYER V1 ;
      RECT 2065 82655 2235 82825 ;
    LAYER V1 ;
      RECT 2065 86855 2235 87025 ;
    LAYER V1 ;
      RECT 2065 88535 2235 88705 ;
    LAYER V1 ;
      RECT 2065 92735 2235 92905 ;
    LAYER V1 ;
      RECT 2065 94415 2235 94585 ;
    LAYER V1 ;
      RECT 2065 98615 2235 98785 ;
    LAYER V1 ;
      RECT 2065 100295 2235 100465 ;
    LAYER V1 ;
      RECT 2065 104495 2235 104665 ;
    LAYER V1 ;
      RECT 2065 106175 2235 106345 ;
    LAYER V1 ;
      RECT 2065 110375 2235 110545 ;
    LAYER V1 ;
      RECT 2065 112055 2235 112225 ;
    LAYER V1 ;
      RECT 2065 116255 2235 116425 ;
    LAYER V1 ;
      RECT 2065 117935 2235 118105 ;
    LAYER V1 ;
      RECT 2065 122135 2235 122305 ;
    LAYER V1 ;
      RECT 2065 123815 2235 123985 ;
    LAYER V1 ;
      RECT 2065 128015 2235 128185 ;
    LAYER V1 ;
      RECT 2065 129695 2235 129865 ;
    LAYER V1 ;
      RECT 2065 133895 2235 134065 ;
    LAYER V1 ;
      RECT 2065 135575 2235 135745 ;
    LAYER V1 ;
      RECT 2065 139775 2235 139945 ;
    LAYER V1 ;
      RECT 2065 141875 2235 142045 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 2495 59555 2665 59725 ;
    LAYER V1 ;
      RECT 2495 65435 2665 65605 ;
    LAYER V1 ;
      RECT 2495 71315 2665 71485 ;
    LAYER V1 ;
      RECT 2495 77195 2665 77365 ;
    LAYER V1 ;
      RECT 2495 83075 2665 83245 ;
    LAYER V1 ;
      RECT 2495 88955 2665 89125 ;
    LAYER V1 ;
      RECT 2495 94835 2665 95005 ;
    LAYER V1 ;
      RECT 2495 100715 2665 100885 ;
    LAYER V1 ;
      RECT 2495 106595 2665 106765 ;
    LAYER V1 ;
      RECT 2495 112475 2665 112645 ;
    LAYER V1 ;
      RECT 2495 118355 2665 118525 ;
    LAYER V1 ;
      RECT 2495 124235 2665 124405 ;
    LAYER V1 ;
      RECT 2495 130115 2665 130285 ;
    LAYER V1 ;
      RECT 2495 135995 2665 136165 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 41915 3525 42085 ;
    LAYER V1 ;
      RECT 3355 47795 3525 47965 ;
    LAYER V1 ;
      RECT 3355 53675 3525 53845 ;
    LAYER V1 ;
      RECT 3355 59555 3525 59725 ;
    LAYER V1 ;
      RECT 3355 65435 3525 65605 ;
    LAYER V1 ;
      RECT 3355 71315 3525 71485 ;
    LAYER V1 ;
      RECT 3355 77195 3525 77365 ;
    LAYER V1 ;
      RECT 3355 83075 3525 83245 ;
    LAYER V1 ;
      RECT 3355 88955 3525 89125 ;
    LAYER V1 ;
      RECT 3355 94835 3525 95005 ;
    LAYER V1 ;
      RECT 3355 100715 3525 100885 ;
    LAYER V1 ;
      RECT 3355 106595 3525 106765 ;
    LAYER V1 ;
      RECT 3355 112475 3525 112645 ;
    LAYER V1 ;
      RECT 3355 118355 3525 118525 ;
    LAYER V1 ;
      RECT 3355 124235 3525 124405 ;
    LAYER V1 ;
      RECT 3355 130115 3525 130285 ;
    LAYER V1 ;
      RECT 3355 135995 3525 136165 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 4215 30155 4385 30325 ;
    LAYER V1 ;
      RECT 4215 36035 4385 36205 ;
    LAYER V1 ;
      RECT 4215 41915 4385 42085 ;
    LAYER V1 ;
      RECT 4215 47795 4385 47965 ;
    LAYER V1 ;
      RECT 4215 53675 4385 53845 ;
    LAYER V1 ;
      RECT 4215 59555 4385 59725 ;
    LAYER V1 ;
      RECT 4215 65435 4385 65605 ;
    LAYER V1 ;
      RECT 4215 71315 4385 71485 ;
    LAYER V1 ;
      RECT 4215 77195 4385 77365 ;
    LAYER V1 ;
      RECT 4215 83075 4385 83245 ;
    LAYER V1 ;
      RECT 4215 88955 4385 89125 ;
    LAYER V1 ;
      RECT 4215 94835 4385 95005 ;
    LAYER V1 ;
      RECT 4215 100715 4385 100885 ;
    LAYER V1 ;
      RECT 4215 106595 4385 106765 ;
    LAYER V1 ;
      RECT 4215 112475 4385 112645 ;
    LAYER V1 ;
      RECT 4215 118355 4385 118525 ;
    LAYER V1 ;
      RECT 4215 124235 4385 124405 ;
    LAYER V1 ;
      RECT 4215 130115 4385 130285 ;
    LAYER V1 ;
      RECT 4215 135995 4385 136165 ;
    LAYER V2 ;
      RECT 2505 345 2655 495 ;
    LAYER V2 ;
      RECT 2505 4545 2655 4695 ;
    LAYER V2 ;
      RECT 2505 6225 2655 6375 ;
    LAYER V2 ;
      RECT 2505 10425 2655 10575 ;
    LAYER V2 ;
      RECT 2505 12105 2655 12255 ;
    LAYER V2 ;
      RECT 2505 16305 2655 16455 ;
    LAYER V2 ;
      RECT 2505 17985 2655 18135 ;
    LAYER V2 ;
      RECT 2505 22185 2655 22335 ;
    LAYER V2 ;
      RECT 2505 23865 2655 24015 ;
    LAYER V2 ;
      RECT 2505 28065 2655 28215 ;
    LAYER V2 ;
      RECT 2505 29745 2655 29895 ;
    LAYER V2 ;
      RECT 2505 33945 2655 34095 ;
    LAYER V2 ;
      RECT 2505 35625 2655 35775 ;
    LAYER V2 ;
      RECT 2505 39825 2655 39975 ;
    LAYER V2 ;
      RECT 2505 41505 2655 41655 ;
    LAYER V2 ;
      RECT 2505 45705 2655 45855 ;
    LAYER V2 ;
      RECT 2505 47385 2655 47535 ;
    LAYER V2 ;
      RECT 2505 51585 2655 51735 ;
    LAYER V2 ;
      RECT 2505 53265 2655 53415 ;
    LAYER V2 ;
      RECT 2505 57465 2655 57615 ;
    LAYER V2 ;
      RECT 2505 59145 2655 59295 ;
    LAYER V2 ;
      RECT 2505 63345 2655 63495 ;
    LAYER V2 ;
      RECT 2505 65025 2655 65175 ;
    LAYER V2 ;
      RECT 2505 69225 2655 69375 ;
    LAYER V2 ;
      RECT 2505 70905 2655 71055 ;
    LAYER V2 ;
      RECT 2505 75105 2655 75255 ;
    LAYER V2 ;
      RECT 2505 76785 2655 76935 ;
    LAYER V2 ;
      RECT 2505 80985 2655 81135 ;
    LAYER V2 ;
      RECT 2505 82665 2655 82815 ;
    LAYER V2 ;
      RECT 2505 86865 2655 87015 ;
    LAYER V2 ;
      RECT 2505 88545 2655 88695 ;
    LAYER V2 ;
      RECT 2505 92745 2655 92895 ;
    LAYER V2 ;
      RECT 2505 94425 2655 94575 ;
    LAYER V2 ;
      RECT 2505 98625 2655 98775 ;
    LAYER V2 ;
      RECT 2505 100305 2655 100455 ;
    LAYER V2 ;
      RECT 2505 104505 2655 104655 ;
    LAYER V2 ;
      RECT 2505 106185 2655 106335 ;
    LAYER V2 ;
      RECT 2505 110385 2655 110535 ;
    LAYER V2 ;
      RECT 2505 112065 2655 112215 ;
    LAYER V2 ;
      RECT 2505 116265 2655 116415 ;
    LAYER V2 ;
      RECT 2505 117945 2655 118095 ;
    LAYER V2 ;
      RECT 2505 122145 2655 122295 ;
    LAYER V2 ;
      RECT 2505 123825 2655 123975 ;
    LAYER V2 ;
      RECT 2505 128025 2655 128175 ;
    LAYER V2 ;
      RECT 2505 129705 2655 129855 ;
    LAYER V2 ;
      RECT 2505 133905 2655 134055 ;
    LAYER V2 ;
      RECT 2505 135585 2655 135735 ;
    LAYER V2 ;
      RECT 2505 139785 2655 139935 ;
    LAYER V2 ;
      RECT 2935 765 3085 915 ;
    LAYER V2 ;
      RECT 2935 6645 3085 6795 ;
    LAYER V2 ;
      RECT 2935 12525 3085 12675 ;
    LAYER V2 ;
      RECT 2935 18405 3085 18555 ;
    LAYER V2 ;
      RECT 2935 24285 3085 24435 ;
    LAYER V2 ;
      RECT 2935 30165 3085 30315 ;
    LAYER V2 ;
      RECT 2935 36045 3085 36195 ;
    LAYER V2 ;
      RECT 2935 41925 3085 42075 ;
    LAYER V2 ;
      RECT 2935 47805 3085 47955 ;
    LAYER V2 ;
      RECT 2935 53685 3085 53835 ;
    LAYER V2 ;
      RECT 2935 59565 3085 59715 ;
    LAYER V2 ;
      RECT 2935 65445 3085 65595 ;
    LAYER V2 ;
      RECT 2935 71325 3085 71475 ;
    LAYER V2 ;
      RECT 2935 77205 3085 77355 ;
    LAYER V2 ;
      RECT 2935 83085 3085 83235 ;
    LAYER V2 ;
      RECT 2935 88965 3085 89115 ;
    LAYER V2 ;
      RECT 2935 94845 3085 94995 ;
    LAYER V2 ;
      RECT 2935 100725 3085 100875 ;
    LAYER V2 ;
      RECT 2935 106605 3085 106755 ;
    LAYER V2 ;
      RECT 2935 112485 3085 112635 ;
    LAYER V2 ;
      RECT 2935 118365 3085 118515 ;
    LAYER V2 ;
      RECT 2935 124245 3085 124395 ;
    LAYER V2 ;
      RECT 2935 130125 3085 130275 ;
    LAYER V2 ;
      RECT 2935 136005 3085 136155 ;
    LAYER V2 ;
      RECT 2935 141885 3085 142035 ;
  END
END DCL_NMOS_S_54772057_X4_Y24
