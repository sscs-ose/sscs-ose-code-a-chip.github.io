* SKY130 Spice File.
.include "../../../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice"
.include "../../../cells/nfet_01v8/sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice"
.include "../../../cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice"
.include "../../../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice"
.include "../../../cells/pfet_01v8/sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice"
.include "../../../cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice"
.include "../../../cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice"
.include "../../../cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice"
.include "../../../cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice"
.include "../../../cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice"
.include "../../../cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice"
.include "../../../cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__subvt_mismatch.corner.spice"
.include "../../../cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice"
.include "../../../cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__subvt_mismatch.corner.spice"
.include "../../../cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice"
.include "../../../cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice"
.include "../../../cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__subvt_mismatch.corner.spice"
.include "../../../cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice"
.include "../../../cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice"
.include "../../../cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../../cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice"
.include "../../../cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice"
.include "nonfet.spice"
.include "../../../cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__subvt_mismatch.corner.spice"
.include "../../../cells/nfet_20v0/sky130_fd_pr__nfet_20v0__tt_discrete.corner.spice"
.include "../../../cells/pfet_20v0/sky130_fd_pr__pfet_20v0__tt_discrete.corner.spice"
.include "../../../cells/nfet_20v0_nvt/sky130_fd_pr__nfet_20v0_nvt__tt_discrete.corner.spice"
.include "../../all.spice"
.include "rf.spice"
