# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.130000 BY  3.540000 ;
  PIN BULK
    ANTENNADIFFAREA  2.145000 ;
    ANTENNAGATEAREA  0.495000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.005000 0.500000 2.535000 ;
        RECT 3.630000 1.005000 3.925000 2.535000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.895000 4.060000 2.535000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.188000 ;
    PORT
      LAYER li1 ;
        RECT 1.190000 0.000000 2.940000 0.695000 ;
        RECT 1.190000 2.845000 2.940000 3.540000 ;
      LAYER mcon ;
        RECT 1.260000 0.095000 2.870000 0.625000 ;
        RECT 1.260000 2.915000 2.870000 3.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.180000 0.000000 2.950000 0.685000 ;
        RECT 1.180000 2.855000 2.950000 3.540000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.005000 4.060000 1.645000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 0.800000 2.615000 ;
      RECT 0.580000 0.455000 0.910000 0.785000 ;
      RECT 0.580000 0.785000 0.800000 0.925000 ;
      RECT 0.580000 2.615000 0.800000 2.755000 ;
      RECT 0.580000 2.755000 0.910000 3.085000 ;
      RECT 1.060000 0.925000 1.230000 2.615000 ;
      RECT 1.520000 0.925000 1.690000 2.615000 ;
      RECT 1.980000 0.925000 2.150000 2.615000 ;
      RECT 2.440000 0.925000 2.610000 2.615000 ;
      RECT 2.900000 0.925000 3.070000 2.615000 ;
      RECT 3.220000 0.455000 3.550000 0.785000 ;
      RECT 3.220000 2.755000 3.550000 3.085000 ;
      RECT 3.330000 0.785000 3.550000 0.925000 ;
      RECT 3.330000 0.925000 3.925000 2.615000 ;
      RECT 3.330000 2.615000 3.550000 2.755000 ;
    LAYER mcon ;
      RECT 0.300000 1.145000 0.470000 1.315000 ;
      RECT 0.300000 1.505000 0.470000 1.675000 ;
      RECT 0.300000 1.865000 0.470000 2.035000 ;
      RECT 0.300000 2.225000 0.470000 2.395000 ;
      RECT 1.060000 1.145000 1.230000 1.315000 ;
      RECT 1.060000 1.505000 1.230000 1.675000 ;
      RECT 1.060000 1.865000 1.230000 2.035000 ;
      RECT 1.060000 2.225000 1.230000 2.395000 ;
      RECT 1.520000 1.145000 1.690000 1.315000 ;
      RECT 1.520000 1.505000 1.690000 1.675000 ;
      RECT 1.520000 1.865000 1.690000 2.035000 ;
      RECT 1.520000 2.225000 1.690000 2.395000 ;
      RECT 1.980000 1.145000 2.150000 1.315000 ;
      RECT 1.980000 1.505000 2.150000 1.675000 ;
      RECT 1.980000 1.865000 2.150000 2.035000 ;
      RECT 1.980000 2.225000 2.150000 2.395000 ;
      RECT 2.440000 1.145000 2.610000 1.315000 ;
      RECT 2.440000 1.505000 2.610000 1.675000 ;
      RECT 2.440000 1.865000 2.610000 2.035000 ;
      RECT 2.440000 2.225000 2.610000 2.395000 ;
      RECT 2.900000 1.145000 3.070000 1.315000 ;
      RECT 2.900000 1.505000 3.070000 1.675000 ;
      RECT 2.900000 1.865000 3.070000 2.035000 ;
      RECT 2.900000 2.225000 3.070000 2.395000 ;
      RECT 3.660000 1.145000 3.830000 1.315000 ;
      RECT 3.660000 1.505000 3.830000 1.675000 ;
      RECT 3.660000 1.865000 3.830000 2.035000 ;
      RECT 3.660000 2.225000 3.830000 2.395000 ;
    LAYER met1 ;
      RECT 1.015000 1.005000 1.275000 2.535000 ;
      RECT 1.475000 1.005000 1.735000 2.535000 ;
      RECT 1.935000 1.005000 2.195000 2.535000 ;
      RECT 2.395000 1.005000 2.655000 2.535000 ;
      RECT 2.855000 1.005000 3.115000 2.535000 ;
    LAYER via ;
      RECT 1.015000 1.035000 1.275000 1.295000 ;
      RECT 1.015000 1.355000 1.275000 1.615000 ;
      RECT 1.475000 1.925000 1.735000 2.185000 ;
      RECT 1.475000 2.245000 1.735000 2.505000 ;
      RECT 1.935000 1.035000 2.195000 1.295000 ;
      RECT 1.935000 1.355000 2.195000 1.615000 ;
      RECT 2.395000 1.925000 2.655000 2.185000 ;
      RECT 2.395000 2.245000 2.655000 2.505000 ;
      RECT 2.855000 1.035000 3.115000 1.295000 ;
      RECT 2.855000 1.355000 3.115000 1.615000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18
END LIBRARY
