# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.700000 BY  6.100000 ;
  PIN C0
    PORT
      LAYER met4 ;
        RECT 0.000000 0.630000 0.300000 5.770000 ;
        RECT 0.000000 5.770000 2.700000 6.100000 ;
        RECT 1.200000 0.630000 1.500000 5.770000 ;
        RECT 2.400000 0.630000 2.700000 5.770000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met4 ;
        RECT 0.300000 0.000000 2.400000 0.330000 ;
        RECT 0.600000 0.330000 0.900000 5.470000 ;
        RECT 1.800000 0.330000 2.100000 5.470000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 1.285000 2.860000 1.390000 3.105000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.065000 0.000000 0.235000 6.100000 ;
      RECT 2.465000 0.000000 2.635000 6.100000 ;
    LAYER met1 ;
      RECT 0.070000 0.630000 0.230000 5.770000 ;
      RECT 0.070000 5.770000 2.630000 6.100000 ;
      RECT 0.300000 0.000000 2.400000 0.330000 ;
      RECT 0.370000 0.330000 0.530000 5.470000 ;
      RECT 0.670000 0.630000 0.830000 5.770000 ;
      RECT 0.970000 0.330000 1.130000 5.470000 ;
      RECT 1.270000 0.630000 1.430000 5.770000 ;
      RECT 1.570000 0.330000 1.730000 5.470000 ;
      RECT 1.870000 0.630000 2.030000 5.770000 ;
      RECT 2.170000 0.330000 2.330000 5.470000 ;
      RECT 2.470000 0.630000 2.630000 5.770000 ;
    LAYER met2 ;
      RECT 0.070000 0.630000 0.230000 5.770000 ;
      RECT 0.070000 5.770000 0.830000 6.100000 ;
      RECT 0.300000 0.000000 2.400000 0.330000 ;
      RECT 0.370000 0.330000 0.530000 5.470000 ;
      RECT 0.670000 0.630000 0.830000 5.770000 ;
      RECT 0.970000 0.330000 1.130000 6.100000 ;
      RECT 1.270000 0.630000 1.430000 5.770000 ;
      RECT 1.270000 5.770000 2.630000 6.100000 ;
      RECT 1.570000 0.330000 1.730000 5.470000 ;
      RECT 1.870000 0.630000 2.030000 5.770000 ;
      RECT 2.170000 0.330000 2.330000 5.470000 ;
      RECT 2.470000 0.630000 2.630000 5.770000 ;
    LAYER met3 ;
      RECT 0.000000 0.630000 0.300000 5.770000 ;
      RECT 0.000000 5.770000 2.700000 6.100000 ;
      RECT 0.300000 0.000000 2.400000 0.330000 ;
      RECT 0.600000 0.330000 0.900000 5.470000 ;
      RECT 1.200000 0.630000 1.500000 5.770000 ;
      RECT 1.800000 0.330000 2.100000 5.470000 ;
      RECT 2.400000 0.630000 2.700000 5.770000 ;
    LAYER via ;
      RECT 0.220000 5.805000 0.480000 6.065000 ;
      RECT 0.420000 0.035000 0.680000 0.295000 ;
      RECT 0.820000 0.035000 1.080000 0.295000 ;
      RECT 1.220000 0.035000 1.480000 0.295000 ;
      RECT 1.420000 5.805000 1.680000 6.065000 ;
      RECT 1.620000 0.035000 1.880000 0.295000 ;
      RECT 1.820000 5.805000 2.080000 6.065000 ;
      RECT 2.020000 0.035000 2.280000 0.295000 ;
      RECT 2.220000 5.805000 2.480000 6.065000 ;
    LAYER via2 ;
      RECT 0.210000 5.795000 0.490000 6.075000 ;
      RECT 0.410000 0.025000 0.690000 0.305000 ;
      RECT 0.810000 0.025000 1.090000 0.305000 ;
      RECT 1.210000 0.025000 1.490000 0.305000 ;
      RECT 1.410000 5.795000 1.690000 6.075000 ;
      RECT 1.610000 0.025000 1.890000 0.305000 ;
      RECT 1.810000 5.795000 2.090000 6.075000 ;
      RECT 2.010000 0.025000 2.290000 0.305000 ;
      RECT 2.210000 5.795000 2.490000 6.075000 ;
    LAYER via3 ;
      RECT 0.190000 5.775000 0.510000 6.095000 ;
      RECT 0.390000 0.005000 0.710000 0.325000 ;
      RECT 0.590000 5.775000 0.910000 6.095000 ;
      RECT 0.790000 0.005000 1.110000 0.325000 ;
      RECT 0.990000 5.775000 1.310000 6.095000 ;
      RECT 1.190000 0.005000 1.510000 0.325000 ;
      RECT 1.390000 5.775000 1.710000 6.095000 ;
      RECT 1.590000 0.005000 1.910000 0.325000 ;
      RECT 1.790000 5.775000 2.110000 6.095000 ;
      RECT 1.990000 0.005000 2.310000 0.325000 ;
      RECT 2.190000 5.775000 2.510000 6.095000 ;
  END
END sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap
END LIBRARY
