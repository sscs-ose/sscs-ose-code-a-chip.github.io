MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 50.47 BY 27.64 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 2.8 23.82 3.08 ;
      LAYER M3 ;
        RECT 30.39 2.78 30.67 7.3 ;
      LAYER M2 ;
        RECT 23.65 2.8 25.37 3.08 ;
      LAYER M3 ;
        RECT 25.23 2.94 25.51 3.36 ;
      LAYER M2 ;
        RECT 25.37 3.22 30.53 3.5 ;
      LAYER M3 ;
        RECT 30.39 3.175 30.67 3.545 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 29.96 7.82 30.24 19.9 ;
      LAYER M3 ;
        RECT 38.99 7.82 39.27 19.9 ;
      LAYER M3 ;
        RECT 29.96 13.675 30.24 14.045 ;
      LAYER M4 ;
        RECT 30.1 13.46 39.13 14.26 ;
      LAYER M3 ;
        RECT 38.99 13.675 39.27 14.045 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 37.67 2.8 46.61 3.08 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.27 2.8 12.21 3.08 ;
    END
  END VINP
  OBS 
  LAYER M2 ;
        RECT 37.67 7 46.61 7.28 ;
  LAYER M3 ;
        RECT 47.16 7.82 47.44 18.22 ;
  LAYER M3 ;
        RECT 39.42 12.02 39.7 24.1 ;
  LAYER M2 ;
        RECT 46.44 7 47.3 7.28 ;
  LAYER M3 ;
        RECT 47.16 7.14 47.44 7.98 ;
  LAYER M2 ;
        RECT 39.4 7 39.72 7.28 ;
  LAYER M3 ;
        RECT 39.42 7.14 39.7 12.18 ;
  LAYER M2 ;
        RECT 47.14 7 47.46 7.28 ;
  LAYER M3 ;
        RECT 47.16 6.98 47.44 7.3 ;
  LAYER M2 ;
        RECT 47.14 7 47.46 7.28 ;
  LAYER M3 ;
        RECT 47.16 6.98 47.44 7.3 ;
  LAYER M2 ;
        RECT 39.4 7 39.72 7.28 ;
  LAYER M3 ;
        RECT 39.42 6.98 39.7 7.3 ;
  LAYER M2 ;
        RECT 47.14 7 47.46 7.28 ;
  LAYER M3 ;
        RECT 47.16 6.98 47.44 7.3 ;
  LAYER M2 ;
        RECT 39.4 7 39.72 7.28 ;
  LAYER M3 ;
        RECT 39.42 6.98 39.7 7.3 ;
  LAYER M2 ;
        RECT 47.14 7 47.46 7.28 ;
  LAYER M3 ;
        RECT 47.16 6.98 47.44 7.3 ;
  LAYER M2 ;
        RECT 3.27 7 12.21 7.28 ;
  LAYER M3 ;
        RECT 2.44 7.82 2.72 18.22 ;
  LAYER M3 ;
        RECT 10.18 12.02 10.46 24.1 ;
  LAYER M2 ;
        RECT 2.58 7 3.44 7.28 ;
  LAYER M3 ;
        RECT 2.44 7.14 2.72 7.98 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 7.14 10.46 12.18 ;
  LAYER M2 ;
        RECT 2.42 7 2.74 7.28 ;
  LAYER M3 ;
        RECT 2.44 6.98 2.72 7.3 ;
  LAYER M2 ;
        RECT 2.42 7 2.74 7.28 ;
  LAYER M3 ;
        RECT 2.44 6.98 2.72 7.3 ;
  LAYER M2 ;
        RECT 2.42 7 2.74 7.28 ;
  LAYER M3 ;
        RECT 2.44 6.98 2.72 7.3 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 2.42 7 2.74 7.28 ;
  LAYER M3 ;
        RECT 2.44 6.98 2.72 7.3 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 2.84 6.58 12.64 6.86 ;
  LAYER M2 ;
        RECT 14.88 7 23.82 7.28 ;
  LAYER M3 ;
        RECT 20.07 8.24 20.35 20.32 ;
  LAYER M3 ;
        RECT 29.1 8.24 29.38 20.32 ;
  LAYER M2 ;
        RECT 37.24 6.58 47.04 6.86 ;
  LAYER M2 ;
        RECT 12.47 6.58 13.76 6.86 ;
  LAYER M1 ;
        RECT 13.635 6.72 13.885 7.14 ;
  LAYER M2 ;
        RECT 13.76 7 15.05 7.28 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 7.14 20.35 8.4 ;
  LAYER M2 ;
        RECT 23.65 7 25.37 7.28 ;
  LAYER M3 ;
        RECT 25.23 7.14 25.51 7.56 ;
  LAYER M2 ;
        RECT 25.37 7.42 29.24 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.56 29.38 8.4 ;
  LAYER M2 ;
        RECT 29.24 7.42 36.12 7.7 ;
  LAYER M1 ;
        RECT 35.995 6.72 36.245 7.56 ;
  LAYER M2 ;
        RECT 36.12 6.58 37.41 6.86 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 25.21 7 25.53 7.28 ;
  LAYER M3 ;
        RECT 25.23 6.98 25.51 7.3 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 25.21 7 25.53 7.28 ;
  LAYER M3 ;
        RECT 25.23 6.98 25.51 7.3 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M1 ;
        RECT 35.995 6.635 36.245 6.805 ;
  LAYER M2 ;
        RECT 35.95 6.58 36.29 6.86 ;
  LAYER M1 ;
        RECT 35.995 7.475 36.245 7.645 ;
  LAYER M2 ;
        RECT 35.95 7.42 36.29 7.7 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 25.21 7 25.53 7.28 ;
  LAYER M3 ;
        RECT 25.23 6.98 25.51 7.3 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M1 ;
        RECT 13.635 6.635 13.885 6.805 ;
  LAYER M2 ;
        RECT 13.59 6.58 13.93 6.86 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 7 13.93 7.28 ;
  LAYER M1 ;
        RECT 35.995 6.635 36.245 6.805 ;
  LAYER M2 ;
        RECT 35.95 6.58 36.29 6.86 ;
  LAYER M1 ;
        RECT 35.995 7.475 36.245 7.645 ;
  LAYER M2 ;
        RECT 35.95 7.42 36.29 7.7 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 25.21 7 25.53 7.28 ;
  LAYER M3 ;
        RECT 25.23 6.98 25.51 7.3 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 19.9 ;
  LAYER M3 ;
        RECT 19.64 7.82 19.92 24.1 ;
  LAYER M3 ;
        RECT 29.53 12.02 29.81 24.1 ;
  LAYER M3 ;
        RECT 10.61 15.775 10.89 16.145 ;
  LAYER M2 ;
        RECT 10.75 15.82 19.78 16.1 ;
  LAYER M3 ;
        RECT 19.64 15.775 19.92 16.145 ;
  LAYER M2 ;
        RECT 19.78 15.82 29.67 16.1 ;
  LAYER M3 ;
        RECT 29.53 15.775 29.81 16.145 ;
  LAYER M2 ;
        RECT 10.59 15.82 10.91 16.1 ;
  LAYER M3 ;
        RECT 10.61 15.8 10.89 16.12 ;
  LAYER M2 ;
        RECT 19.62 15.82 19.94 16.1 ;
  LAYER M3 ;
        RECT 19.64 15.8 19.92 16.12 ;
  LAYER M2 ;
        RECT 10.59 15.82 10.91 16.1 ;
  LAYER M3 ;
        RECT 10.61 15.8 10.89 16.12 ;
  LAYER M2 ;
        RECT 19.62 15.82 19.94 16.1 ;
  LAYER M3 ;
        RECT 19.64 15.8 19.92 16.12 ;
  LAYER M2 ;
        RECT 10.59 15.82 10.91 16.1 ;
  LAYER M3 ;
        RECT 10.61 15.8 10.89 16.12 ;
  LAYER M2 ;
        RECT 19.62 15.82 19.94 16.1 ;
  LAYER M3 ;
        RECT 19.64 15.8 19.92 16.12 ;
  LAYER M2 ;
        RECT 29.51 15.82 29.83 16.1 ;
  LAYER M3 ;
        RECT 29.53 15.8 29.81 16.12 ;
  LAYER M2 ;
        RECT 10.59 15.82 10.91 16.1 ;
  LAYER M3 ;
        RECT 10.61 15.8 10.89 16.12 ;
  LAYER M2 ;
        RECT 19.62 15.82 19.94 16.1 ;
  LAYER M3 ;
        RECT 19.64 15.8 19.92 16.12 ;
  LAYER M2 ;
        RECT 29.51 15.82 29.83 16.1 ;
  LAYER M3 ;
        RECT 29.53 15.8 29.81 16.12 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 33.845 3.695 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.845 2.435 34.095 3.445 ;
  LAYER M1 ;
        RECT 33.845 0.335 34.095 1.345 ;
  LAYER M1 ;
        RECT 34.275 3.695 34.525 7.225 ;
  LAYER M1 ;
        RECT 34.705 3.695 34.955 7.225 ;
  LAYER M1 ;
        RECT 34.705 2.435 34.955 3.445 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 1.345 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M2 ;
        RECT 26.06 2.8 35 3.08 ;
  LAYER M2 ;
        RECT 26.06 7 35 7.28 ;
  LAYER M2 ;
        RECT 25.63 6.58 35.43 6.86 ;
  LAYER M2 ;
        RECT 26.06 0.7 35 0.98 ;
  LAYER M3 ;
        RECT 30.39 2.78 30.67 7.3 ;
  LAYER M3 ;
        RECT 30.82 0.68 31.1 6.88 ;
  LAYER M1 ;
        RECT 48.465 7.895 48.715 11.425 ;
  LAYER M1 ;
        RECT 48.465 11.675 48.715 12.685 ;
  LAYER M1 ;
        RECT 48.465 13.775 48.715 17.305 ;
  LAYER M1 ;
        RECT 48.465 17.555 48.715 18.565 ;
  LAYER M1 ;
        RECT 48.465 19.655 48.715 20.665 ;
  LAYER M1 ;
        RECT 48.895 7.895 49.145 11.425 ;
  LAYER M1 ;
        RECT 48.895 13.775 49.145 17.305 ;
  LAYER M1 ;
        RECT 48.035 7.895 48.285 11.425 ;
  LAYER M1 ;
        RECT 48.035 13.775 48.285 17.305 ;
  LAYER M1 ;
        RECT 47.605 7.895 47.855 11.425 ;
  LAYER M1 ;
        RECT 47.605 11.675 47.855 12.685 ;
  LAYER M1 ;
        RECT 47.605 13.775 47.855 17.305 ;
  LAYER M1 ;
        RECT 47.605 17.555 47.855 18.565 ;
  LAYER M1 ;
        RECT 47.605 19.655 47.855 20.665 ;
  LAYER M1 ;
        RECT 47.175 7.895 47.425 11.425 ;
  LAYER M1 ;
        RECT 47.175 13.775 47.425 17.305 ;
  LAYER M1 ;
        RECT 46.745 7.895 46.995 11.425 ;
  LAYER M1 ;
        RECT 46.745 11.675 46.995 12.685 ;
  LAYER M1 ;
        RECT 46.745 13.775 46.995 17.305 ;
  LAYER M1 ;
        RECT 46.745 17.555 46.995 18.565 ;
  LAYER M1 ;
        RECT 46.745 19.655 46.995 20.665 ;
  LAYER M1 ;
        RECT 46.315 7.895 46.565 11.425 ;
  LAYER M1 ;
        RECT 46.315 13.775 46.565 17.305 ;
  LAYER M1 ;
        RECT 45.885 7.895 46.135 11.425 ;
  LAYER M1 ;
        RECT 45.885 11.675 46.135 12.685 ;
  LAYER M1 ;
        RECT 45.885 13.775 46.135 17.305 ;
  LAYER M1 ;
        RECT 45.885 17.555 46.135 18.565 ;
  LAYER M1 ;
        RECT 45.885 19.655 46.135 20.665 ;
  LAYER M1 ;
        RECT 45.455 7.895 45.705 11.425 ;
  LAYER M1 ;
        RECT 45.455 13.775 45.705 17.305 ;
  LAYER M2 ;
        RECT 45.84 12.04 48.76 12.32 ;
  LAYER M2 ;
        RECT 45.84 7.84 48.76 8.12 ;
  LAYER M2 ;
        RECT 45.41 8.26 49.19 8.54 ;
  LAYER M2 ;
        RECT 45.84 17.92 48.76 18.2 ;
  LAYER M2 ;
        RECT 45.84 13.72 48.76 14 ;
  LAYER M2 ;
        RECT 45.41 14.14 49.19 14.42 ;
  LAYER M2 ;
        RECT 45.84 20.02 48.76 20.3 ;
  LAYER M3 ;
        RECT 47.16 7.82 47.44 18.22 ;
  LAYER M3 ;
        RECT 46.73 8.24 47.01 20.32 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 17.305 ;
  LAYER M1 ;
        RECT 1.165 17.555 1.415 18.565 ;
  LAYER M1 ;
        RECT 1.165 19.655 1.415 20.665 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 0.735 13.775 0.985 17.305 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 1.595 13.775 1.845 17.305 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 17.305 ;
  LAYER M1 ;
        RECT 2.025 17.555 2.275 18.565 ;
  LAYER M1 ;
        RECT 2.025 19.655 2.275 20.665 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.455 13.775 2.705 17.305 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 17.305 ;
  LAYER M1 ;
        RECT 2.885 17.555 3.135 18.565 ;
  LAYER M1 ;
        RECT 2.885 19.655 3.135 20.665 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.315 13.775 3.565 17.305 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 17.305 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 19.655 3.995 20.665 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.175 13.775 4.425 17.305 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 0.69 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 1.12 17.92 4.04 18.2 ;
  LAYER M2 ;
        RECT 1.12 13.72 4.04 14 ;
  LAYER M2 ;
        RECT 0.69 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 1.12 20.02 4.04 20.3 ;
  LAYER M3 ;
        RECT 2.44 7.82 2.72 18.22 ;
  LAYER M3 ;
        RECT 2.87 8.24 3.15 20.32 ;
  LAYER M1 ;
        RECT 23.525 3.695 23.775 7.225 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.525 0.335 23.775 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M2 ;
        RECT 14.45 6.58 24.25 6.86 ;
  LAYER M2 ;
        RECT 14.88 0.7 23.82 0.98 ;
  LAYER M2 ;
        RECT 14.88 7 23.82 7.28 ;
  LAYER M2 ;
        RECT 14.88 2.8 23.82 3.08 ;
  LAYER M3 ;
        RECT 18.78 0.68 19.06 6.88 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 17.305 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 19.655 14.315 23.185 ;
  LAYER M1 ;
        RECT 14.065 23.435 14.315 24.445 ;
  LAYER M1 ;
        RECT 14.065 25.535 14.315 26.545 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 17.305 ;
  LAYER M1 ;
        RECT 14.495 19.655 14.745 23.185 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 13.635 19.655 13.885 23.185 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 17.305 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 19.655 13.455 23.185 ;
  LAYER M1 ;
        RECT 13.205 23.435 13.455 24.445 ;
  LAYER M1 ;
        RECT 13.205 25.535 13.455 26.545 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M1 ;
        RECT 12.775 13.775 13.025 17.305 ;
  LAYER M1 ;
        RECT 12.775 19.655 13.025 23.185 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 11.425 ;
  LAYER M1 ;
        RECT 12.345 11.675 12.595 12.685 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 17.305 ;
  LAYER M1 ;
        RECT 12.345 17.555 12.595 18.565 ;
  LAYER M1 ;
        RECT 12.345 19.655 12.595 23.185 ;
  LAYER M1 ;
        RECT 12.345 23.435 12.595 24.445 ;
  LAYER M1 ;
        RECT 12.345 25.535 12.595 26.545 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.915 13.775 12.165 17.305 ;
  LAYER M1 ;
        RECT 11.915 19.655 12.165 23.185 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 17.305 ;
  LAYER M1 ;
        RECT 11.485 17.555 11.735 18.565 ;
  LAYER M1 ;
        RECT 11.485 19.655 11.735 23.185 ;
  LAYER M1 ;
        RECT 11.485 23.435 11.735 24.445 ;
  LAYER M1 ;
        RECT 11.485 25.535 11.735 26.545 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.055 13.775 11.305 17.305 ;
  LAYER M1 ;
        RECT 11.055 19.655 11.305 23.185 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 17.305 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 19.655 10.875 23.185 ;
  LAYER M1 ;
        RECT 10.625 23.435 10.875 24.445 ;
  LAYER M1 ;
        RECT 10.625 25.535 10.875 26.545 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 10.195 13.775 10.445 17.305 ;
  LAYER M1 ;
        RECT 10.195 19.655 10.445 23.185 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 17.305 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 19.655 10.015 23.185 ;
  LAYER M1 ;
        RECT 9.765 23.435 10.015 24.445 ;
  LAYER M1 ;
        RECT 9.765 25.535 10.015 26.545 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 9.335 13.775 9.585 17.305 ;
  LAYER M1 ;
        RECT 9.335 19.655 9.585 23.185 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 17.305 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 19.655 9.155 23.185 ;
  LAYER M1 ;
        RECT 8.905 23.435 9.155 24.445 ;
  LAYER M1 ;
        RECT 8.905 25.535 9.155 26.545 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.475 13.775 8.725 17.305 ;
  LAYER M1 ;
        RECT 8.475 19.655 8.725 23.185 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 17.305 ;
  LAYER M1 ;
        RECT 8.045 17.555 8.295 18.565 ;
  LAYER M1 ;
        RECT 8.045 19.655 8.295 23.185 ;
  LAYER M1 ;
        RECT 8.045 23.435 8.295 24.445 ;
  LAYER M1 ;
        RECT 8.045 25.535 8.295 26.545 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 7.615 19.655 7.865 23.185 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 17.305 ;
  LAYER M1 ;
        RECT 7.185 17.555 7.435 18.565 ;
  LAYER M1 ;
        RECT 7.185 19.655 7.435 23.185 ;
  LAYER M1 ;
        RECT 7.185 23.435 7.435 24.445 ;
  LAYER M1 ;
        RECT 7.185 25.535 7.435 26.545 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.755 13.775 7.005 17.305 ;
  LAYER M1 ;
        RECT 6.755 19.655 7.005 23.185 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 19.655 6.575 23.185 ;
  LAYER M1 ;
        RECT 6.325 23.435 6.575 24.445 ;
  LAYER M1 ;
        RECT 6.325 25.535 6.575 26.545 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 5.895 19.655 6.145 23.185 ;
  LAYER M2 ;
        RECT 6.28 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 14.36 12.32 ;
  LAYER M2 ;
        RECT 5.85 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 6.28 13.72 14.36 14 ;
  LAYER M2 ;
        RECT 6.28 17.92 14.36 18.2 ;
  LAYER M2 ;
        RECT 5.85 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 6.28 19.6 14.36 19.88 ;
  LAYER M2 ;
        RECT 6.28 23.8 14.36 24.08 ;
  LAYER M2 ;
        RECT 5.85 20.02 14.79 20.3 ;
  LAYER M2 ;
        RECT 6.28 25.9 14.36 26.18 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 19.9 ;
  LAYER M3 ;
        RECT 10.18 12.02 10.46 24.1 ;
  LAYER M3 ;
        RECT 9.75 8.24 10.03 26.2 ;
  LAYER M1 ;
        RECT 35.565 7.895 35.815 11.425 ;
  LAYER M1 ;
        RECT 35.565 11.675 35.815 12.685 ;
  LAYER M1 ;
        RECT 35.565 13.775 35.815 17.305 ;
  LAYER M1 ;
        RECT 35.565 17.555 35.815 18.565 ;
  LAYER M1 ;
        RECT 35.565 19.655 35.815 23.185 ;
  LAYER M1 ;
        RECT 35.565 23.435 35.815 24.445 ;
  LAYER M1 ;
        RECT 35.565 25.535 35.815 26.545 ;
  LAYER M1 ;
        RECT 35.135 7.895 35.385 11.425 ;
  LAYER M1 ;
        RECT 35.135 13.775 35.385 17.305 ;
  LAYER M1 ;
        RECT 35.135 19.655 35.385 23.185 ;
  LAYER M1 ;
        RECT 35.995 7.895 36.245 11.425 ;
  LAYER M1 ;
        RECT 35.995 13.775 36.245 17.305 ;
  LAYER M1 ;
        RECT 35.995 19.655 36.245 23.185 ;
  LAYER M1 ;
        RECT 36.425 7.895 36.675 11.425 ;
  LAYER M1 ;
        RECT 36.425 11.675 36.675 12.685 ;
  LAYER M1 ;
        RECT 36.425 13.775 36.675 17.305 ;
  LAYER M1 ;
        RECT 36.425 17.555 36.675 18.565 ;
  LAYER M1 ;
        RECT 36.425 19.655 36.675 23.185 ;
  LAYER M1 ;
        RECT 36.425 23.435 36.675 24.445 ;
  LAYER M1 ;
        RECT 36.425 25.535 36.675 26.545 ;
  LAYER M1 ;
        RECT 36.855 7.895 37.105 11.425 ;
  LAYER M1 ;
        RECT 36.855 13.775 37.105 17.305 ;
  LAYER M1 ;
        RECT 36.855 19.655 37.105 23.185 ;
  LAYER M1 ;
        RECT 37.285 7.895 37.535 11.425 ;
  LAYER M1 ;
        RECT 37.285 11.675 37.535 12.685 ;
  LAYER M1 ;
        RECT 37.285 13.775 37.535 17.305 ;
  LAYER M1 ;
        RECT 37.285 17.555 37.535 18.565 ;
  LAYER M1 ;
        RECT 37.285 19.655 37.535 23.185 ;
  LAYER M1 ;
        RECT 37.285 23.435 37.535 24.445 ;
  LAYER M1 ;
        RECT 37.285 25.535 37.535 26.545 ;
  LAYER M1 ;
        RECT 37.715 7.895 37.965 11.425 ;
  LAYER M1 ;
        RECT 37.715 13.775 37.965 17.305 ;
  LAYER M1 ;
        RECT 37.715 19.655 37.965 23.185 ;
  LAYER M1 ;
        RECT 38.145 7.895 38.395 11.425 ;
  LAYER M1 ;
        RECT 38.145 11.675 38.395 12.685 ;
  LAYER M1 ;
        RECT 38.145 13.775 38.395 17.305 ;
  LAYER M1 ;
        RECT 38.145 17.555 38.395 18.565 ;
  LAYER M1 ;
        RECT 38.145 19.655 38.395 23.185 ;
  LAYER M1 ;
        RECT 38.145 23.435 38.395 24.445 ;
  LAYER M1 ;
        RECT 38.145 25.535 38.395 26.545 ;
  LAYER M1 ;
        RECT 38.575 7.895 38.825 11.425 ;
  LAYER M1 ;
        RECT 38.575 13.775 38.825 17.305 ;
  LAYER M1 ;
        RECT 38.575 19.655 38.825 23.185 ;
  LAYER M1 ;
        RECT 39.005 7.895 39.255 11.425 ;
  LAYER M1 ;
        RECT 39.005 11.675 39.255 12.685 ;
  LAYER M1 ;
        RECT 39.005 13.775 39.255 17.305 ;
  LAYER M1 ;
        RECT 39.005 17.555 39.255 18.565 ;
  LAYER M1 ;
        RECT 39.005 19.655 39.255 23.185 ;
  LAYER M1 ;
        RECT 39.005 23.435 39.255 24.445 ;
  LAYER M1 ;
        RECT 39.005 25.535 39.255 26.545 ;
  LAYER M1 ;
        RECT 39.435 7.895 39.685 11.425 ;
  LAYER M1 ;
        RECT 39.435 13.775 39.685 17.305 ;
  LAYER M1 ;
        RECT 39.435 19.655 39.685 23.185 ;
  LAYER M1 ;
        RECT 39.865 7.895 40.115 11.425 ;
  LAYER M1 ;
        RECT 39.865 11.675 40.115 12.685 ;
  LAYER M1 ;
        RECT 39.865 13.775 40.115 17.305 ;
  LAYER M1 ;
        RECT 39.865 17.555 40.115 18.565 ;
  LAYER M1 ;
        RECT 39.865 19.655 40.115 23.185 ;
  LAYER M1 ;
        RECT 39.865 23.435 40.115 24.445 ;
  LAYER M1 ;
        RECT 39.865 25.535 40.115 26.545 ;
  LAYER M1 ;
        RECT 40.295 7.895 40.545 11.425 ;
  LAYER M1 ;
        RECT 40.295 13.775 40.545 17.305 ;
  LAYER M1 ;
        RECT 40.295 19.655 40.545 23.185 ;
  LAYER M1 ;
        RECT 40.725 7.895 40.975 11.425 ;
  LAYER M1 ;
        RECT 40.725 11.675 40.975 12.685 ;
  LAYER M1 ;
        RECT 40.725 13.775 40.975 17.305 ;
  LAYER M1 ;
        RECT 40.725 17.555 40.975 18.565 ;
  LAYER M1 ;
        RECT 40.725 19.655 40.975 23.185 ;
  LAYER M1 ;
        RECT 40.725 23.435 40.975 24.445 ;
  LAYER M1 ;
        RECT 40.725 25.535 40.975 26.545 ;
  LAYER M1 ;
        RECT 41.155 7.895 41.405 11.425 ;
  LAYER M1 ;
        RECT 41.155 13.775 41.405 17.305 ;
  LAYER M1 ;
        RECT 41.155 19.655 41.405 23.185 ;
  LAYER M1 ;
        RECT 41.585 7.895 41.835 11.425 ;
  LAYER M1 ;
        RECT 41.585 11.675 41.835 12.685 ;
  LAYER M1 ;
        RECT 41.585 13.775 41.835 17.305 ;
  LAYER M1 ;
        RECT 41.585 17.555 41.835 18.565 ;
  LAYER M1 ;
        RECT 41.585 19.655 41.835 23.185 ;
  LAYER M1 ;
        RECT 41.585 23.435 41.835 24.445 ;
  LAYER M1 ;
        RECT 41.585 25.535 41.835 26.545 ;
  LAYER M1 ;
        RECT 42.015 7.895 42.265 11.425 ;
  LAYER M1 ;
        RECT 42.015 13.775 42.265 17.305 ;
  LAYER M1 ;
        RECT 42.015 19.655 42.265 23.185 ;
  LAYER M1 ;
        RECT 42.445 7.895 42.695 11.425 ;
  LAYER M1 ;
        RECT 42.445 11.675 42.695 12.685 ;
  LAYER M1 ;
        RECT 42.445 13.775 42.695 17.305 ;
  LAYER M1 ;
        RECT 42.445 17.555 42.695 18.565 ;
  LAYER M1 ;
        RECT 42.445 19.655 42.695 23.185 ;
  LAYER M1 ;
        RECT 42.445 23.435 42.695 24.445 ;
  LAYER M1 ;
        RECT 42.445 25.535 42.695 26.545 ;
  LAYER M1 ;
        RECT 42.875 7.895 43.125 11.425 ;
  LAYER M1 ;
        RECT 42.875 13.775 43.125 17.305 ;
  LAYER M1 ;
        RECT 42.875 19.655 43.125 23.185 ;
  LAYER M1 ;
        RECT 43.305 7.895 43.555 11.425 ;
  LAYER M1 ;
        RECT 43.305 11.675 43.555 12.685 ;
  LAYER M1 ;
        RECT 43.305 13.775 43.555 17.305 ;
  LAYER M1 ;
        RECT 43.305 17.555 43.555 18.565 ;
  LAYER M1 ;
        RECT 43.305 19.655 43.555 23.185 ;
  LAYER M1 ;
        RECT 43.305 23.435 43.555 24.445 ;
  LAYER M1 ;
        RECT 43.305 25.535 43.555 26.545 ;
  LAYER M1 ;
        RECT 43.735 7.895 43.985 11.425 ;
  LAYER M1 ;
        RECT 43.735 13.775 43.985 17.305 ;
  LAYER M1 ;
        RECT 43.735 19.655 43.985 23.185 ;
  LAYER M2 ;
        RECT 35.52 7.84 43.6 8.12 ;
  LAYER M2 ;
        RECT 35.52 12.04 43.6 12.32 ;
  LAYER M2 ;
        RECT 35.09 8.26 44.03 8.54 ;
  LAYER M2 ;
        RECT 35.52 13.72 43.6 14 ;
  LAYER M2 ;
        RECT 35.52 17.92 43.6 18.2 ;
  LAYER M2 ;
        RECT 35.09 14.14 44.03 14.42 ;
  LAYER M2 ;
        RECT 35.52 19.6 43.6 19.88 ;
  LAYER M2 ;
        RECT 35.52 23.8 43.6 24.08 ;
  LAYER M2 ;
        RECT 35.09 20.02 44.03 20.3 ;
  LAYER M2 ;
        RECT 35.52 25.9 43.6 26.18 ;
  LAYER M3 ;
        RECT 38.99 7.82 39.27 19.9 ;
  LAYER M3 ;
        RECT 39.42 12.02 39.7 24.1 ;
  LAYER M3 ;
        RECT 39.85 8.24 40.13 26.2 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 17.305 ;
  LAYER M1 ;
        RECT 16.645 17.555 16.895 18.565 ;
  LAYER M1 ;
        RECT 16.645 19.655 16.895 23.185 ;
  LAYER M1 ;
        RECT 16.645 23.435 16.895 24.445 ;
  LAYER M1 ;
        RECT 16.645 25.535 16.895 26.545 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.215 13.775 16.465 17.305 ;
  LAYER M1 ;
        RECT 16.215 19.655 16.465 23.185 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M1 ;
        RECT 17.075 19.655 17.325 23.185 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.505 17.555 17.755 18.565 ;
  LAYER M1 ;
        RECT 17.505 19.655 17.755 23.185 ;
  LAYER M1 ;
        RECT 17.505 23.435 17.755 24.445 ;
  LAYER M1 ;
        RECT 17.505 25.535 17.755 26.545 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M1 ;
        RECT 17.935 13.775 18.185 17.305 ;
  LAYER M1 ;
        RECT 17.935 19.655 18.185 23.185 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.365 11.675 18.615 12.685 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 17.305 ;
  LAYER M1 ;
        RECT 18.365 17.555 18.615 18.565 ;
  LAYER M1 ;
        RECT 18.365 19.655 18.615 23.185 ;
  LAYER M1 ;
        RECT 18.365 23.435 18.615 24.445 ;
  LAYER M1 ;
        RECT 18.365 25.535 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 18.795 13.775 19.045 17.305 ;
  LAYER M1 ;
        RECT 18.795 19.655 19.045 23.185 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 17.305 ;
  LAYER M1 ;
        RECT 19.225 17.555 19.475 18.565 ;
  LAYER M1 ;
        RECT 19.225 19.655 19.475 23.185 ;
  LAYER M1 ;
        RECT 19.225 23.435 19.475 24.445 ;
  LAYER M1 ;
        RECT 19.225 25.535 19.475 26.545 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 19.655 13.775 19.905 17.305 ;
  LAYER M1 ;
        RECT 19.655 19.655 19.905 23.185 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M1 ;
        RECT 20.085 11.675 20.335 12.685 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 17.305 ;
  LAYER M1 ;
        RECT 20.085 17.555 20.335 18.565 ;
  LAYER M1 ;
        RECT 20.085 19.655 20.335 23.185 ;
  LAYER M1 ;
        RECT 20.085 23.435 20.335 24.445 ;
  LAYER M1 ;
        RECT 20.085 25.535 20.335 26.545 ;
  LAYER M1 ;
        RECT 20.515 7.895 20.765 11.425 ;
  LAYER M1 ;
        RECT 20.515 13.775 20.765 17.305 ;
  LAYER M1 ;
        RECT 20.515 19.655 20.765 23.185 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 11.425 ;
  LAYER M1 ;
        RECT 20.945 11.675 21.195 12.685 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 17.305 ;
  LAYER M1 ;
        RECT 20.945 17.555 21.195 18.565 ;
  LAYER M1 ;
        RECT 20.945 19.655 21.195 23.185 ;
  LAYER M1 ;
        RECT 20.945 23.435 21.195 24.445 ;
  LAYER M1 ;
        RECT 20.945 25.535 21.195 26.545 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M1 ;
        RECT 21.375 13.775 21.625 17.305 ;
  LAYER M1 ;
        RECT 21.375 19.655 21.625 23.185 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 17.305 ;
  LAYER M1 ;
        RECT 21.805 17.555 22.055 18.565 ;
  LAYER M1 ;
        RECT 21.805 19.655 22.055 23.185 ;
  LAYER M1 ;
        RECT 21.805 23.435 22.055 24.445 ;
  LAYER M1 ;
        RECT 21.805 25.535 22.055 26.545 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 22.235 19.655 22.485 23.185 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 22.665 11.675 22.915 12.685 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 17.305 ;
  LAYER M1 ;
        RECT 22.665 17.555 22.915 18.565 ;
  LAYER M1 ;
        RECT 22.665 19.655 22.915 23.185 ;
  LAYER M1 ;
        RECT 22.665 23.435 22.915 24.445 ;
  LAYER M1 ;
        RECT 22.665 25.535 22.915 26.545 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 23.095 13.775 23.345 17.305 ;
  LAYER M1 ;
        RECT 23.095 19.655 23.345 23.185 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 11.425 ;
  LAYER M1 ;
        RECT 23.525 11.675 23.775 12.685 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 17.305 ;
  LAYER M1 ;
        RECT 23.525 17.555 23.775 18.565 ;
  LAYER M1 ;
        RECT 23.525 19.655 23.775 23.185 ;
  LAYER M1 ;
        RECT 23.525 23.435 23.775 24.445 ;
  LAYER M1 ;
        RECT 23.525 25.535 23.775 26.545 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M1 ;
        RECT 23.955 13.775 24.205 17.305 ;
  LAYER M1 ;
        RECT 23.955 19.655 24.205 23.185 ;
  LAYER M2 ;
        RECT 16.6 12.04 23.82 12.32 ;
  LAYER M2 ;
        RECT 16.6 7.84 23.82 8.12 ;
  LAYER M2 ;
        RECT 16.17 8.26 24.25 8.54 ;
  LAYER M2 ;
        RECT 16.6 17.92 23.82 18.2 ;
  LAYER M2 ;
        RECT 16.6 13.72 23.82 14 ;
  LAYER M2 ;
        RECT 16.17 14.14 24.25 14.42 ;
  LAYER M2 ;
        RECT 16.6 23.8 23.82 24.08 ;
  LAYER M2 ;
        RECT 16.6 19.6 23.82 19.88 ;
  LAYER M2 ;
        RECT 16.17 20.02 24.25 20.3 ;
  LAYER M2 ;
        RECT 16.6 25.9 23.82 26.18 ;
  LAYER M3 ;
        RECT 19.64 7.82 19.92 24.1 ;
  LAYER M3 ;
        RECT 20.07 8.24 20.35 20.32 ;
  LAYER M1 ;
        RECT 46.315 3.695 46.565 7.225 ;
  LAYER M1 ;
        RECT 46.315 2.435 46.565 3.445 ;
  LAYER M1 ;
        RECT 46.315 0.335 46.565 1.345 ;
  LAYER M1 ;
        RECT 46.745 3.695 46.995 7.225 ;
  LAYER M1 ;
        RECT 45.885 3.695 46.135 7.225 ;
  LAYER M1 ;
        RECT 45.455 3.695 45.705 7.225 ;
  LAYER M1 ;
        RECT 45.455 2.435 45.705 3.445 ;
  LAYER M1 ;
        RECT 45.455 0.335 45.705 1.345 ;
  LAYER M1 ;
        RECT 45.025 3.695 45.275 7.225 ;
  LAYER M1 ;
        RECT 44.595 3.695 44.845 7.225 ;
  LAYER M1 ;
        RECT 44.595 2.435 44.845 3.445 ;
  LAYER M1 ;
        RECT 44.595 0.335 44.845 1.345 ;
  LAYER M1 ;
        RECT 44.165 3.695 44.415 7.225 ;
  LAYER M1 ;
        RECT 43.735 3.695 43.985 7.225 ;
  LAYER M1 ;
        RECT 43.735 2.435 43.985 3.445 ;
  LAYER M1 ;
        RECT 43.735 0.335 43.985 1.345 ;
  LAYER M1 ;
        RECT 43.305 3.695 43.555 7.225 ;
  LAYER M1 ;
        RECT 42.875 3.695 43.125 7.225 ;
  LAYER M1 ;
        RECT 42.875 2.435 43.125 3.445 ;
  LAYER M1 ;
        RECT 42.875 0.335 43.125 1.345 ;
  LAYER M1 ;
        RECT 42.445 3.695 42.695 7.225 ;
  LAYER M1 ;
        RECT 42.015 3.695 42.265 7.225 ;
  LAYER M1 ;
        RECT 42.015 2.435 42.265 3.445 ;
  LAYER M1 ;
        RECT 42.015 0.335 42.265 1.345 ;
  LAYER M1 ;
        RECT 41.585 3.695 41.835 7.225 ;
  LAYER M1 ;
        RECT 41.155 3.695 41.405 7.225 ;
  LAYER M1 ;
        RECT 41.155 2.435 41.405 3.445 ;
  LAYER M1 ;
        RECT 41.155 0.335 41.405 1.345 ;
  LAYER M1 ;
        RECT 40.725 3.695 40.975 7.225 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M1 ;
        RECT 40.295 2.435 40.545 3.445 ;
  LAYER M1 ;
        RECT 40.295 0.335 40.545 1.345 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 39.435 2.435 39.685 3.445 ;
  LAYER M1 ;
        RECT 39.435 0.335 39.685 1.345 ;
  LAYER M1 ;
        RECT 39.005 3.695 39.255 7.225 ;
  LAYER M1 ;
        RECT 38.575 3.695 38.825 7.225 ;
  LAYER M1 ;
        RECT 38.575 2.435 38.825 3.445 ;
  LAYER M1 ;
        RECT 38.575 0.335 38.825 1.345 ;
  LAYER M1 ;
        RECT 38.145 3.695 38.395 7.225 ;
  LAYER M1 ;
        RECT 37.715 3.695 37.965 7.225 ;
  LAYER M1 ;
        RECT 37.715 2.435 37.965 3.445 ;
  LAYER M1 ;
        RECT 37.715 0.335 37.965 1.345 ;
  LAYER M1 ;
        RECT 37.285 3.695 37.535 7.225 ;
  LAYER M2 ;
        RECT 37.67 0.7 46.61 0.98 ;
  LAYER M2 ;
        RECT 37.67 7 46.61 7.28 ;
  LAYER M2 ;
        RECT 37.67 2.8 46.61 3.08 ;
  LAYER M2 ;
        RECT 37.24 6.58 47.04 6.86 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.315 2.435 3.565 3.445 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 1.345 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.175 2.435 4.425 3.445 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 1.345 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.035 2.435 5.285 3.445 ;
  LAYER M1 ;
        RECT 5.035 0.335 5.285 1.345 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 5.895 2.435 6.145 3.445 ;
  LAYER M1 ;
        RECT 5.895 0.335 6.145 1.345 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 6.755 2.435 7.005 3.445 ;
  LAYER M1 ;
        RECT 6.755 0.335 7.005 1.345 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.615 2.435 7.865 3.445 ;
  LAYER M1 ;
        RECT 7.615 0.335 7.865 1.345 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.475 2.435 8.725 3.445 ;
  LAYER M1 ;
        RECT 8.475 0.335 8.725 1.345 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.335 2.435 9.585 3.445 ;
  LAYER M1 ;
        RECT 9.335 0.335 9.585 1.345 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.195 2.435 10.445 3.445 ;
  LAYER M1 ;
        RECT 10.195 0.335 10.445 1.345 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.055 2.435 11.305 3.445 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 1.345 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.915 2.435 12.165 3.445 ;
  LAYER M1 ;
        RECT 11.915 0.335 12.165 1.345 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M2 ;
        RECT 3.27 0.7 12.21 0.98 ;
  LAYER M2 ;
        RECT 3.27 7 12.21 7.28 ;
  LAYER M2 ;
        RECT 3.27 2.8 12.21 3.08 ;
  LAYER M2 ;
        RECT 2.84 6.58 12.64 6.86 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 11.425 ;
  LAYER M1 ;
        RECT 32.985 11.675 33.235 12.685 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 17.305 ;
  LAYER M1 ;
        RECT 32.985 17.555 33.235 18.565 ;
  LAYER M1 ;
        RECT 32.985 19.655 33.235 23.185 ;
  LAYER M1 ;
        RECT 32.985 23.435 33.235 24.445 ;
  LAYER M1 ;
        RECT 32.985 25.535 33.235 26.545 ;
  LAYER M1 ;
        RECT 33.415 7.895 33.665 11.425 ;
  LAYER M1 ;
        RECT 33.415 13.775 33.665 17.305 ;
  LAYER M1 ;
        RECT 33.415 19.655 33.665 23.185 ;
  LAYER M1 ;
        RECT 32.555 7.895 32.805 11.425 ;
  LAYER M1 ;
        RECT 32.555 13.775 32.805 17.305 ;
  LAYER M1 ;
        RECT 32.555 19.655 32.805 23.185 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 11.425 ;
  LAYER M1 ;
        RECT 32.125 11.675 32.375 12.685 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 17.305 ;
  LAYER M1 ;
        RECT 32.125 17.555 32.375 18.565 ;
  LAYER M1 ;
        RECT 32.125 19.655 32.375 23.185 ;
  LAYER M1 ;
        RECT 32.125 23.435 32.375 24.445 ;
  LAYER M1 ;
        RECT 32.125 25.535 32.375 26.545 ;
  LAYER M1 ;
        RECT 31.695 7.895 31.945 11.425 ;
  LAYER M1 ;
        RECT 31.695 13.775 31.945 17.305 ;
  LAYER M1 ;
        RECT 31.695 19.655 31.945 23.185 ;
  LAYER M1 ;
        RECT 31.265 7.895 31.515 11.425 ;
  LAYER M1 ;
        RECT 31.265 11.675 31.515 12.685 ;
  LAYER M1 ;
        RECT 31.265 13.775 31.515 17.305 ;
  LAYER M1 ;
        RECT 31.265 17.555 31.515 18.565 ;
  LAYER M1 ;
        RECT 31.265 19.655 31.515 23.185 ;
  LAYER M1 ;
        RECT 31.265 23.435 31.515 24.445 ;
  LAYER M1 ;
        RECT 31.265 25.535 31.515 26.545 ;
  LAYER M1 ;
        RECT 30.835 7.895 31.085 11.425 ;
  LAYER M1 ;
        RECT 30.835 13.775 31.085 17.305 ;
  LAYER M1 ;
        RECT 30.835 19.655 31.085 23.185 ;
  LAYER M1 ;
        RECT 30.405 7.895 30.655 11.425 ;
  LAYER M1 ;
        RECT 30.405 11.675 30.655 12.685 ;
  LAYER M1 ;
        RECT 30.405 13.775 30.655 17.305 ;
  LAYER M1 ;
        RECT 30.405 17.555 30.655 18.565 ;
  LAYER M1 ;
        RECT 30.405 19.655 30.655 23.185 ;
  LAYER M1 ;
        RECT 30.405 23.435 30.655 24.445 ;
  LAYER M1 ;
        RECT 30.405 25.535 30.655 26.545 ;
  LAYER M1 ;
        RECT 29.975 7.895 30.225 11.425 ;
  LAYER M1 ;
        RECT 29.975 13.775 30.225 17.305 ;
  LAYER M1 ;
        RECT 29.975 19.655 30.225 23.185 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 11.425 ;
  LAYER M1 ;
        RECT 29.545 11.675 29.795 12.685 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 17.305 ;
  LAYER M1 ;
        RECT 29.545 17.555 29.795 18.565 ;
  LAYER M1 ;
        RECT 29.545 19.655 29.795 23.185 ;
  LAYER M1 ;
        RECT 29.545 23.435 29.795 24.445 ;
  LAYER M1 ;
        RECT 29.545 25.535 29.795 26.545 ;
  LAYER M1 ;
        RECT 29.115 7.895 29.365 11.425 ;
  LAYER M1 ;
        RECT 29.115 13.775 29.365 17.305 ;
  LAYER M1 ;
        RECT 29.115 19.655 29.365 23.185 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 11.425 ;
  LAYER M1 ;
        RECT 28.685 11.675 28.935 12.685 ;
  LAYER M1 ;
        RECT 28.685 13.775 28.935 17.305 ;
  LAYER M1 ;
        RECT 28.685 17.555 28.935 18.565 ;
  LAYER M1 ;
        RECT 28.685 19.655 28.935 23.185 ;
  LAYER M1 ;
        RECT 28.685 23.435 28.935 24.445 ;
  LAYER M1 ;
        RECT 28.685 25.535 28.935 26.545 ;
  LAYER M1 ;
        RECT 28.255 7.895 28.505 11.425 ;
  LAYER M1 ;
        RECT 28.255 13.775 28.505 17.305 ;
  LAYER M1 ;
        RECT 28.255 19.655 28.505 23.185 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 11.425 ;
  LAYER M1 ;
        RECT 27.825 11.675 28.075 12.685 ;
  LAYER M1 ;
        RECT 27.825 13.775 28.075 17.305 ;
  LAYER M1 ;
        RECT 27.825 17.555 28.075 18.565 ;
  LAYER M1 ;
        RECT 27.825 19.655 28.075 23.185 ;
  LAYER M1 ;
        RECT 27.825 23.435 28.075 24.445 ;
  LAYER M1 ;
        RECT 27.825 25.535 28.075 26.545 ;
  LAYER M1 ;
        RECT 27.395 7.895 27.645 11.425 ;
  LAYER M1 ;
        RECT 27.395 13.775 27.645 17.305 ;
  LAYER M1 ;
        RECT 27.395 19.655 27.645 23.185 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 11.425 ;
  LAYER M1 ;
        RECT 26.965 11.675 27.215 12.685 ;
  LAYER M1 ;
        RECT 26.965 13.775 27.215 17.305 ;
  LAYER M1 ;
        RECT 26.965 17.555 27.215 18.565 ;
  LAYER M1 ;
        RECT 26.965 19.655 27.215 23.185 ;
  LAYER M1 ;
        RECT 26.965 23.435 27.215 24.445 ;
  LAYER M1 ;
        RECT 26.965 25.535 27.215 26.545 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M1 ;
        RECT 26.535 13.775 26.785 17.305 ;
  LAYER M1 ;
        RECT 26.535 19.655 26.785 23.185 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 11.425 ;
  LAYER M1 ;
        RECT 26.105 11.675 26.355 12.685 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 17.305 ;
  LAYER M1 ;
        RECT 26.105 17.555 26.355 18.565 ;
  LAYER M1 ;
        RECT 26.105 19.655 26.355 23.185 ;
  LAYER M1 ;
        RECT 26.105 23.435 26.355 24.445 ;
  LAYER M1 ;
        RECT 26.105 25.535 26.355 26.545 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 25.675 13.775 25.925 17.305 ;
  LAYER M1 ;
        RECT 25.675 19.655 25.925 23.185 ;
  LAYER M2 ;
        RECT 26.06 7.84 33.28 8.12 ;
  LAYER M2 ;
        RECT 26.06 12.04 33.28 12.32 ;
  LAYER M2 ;
        RECT 25.63 8.26 33.71 8.54 ;
  LAYER M2 ;
        RECT 26.06 13.72 33.28 14 ;
  LAYER M2 ;
        RECT 26.06 17.92 33.28 18.2 ;
  LAYER M2 ;
        RECT 25.63 14.14 33.71 14.42 ;
  LAYER M2 ;
        RECT 26.06 19.6 33.28 19.88 ;
  LAYER M2 ;
        RECT 26.06 23.8 33.28 24.08 ;
  LAYER M2 ;
        RECT 25.63 20.02 33.71 20.3 ;
  LAYER M2 ;
        RECT 26.06 25.9 33.28 26.18 ;
  LAYER M3 ;
        RECT 29.96 7.82 30.24 19.9 ;
  LAYER M3 ;
        RECT 29.53 12.02 29.81 24.1 ;
  LAYER M3 ;
        RECT 29.1 8.24 29.38 20.32 ;
  END 
END CURRENT_MIRROR_OTA
