* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 9
.param
+ sky130_fd_pr__nfet_03v3_nvt__toxe_mult = 0.9635
+ sky130_fd_pr__nfet_03v3_nvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_03v3_nvt__overlap_mult = 0.51025
+ sky130_fd_pr__nfet_03v3_nvt__ajunction_mult = 0.68772
+ sky130_fd_pr__nfet_03v3_nvt__pjunction_mult = 0.9019
+ sky130_fd_pr__nfet_03v3_nvt__lint_diff = 1.21275e-8
+ sky130_fd_pr__nfet_03v3_nvt__wint_diff = -2.252e-8
+ sky130_fd_pr__nfet_03v3_nvt__dlc_diff = 1.6112e-8
+ sky130_fd_pr__nfet_03v3_nvt__dwc_diff = -2.252e-8
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_0 = 0.017139
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_0 = -0.016856
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0 = -1.0949
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0 = -0.041263
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_0 = 0.00079908
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0 = -1877.8
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_0 = -8.8355e-20
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_0 = 1.2237e-11
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_1 = 3.5287e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_1 = 0.010252
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_1 = -0.00051272
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1 = -1.3847
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1 = -0.0485
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_1 = -7.0468e-5
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1 = -9793.6
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_1 = 2.2579e-19
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_2 = 1.2013e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_2 = 1.1421e-10
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_2 = 0.0012159
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2 = -0.49031
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2 = -0.034235
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_2 = 0.0043842
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2 = -8139.1
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_2 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_3 = 6.5751e-20
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_3 = 2.2944e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_3 = 0.0177
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_3 = -0.01428
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3 = -1.0283
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3 = -0.04376
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_3 = 0.0014903
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3 = -3761.4
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_3 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_4 = -4.2142e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_4 = -1.3052e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_4 = 0.044934
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_4 = 0.0083971
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4 = -1.5502
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4 = -0.068861
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_4 = 0.0016304
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4 = -6110.3
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_5 = 0.01509
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5 = -5015.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_5 = 2.0257e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_5 = 4.4064e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_5 = 0.0059498
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5 = -1.6314
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5 = 0.014604
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6 = -0.77252
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6 = -0.0039098
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_6 = 0.011371
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6 = -3438.4
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_6 = 1.7785e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_6 = 5.037e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_6 = 0.0058775
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_7 = 0.021791
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_7 = 0.0022917
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7 = -1.3041
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7 = -0.046002
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_7 = 0.00087134
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7 = -9538.4
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_7 = 4.1235e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_7 = 2.4503e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_7 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_8 = 0.0038297
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8 = -0.51817
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8 = -0.040702
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_8 = 0.006163
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8 = -7789.7
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_8 = 1.381e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_8 = 1.3573e-10
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8 = 0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"
