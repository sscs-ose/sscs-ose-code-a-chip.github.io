MACRO SCM_NMOS_B_90984876_X11_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_90984876_X11_Y1 0 0 ;
  SIZE 20640 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 19520 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 9750 260 10030 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 700 19520 980 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 19950 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 7225 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 7225 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 7225 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 7225 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 7225 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 7225 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 7225 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 7225 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 7225 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 7225 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 7225 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 7225 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 7225 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 7225 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 7225 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 7225 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 7225 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 7225 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 7225 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M2 ;
      RECT 1120 4480 19520 4760 ;
    LAYER M2 ;
      RECT 1120 280 18660 560 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 3785 755 3955 925 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6635 3955 6805 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 5505 755 5675 925 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6635 5675 6805 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6635 6535 6805 ;
    LAYER V1 ;
      RECT 7225 755 7395 925 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6635 7395 6805 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6635 8255 6805 ;
    LAYER V1 ;
      RECT 8945 755 9115 925 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6635 9115 6805 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6635 9975 6805 ;
    LAYER V1 ;
      RECT 10665 755 10835 925 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6635 10835 6805 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6635 11695 6805 ;
    LAYER V1 ;
      RECT 12385 755 12555 925 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6635 12555 6805 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6635 13415 6805 ;
    LAYER V1 ;
      RECT 14105 755 14275 925 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6635 14275 6805 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6635 15135 6805 ;
    LAYER V1 ;
      RECT 15825 755 15995 925 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6635 15995 6805 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6635 16855 6805 ;
    LAYER V1 ;
      RECT 17545 755 17715 925 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6635 17715 6805 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6635 18575 6805 ;
    LAYER V1 ;
      RECT 19265 755 19435 925 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6635 19435 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 3355 1175 3525 1345 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 5075 1175 5245 1345 ;
    LAYER V1 ;
      RECT 5935 1175 6105 1345 ;
    LAYER V1 ;
      RECT 6795 1175 6965 1345 ;
    LAYER V1 ;
      RECT 7655 1175 7825 1345 ;
    LAYER V1 ;
      RECT 8515 1175 8685 1345 ;
    LAYER V1 ;
      RECT 9375 1175 9545 1345 ;
    LAYER V1 ;
      RECT 10235 1175 10405 1345 ;
    LAYER V1 ;
      RECT 11095 1175 11265 1345 ;
    LAYER V1 ;
      RECT 11955 1175 12125 1345 ;
    LAYER V1 ;
      RECT 12815 1175 12985 1345 ;
    LAYER V1 ;
      RECT 13675 1175 13845 1345 ;
    LAYER V1 ;
      RECT 14535 1175 14705 1345 ;
    LAYER V1 ;
      RECT 15395 1175 15565 1345 ;
    LAYER V1 ;
      RECT 16255 1175 16425 1345 ;
    LAYER V1 ;
      RECT 17115 1175 17285 1345 ;
    LAYER V1 ;
      RECT 17975 1175 18145 1345 ;
    LAYER V1 ;
      RECT 18835 1175 19005 1345 ;
    LAYER V1 ;
      RECT 19695 1175 19865 1345 ;
    LAYER V2 ;
      RECT 9815 345 9965 495 ;
    LAYER V2 ;
      RECT 9815 4545 9965 4695 ;
  END
END SCM_NMOS_B_90984876_X11_Y1
