# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_npn_05v5_W5p00L5p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_npn_05v5_W5p00L5p00 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  13.70000 BY  13.70000 ;
  OBS
    LAYER li1 ;
      RECT  0.170000  0.170000 13.790000  0.500000 ;
      RECT  0.170000  0.500000  0.500000 13.460000 ;
      RECT  0.170000 13.460000 13.790000 13.790000 ;
      RECT  1.300000  1.300000 12.660000  1.630000 ;
      RECT  1.300000  1.630000  1.630000 12.330000 ;
      RECT  1.300000 12.330000 12.660000 12.660000 ;
      RECT  3.310000  3.310000 10.650000  3.640000 ;
      RECT  3.310000  3.640000  3.640000 10.320000 ;
      RECT  3.310000 10.320000 10.650000 10.650000 ;
      RECT  4.605000  4.605000  9.355000  9.355000 ;
      RECT 10.320000  3.640000 10.650000 10.320000 ;
      RECT 12.330000  1.630000 12.660000 12.330000 ;
      RECT 13.460000  0.500000 13.790000 13.460000 ;
    LAYER mcon ;
      RECT  0.250000  0.250000  0.420000  0.420000 ;
      RECT  0.250000  0.775000  0.420000  0.945000 ;
      RECT  0.250000  1.135000  0.420000  1.305000 ;
      RECT  0.250000  1.495000  0.420000  1.665000 ;
      RECT  0.250000  1.855000  0.420000  2.025000 ;
      RECT  0.250000  2.215000  0.420000  2.385000 ;
      RECT  0.250000  2.575000  0.420000  2.745000 ;
      RECT  0.250000  2.935000  0.420000  3.105000 ;
      RECT  0.250000  3.295000  0.420000  3.465000 ;
      RECT  0.250000  3.655000  0.420000  3.825000 ;
      RECT  0.250000  4.015000  0.420000  4.185000 ;
      RECT  0.250000  4.375000  0.420000  4.545000 ;
      RECT  0.250000  4.735000  0.420000  4.905000 ;
      RECT  0.250000  5.095000  0.420000  5.265000 ;
      RECT  0.250000  5.455000  0.420000  5.625000 ;
      RECT  0.250000  5.815000  0.420000  5.985000 ;
      RECT  0.250000  6.175000  0.420000  6.345000 ;
      RECT  0.250000  6.535000  0.420000  6.705000 ;
      RECT  0.250000  6.895000  0.420000  7.065000 ;
      RECT  0.250000  7.255000  0.420000  7.425000 ;
      RECT  0.250000  7.615000  0.420000  7.785000 ;
      RECT  0.250000  7.975000  0.420000  8.145000 ;
      RECT  0.250000  8.335000  0.420000  8.505000 ;
      RECT  0.250000  8.695000  0.420000  8.865000 ;
      RECT  0.250000  9.055000  0.420000  9.225000 ;
      RECT  0.250000  9.415000  0.420000  9.585000 ;
      RECT  0.250000  9.775000  0.420000  9.945000 ;
      RECT  0.250000 10.135000  0.420000 10.305000 ;
      RECT  0.250000 10.495000  0.420000 10.665000 ;
      RECT  0.250000 10.855000  0.420000 11.025000 ;
      RECT  0.250000 11.215000  0.420000 11.385000 ;
      RECT  0.250000 11.575000  0.420000 11.745000 ;
      RECT  0.250000 11.935000  0.420000 12.105000 ;
      RECT  0.250000 12.295000  0.420000 12.465000 ;
      RECT  0.250000 12.655000  0.420000 12.825000 ;
      RECT  0.250000 13.015000  0.420000 13.185000 ;
      RECT  0.250000 13.540000  0.420000 13.710000 ;
      RECT  0.775000  0.250000  0.945000  0.420000 ;
      RECT  0.775000 13.540000  0.945000 13.710000 ;
      RECT  1.135000  0.250000  1.305000  0.420000 ;
      RECT  1.135000 13.540000  1.305000 13.710000 ;
      RECT  1.380000  1.380000  1.550000  1.550000 ;
      RECT  1.380000  1.855000  1.550000  2.025000 ;
      RECT  1.380000  2.215000  1.550000  2.385000 ;
      RECT  1.380000  2.575000  1.550000  2.745000 ;
      RECT  1.380000  2.935000  1.550000  3.105000 ;
      RECT  1.380000  3.295000  1.550000  3.465000 ;
      RECT  1.380000  3.655000  1.550000  3.825000 ;
      RECT  1.380000  4.015000  1.550000  4.185000 ;
      RECT  1.380000  4.375000  1.550000  4.545000 ;
      RECT  1.380000  4.735000  1.550000  4.905000 ;
      RECT  1.380000  5.095000  1.550000  5.265000 ;
      RECT  1.380000  5.455000  1.550000  5.625000 ;
      RECT  1.380000  5.815000  1.550000  5.985000 ;
      RECT  1.380000  6.175000  1.550000  6.345000 ;
      RECT  1.380000  6.535000  1.550000  6.705000 ;
      RECT  1.380000  6.895000  1.550000  7.065000 ;
      RECT  1.380000  7.255000  1.550000  7.425000 ;
      RECT  1.380000  7.615000  1.550000  7.785000 ;
      RECT  1.380000  7.975000  1.550000  8.145000 ;
      RECT  1.380000  8.335000  1.550000  8.505000 ;
      RECT  1.380000  8.695000  1.550000  8.865000 ;
      RECT  1.380000  9.055000  1.550000  9.225000 ;
      RECT  1.380000  9.415000  1.550000  9.585000 ;
      RECT  1.380000  9.775000  1.550000  9.945000 ;
      RECT  1.380000 10.135000  1.550000 10.305000 ;
      RECT  1.380000 10.495000  1.550000 10.665000 ;
      RECT  1.380000 10.855000  1.550000 11.025000 ;
      RECT  1.380000 11.215000  1.550000 11.385000 ;
      RECT  1.380000 11.575000  1.550000 11.745000 ;
      RECT  1.380000 11.935000  1.550000 12.105000 ;
      RECT  1.380000 12.410000  1.550000 12.580000 ;
      RECT  1.495000  0.250000  1.665000  0.420000 ;
      RECT  1.495000 13.540000  1.665000 13.710000 ;
      RECT  1.855000  0.250000  2.025000  0.420000 ;
      RECT  1.855000  1.380000  2.025000  1.550000 ;
      RECT  1.855000 12.410000  2.025000 12.580000 ;
      RECT  1.855000 13.540000  2.025000 13.710000 ;
      RECT  2.215000  0.250000  2.385000  0.420000 ;
      RECT  2.215000  1.380000  2.385000  1.550000 ;
      RECT  2.215000 12.410000  2.385000 12.580000 ;
      RECT  2.215000 13.540000  2.385000 13.710000 ;
      RECT  2.575000  0.250000  2.745000  0.420000 ;
      RECT  2.575000  1.380000  2.745000  1.550000 ;
      RECT  2.575000 12.410000  2.745000 12.580000 ;
      RECT  2.575000 13.540000  2.745000 13.710000 ;
      RECT  2.935000  0.250000  3.105000  0.420000 ;
      RECT  2.935000  1.380000  3.105000  1.550000 ;
      RECT  2.935000 12.410000  3.105000 12.580000 ;
      RECT  2.935000 13.540000  3.105000 13.710000 ;
      RECT  3.295000  0.250000  3.465000  0.420000 ;
      RECT  3.295000  1.380000  3.465000  1.550000 ;
      RECT  3.295000 12.410000  3.465000 12.580000 ;
      RECT  3.295000 13.540000  3.465000 13.710000 ;
      RECT  3.390000  3.390000  3.560000  3.560000 ;
      RECT  3.390000  3.835000  3.560000  4.005000 ;
      RECT  3.390000  4.195000  3.560000  4.365000 ;
      RECT  3.390000  4.555000  3.560000  4.725000 ;
      RECT  3.390000  4.915000  3.560000  5.085000 ;
      RECT  3.390000  5.275000  3.560000  5.445000 ;
      RECT  3.390000  5.635000  3.560000  5.805000 ;
      RECT  3.390000  5.995000  3.560000  6.165000 ;
      RECT  3.390000  6.355000  3.560000  6.525000 ;
      RECT  3.390000  6.715000  3.560000  6.885000 ;
      RECT  3.390000  7.075000  3.560000  7.245000 ;
      RECT  3.390000  7.435000  3.560000  7.605000 ;
      RECT  3.390000  7.795000  3.560000  7.965000 ;
      RECT  3.390000  8.155000  3.560000  8.325000 ;
      RECT  3.390000  8.515000  3.560000  8.685000 ;
      RECT  3.390000  8.875000  3.560000  9.045000 ;
      RECT  3.390000  9.235000  3.560000  9.405000 ;
      RECT  3.390000  9.595000  3.560000  9.765000 ;
      RECT  3.390000  9.955000  3.560000 10.125000 ;
      RECT  3.390000 10.400000  3.560000 10.570000 ;
      RECT  3.655000  0.250000  3.825000  0.420000 ;
      RECT  3.655000  1.380000  3.825000  1.550000 ;
      RECT  3.655000 12.410000  3.825000 12.580000 ;
      RECT  3.655000 13.540000  3.825000 13.710000 ;
      RECT  3.835000  3.390000  4.005000  3.560000 ;
      RECT  3.835000 10.400000  4.005000 10.570000 ;
      RECT  4.015000  0.250000  4.185000  0.420000 ;
      RECT  4.015000  1.380000  4.185000  1.550000 ;
      RECT  4.015000 12.410000  4.185000 12.580000 ;
      RECT  4.015000 13.540000  4.185000 13.710000 ;
      RECT  4.195000  3.390000  4.365000  3.560000 ;
      RECT  4.195000 10.400000  4.365000 10.570000 ;
      RECT  4.375000  0.250000  4.545000  0.420000 ;
      RECT  4.375000  1.380000  4.545000  1.550000 ;
      RECT  4.375000 12.410000  4.545000 12.580000 ;
      RECT  4.375000 13.540000  4.545000 13.710000 ;
      RECT  4.555000  3.390000  4.725000  3.560000 ;
      RECT  4.555000 10.400000  4.725000 10.570000 ;
      RECT  4.735000  0.250000  4.905000  0.420000 ;
      RECT  4.735000  1.380000  4.905000  1.550000 ;
      RECT  4.735000  4.735000  9.225000  9.225000 ;
      RECT  4.735000 12.410000  4.905000 12.580000 ;
      RECT  4.735000 13.540000  4.905000 13.710000 ;
      RECT  4.915000  3.390000  5.085000  3.560000 ;
      RECT  4.915000 10.400000  5.085000 10.570000 ;
      RECT  5.095000  0.250000  5.265000  0.420000 ;
      RECT  5.095000  1.380000  5.265000  1.550000 ;
      RECT  5.095000 12.410000  5.265000 12.580000 ;
      RECT  5.095000 13.540000  5.265000 13.710000 ;
      RECT  5.275000  3.390000  5.445000  3.560000 ;
      RECT  5.275000 10.400000  5.445000 10.570000 ;
      RECT  5.455000  0.250000  5.625000  0.420000 ;
      RECT  5.455000  1.380000  5.625000  1.550000 ;
      RECT  5.455000 12.410000  5.625000 12.580000 ;
      RECT  5.455000 13.540000  5.625000 13.710000 ;
      RECT  5.635000  3.390000  5.805000  3.560000 ;
      RECT  5.635000 10.400000  5.805000 10.570000 ;
      RECT  5.815000  0.250000  5.985000  0.420000 ;
      RECT  5.815000  1.380000  5.985000  1.550000 ;
      RECT  5.815000 12.410000  5.985000 12.580000 ;
      RECT  5.815000 13.540000  5.985000 13.710000 ;
      RECT  5.995000  3.390000  6.165000  3.560000 ;
      RECT  5.995000 10.400000  6.165000 10.570000 ;
      RECT  6.175000  0.250000  6.345000  0.420000 ;
      RECT  6.175000  1.380000  6.345000  1.550000 ;
      RECT  6.175000 12.410000  6.345000 12.580000 ;
      RECT  6.175000 13.540000  6.345000 13.710000 ;
      RECT  6.355000  3.390000  6.525000  3.560000 ;
      RECT  6.355000 10.400000  6.525000 10.570000 ;
      RECT  6.535000  0.250000  6.705000  0.420000 ;
      RECT  6.535000  1.380000  6.705000  1.550000 ;
      RECT  6.535000 12.410000  6.705000 12.580000 ;
      RECT  6.535000 13.540000  6.705000 13.710000 ;
      RECT  6.715000  3.390000  6.885000  3.560000 ;
      RECT  6.715000 10.400000  6.885000 10.570000 ;
      RECT  6.895000  0.250000  7.065000  0.420000 ;
      RECT  6.895000  1.380000  7.065000  1.550000 ;
      RECT  6.895000 12.410000  7.065000 12.580000 ;
      RECT  6.895000 13.540000  7.065000 13.710000 ;
      RECT  7.075000  3.390000  7.245000  3.560000 ;
      RECT  7.075000 10.400000  7.245000 10.570000 ;
      RECT  7.255000  0.250000  7.425000  0.420000 ;
      RECT  7.255000  1.380000  7.425000  1.550000 ;
      RECT  7.255000 12.410000  7.425000 12.580000 ;
      RECT  7.255000 13.540000  7.425000 13.710000 ;
      RECT  7.435000  3.390000  7.605000  3.560000 ;
      RECT  7.435000 10.400000  7.605000 10.570000 ;
      RECT  7.615000  0.250000  7.785000  0.420000 ;
      RECT  7.615000  1.380000  7.785000  1.550000 ;
      RECT  7.615000 12.410000  7.785000 12.580000 ;
      RECT  7.615000 13.540000  7.785000 13.710000 ;
      RECT  7.795000  3.390000  7.965000  3.560000 ;
      RECT  7.795000 10.400000  7.965000 10.570000 ;
      RECT  7.975000  0.250000  8.145000  0.420000 ;
      RECT  7.975000  1.380000  8.145000  1.550000 ;
      RECT  7.975000 12.410000  8.145000 12.580000 ;
      RECT  7.975000 13.540000  8.145000 13.710000 ;
      RECT  8.155000  3.390000  8.325000  3.560000 ;
      RECT  8.155000 10.400000  8.325000 10.570000 ;
      RECT  8.335000  0.250000  8.505000  0.420000 ;
      RECT  8.335000  1.380000  8.505000  1.550000 ;
      RECT  8.335000 12.410000  8.505000 12.580000 ;
      RECT  8.335000 13.540000  8.505000 13.710000 ;
      RECT  8.515000  3.390000  8.685000  3.560000 ;
      RECT  8.515000 10.400000  8.685000 10.570000 ;
      RECT  8.695000  0.250000  8.865000  0.420000 ;
      RECT  8.695000  1.380000  8.865000  1.550000 ;
      RECT  8.695000 12.410000  8.865000 12.580000 ;
      RECT  8.695000 13.540000  8.865000 13.710000 ;
      RECT  8.875000  3.390000  9.045000  3.560000 ;
      RECT  8.875000 10.400000  9.045000 10.570000 ;
      RECT  9.055000  0.250000  9.225000  0.420000 ;
      RECT  9.055000  1.380000  9.225000  1.550000 ;
      RECT  9.055000 12.410000  9.225000 12.580000 ;
      RECT  9.055000 13.540000  9.225000 13.710000 ;
      RECT  9.235000  3.390000  9.405000  3.560000 ;
      RECT  9.235000 10.400000  9.405000 10.570000 ;
      RECT  9.415000  0.250000  9.585000  0.420000 ;
      RECT  9.415000  1.380000  9.585000  1.550000 ;
      RECT  9.415000 12.410000  9.585000 12.580000 ;
      RECT  9.415000 13.540000  9.585000 13.710000 ;
      RECT  9.595000  3.390000  9.765000  3.560000 ;
      RECT  9.595000 10.400000  9.765000 10.570000 ;
      RECT  9.775000  0.250000  9.945000  0.420000 ;
      RECT  9.775000  1.380000  9.945000  1.550000 ;
      RECT  9.775000 12.410000  9.945000 12.580000 ;
      RECT  9.775000 13.540000  9.945000 13.710000 ;
      RECT  9.955000  3.390000 10.125000  3.560000 ;
      RECT  9.955000 10.400000 10.125000 10.570000 ;
      RECT 10.135000  0.250000 10.305000  0.420000 ;
      RECT 10.135000  1.380000 10.305000  1.550000 ;
      RECT 10.135000 12.410000 10.305000 12.580000 ;
      RECT 10.135000 13.540000 10.305000 13.710000 ;
      RECT 10.400000  3.390000 10.570000  3.560000 ;
      RECT 10.400000  3.835000 10.570000  4.005000 ;
      RECT 10.400000  4.195000 10.570000  4.365000 ;
      RECT 10.400000  4.555000 10.570000  4.725000 ;
      RECT 10.400000  4.915000 10.570000  5.085000 ;
      RECT 10.400000  5.275000 10.570000  5.445000 ;
      RECT 10.400000  5.635000 10.570000  5.805000 ;
      RECT 10.400000  5.995000 10.570000  6.165000 ;
      RECT 10.400000  6.355000 10.570000  6.525000 ;
      RECT 10.400000  6.715000 10.570000  6.885000 ;
      RECT 10.400000  7.075000 10.570000  7.245000 ;
      RECT 10.400000  7.435000 10.570000  7.605000 ;
      RECT 10.400000  7.795000 10.570000  7.965000 ;
      RECT 10.400000  8.155000 10.570000  8.325000 ;
      RECT 10.400000  8.515000 10.570000  8.685000 ;
      RECT 10.400000  8.875000 10.570000  9.045000 ;
      RECT 10.400000  9.235000 10.570000  9.405000 ;
      RECT 10.400000  9.595000 10.570000  9.765000 ;
      RECT 10.400000  9.955000 10.570000 10.125000 ;
      RECT 10.400000 10.400000 10.570000 10.570000 ;
      RECT 10.495000  0.250000 10.665000  0.420000 ;
      RECT 10.495000  1.380000 10.665000  1.550000 ;
      RECT 10.495000 12.410000 10.665000 12.580000 ;
      RECT 10.495000 13.540000 10.665000 13.710000 ;
      RECT 10.855000  0.250000 11.025000  0.420000 ;
      RECT 10.855000  1.380000 11.025000  1.550000 ;
      RECT 10.855000 12.410000 11.025000 12.580000 ;
      RECT 10.855000 13.540000 11.025000 13.710000 ;
      RECT 11.215000  0.250000 11.385000  0.420000 ;
      RECT 11.215000  1.380000 11.385000  1.550000 ;
      RECT 11.215000 12.410000 11.385000 12.580000 ;
      RECT 11.215000 13.540000 11.385000 13.710000 ;
      RECT 11.575000  0.250000 11.745000  0.420000 ;
      RECT 11.575000  1.380000 11.745000  1.550000 ;
      RECT 11.575000 12.410000 11.745000 12.580000 ;
      RECT 11.575000 13.540000 11.745000 13.710000 ;
      RECT 11.935000  0.250000 12.105000  0.420000 ;
      RECT 11.935000  1.380000 12.105000  1.550000 ;
      RECT 11.935000 12.410000 12.105000 12.580000 ;
      RECT 11.935000 13.540000 12.105000 13.710000 ;
      RECT 12.295000  0.250000 12.465000  0.420000 ;
      RECT 12.295000 13.540000 12.465000 13.710000 ;
      RECT 12.410000  1.380000 12.580000  1.550000 ;
      RECT 12.410000  1.855000 12.580000  2.025000 ;
      RECT 12.410000  2.215000 12.580000  2.385000 ;
      RECT 12.410000  2.575000 12.580000  2.745000 ;
      RECT 12.410000  2.935000 12.580000  3.105000 ;
      RECT 12.410000  3.295000 12.580000  3.465000 ;
      RECT 12.410000  3.655000 12.580000  3.825000 ;
      RECT 12.410000  4.015000 12.580000  4.185000 ;
      RECT 12.410000  4.375000 12.580000  4.545000 ;
      RECT 12.410000  4.735000 12.580000  4.905000 ;
      RECT 12.410000  5.095000 12.580000  5.265000 ;
      RECT 12.410000  5.455000 12.580000  5.625000 ;
      RECT 12.410000  5.815000 12.580000  5.985000 ;
      RECT 12.410000  6.175000 12.580000  6.345000 ;
      RECT 12.410000  6.535000 12.580000  6.705000 ;
      RECT 12.410000  6.895000 12.580000  7.065000 ;
      RECT 12.410000  7.255000 12.580000  7.425000 ;
      RECT 12.410000  7.615000 12.580000  7.785000 ;
      RECT 12.410000  7.975000 12.580000  8.145000 ;
      RECT 12.410000  8.335000 12.580000  8.505000 ;
      RECT 12.410000  8.695000 12.580000  8.865000 ;
      RECT 12.410000  9.055000 12.580000  9.225000 ;
      RECT 12.410000  9.415000 12.580000  9.585000 ;
      RECT 12.410000  9.775000 12.580000  9.945000 ;
      RECT 12.410000 10.135000 12.580000 10.305000 ;
      RECT 12.410000 10.495000 12.580000 10.665000 ;
      RECT 12.410000 10.855000 12.580000 11.025000 ;
      RECT 12.410000 11.215000 12.580000 11.385000 ;
      RECT 12.410000 11.575000 12.580000 11.745000 ;
      RECT 12.410000 11.935000 12.580000 12.105000 ;
      RECT 12.410000 12.410000 12.580000 12.580000 ;
      RECT 12.655000  0.250000 12.825000  0.420000 ;
      RECT 12.655000 13.540000 12.825000 13.710000 ;
      RECT 13.015000  0.250000 13.185000  0.420000 ;
      RECT 13.015000 13.540000 13.185000 13.710000 ;
      RECT 13.540000  0.250000 13.710000  0.420000 ;
      RECT 13.540000  0.775000 13.710000  0.945000 ;
      RECT 13.540000  1.135000 13.710000  1.305000 ;
      RECT 13.540000  1.495000 13.710000  1.665000 ;
      RECT 13.540000  1.855000 13.710000  2.025000 ;
      RECT 13.540000  2.215000 13.710000  2.385000 ;
      RECT 13.540000  2.575000 13.710000  2.745000 ;
      RECT 13.540000  2.935000 13.710000  3.105000 ;
      RECT 13.540000  3.295000 13.710000  3.465000 ;
      RECT 13.540000  3.655000 13.710000  3.825000 ;
      RECT 13.540000  4.015000 13.710000  4.185000 ;
      RECT 13.540000  4.375000 13.710000  4.545000 ;
      RECT 13.540000  4.735000 13.710000  4.905000 ;
      RECT 13.540000  5.095000 13.710000  5.265000 ;
      RECT 13.540000  5.455000 13.710000  5.625000 ;
      RECT 13.540000  5.815000 13.710000  5.985000 ;
      RECT 13.540000  6.175000 13.710000  6.345000 ;
      RECT 13.540000  6.535000 13.710000  6.705000 ;
      RECT 13.540000  6.895000 13.710000  7.065000 ;
      RECT 13.540000  7.255000 13.710000  7.425000 ;
      RECT 13.540000  7.615000 13.710000  7.785000 ;
      RECT 13.540000  7.975000 13.710000  8.145000 ;
      RECT 13.540000  8.335000 13.710000  8.505000 ;
      RECT 13.540000  8.695000 13.710000  8.865000 ;
      RECT 13.540000  9.055000 13.710000  9.225000 ;
      RECT 13.540000  9.415000 13.710000  9.585000 ;
      RECT 13.540000  9.775000 13.710000  9.945000 ;
      RECT 13.540000 10.135000 13.710000 10.305000 ;
      RECT 13.540000 10.495000 13.710000 10.665000 ;
      RECT 13.540000 10.855000 13.710000 11.025000 ;
      RECT 13.540000 11.215000 13.710000 11.385000 ;
      RECT 13.540000 11.575000 13.710000 11.745000 ;
      RECT 13.540000 11.935000 13.710000 12.105000 ;
      RECT 13.540000 12.295000 13.710000 12.465000 ;
      RECT 13.540000 12.655000 13.710000 12.825000 ;
      RECT 13.540000 13.015000 13.710000 13.185000 ;
      RECT 13.540000 13.540000 13.710000 13.710000 ;
    LAYER met1 ;
      RECT  0.190000  0.190000 13.770000  0.480000 ;
      RECT  0.190000  0.480000  0.480000 13.480000 ;
      RECT  0.190000 13.480000 13.770000 13.770000 ;
      RECT  1.320000  1.320000 12.640000  1.610000 ;
      RECT  1.320000  1.610000  1.610000 12.350000 ;
      RECT  1.320000 12.350000 12.640000 12.640000 ;
      RECT  3.330000  3.330000 10.630000  3.620000 ;
      RECT  3.330000  3.620000  3.620000 10.340000 ;
      RECT  3.330000 10.340000 10.630000 10.630000 ;
      RECT  4.675000  4.675000  9.285000  9.285000 ;
      RECT 10.340000  3.620000 10.630000 10.340000 ;
      RECT 12.350000  1.610000 12.640000 12.350000 ;
      RECT 13.480000  0.480000 13.770000 13.480000 ;
  END
END sky130_fd_pr__rf_npn_05v5_W5p00L5p00
END LIBRARY
