module MyVerilogModule(
  input wire in_signal,
  output wire out_signal
);
  assign out_signal = in_signal;
endmodule
