MACRO PMOS_S_24460802_X3_Y12
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_24460802_X3_Y12 0 0 ;
  SIZE 4300 BY 72240 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 260 1860 65260 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 4460 2290 69460 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 680 2720 71560 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 71905 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 68545 ;
    LAYER M1 ;
      RECT 2025 68795 2275 69805 ;
    LAYER M1 ;
      RECT 2025 70895 2275 71905 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M1 ;
      RECT 2455 65015 2705 68545 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 39145 ;
    LAYER M1 ;
      RECT 2885 39395 3135 40405 ;
    LAYER M1 ;
      RECT 2885 41495 3135 45025 ;
    LAYER M1 ;
      RECT 2885 45275 3135 46285 ;
    LAYER M1 ;
      RECT 2885 47375 3135 50905 ;
    LAYER M1 ;
      RECT 2885 51155 3135 52165 ;
    LAYER M1 ;
      RECT 2885 53255 3135 56785 ;
    LAYER M1 ;
      RECT 2885 57035 3135 58045 ;
    LAYER M1 ;
      RECT 2885 59135 3135 62665 ;
    LAYER M1 ;
      RECT 2885 62915 3135 63925 ;
    LAYER M1 ;
      RECT 2885 65015 3135 68545 ;
    LAYER M1 ;
      RECT 2885 68795 3135 69805 ;
    LAYER M1 ;
      RECT 2885 70895 3135 71905 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3315 47375 3565 50905 ;
    LAYER M1 ;
      RECT 3315 53255 3565 56785 ;
    LAYER M1 ;
      RECT 3315 59135 3565 62665 ;
    LAYER M1 ;
      RECT 3315 65015 3565 68545 ;
    LAYER M2 ;
      RECT 1120 280 3180 560 ;
    LAYER M2 ;
      RECT 1120 4480 3180 4760 ;
    LAYER M2 ;
      RECT 690 700 3610 980 ;
    LAYER M2 ;
      RECT 1120 6160 3180 6440 ;
    LAYER M2 ;
      RECT 1120 10360 3180 10640 ;
    LAYER M2 ;
      RECT 690 6580 3610 6860 ;
    LAYER M2 ;
      RECT 1120 12040 3180 12320 ;
    LAYER M2 ;
      RECT 1120 16240 3180 16520 ;
    LAYER M2 ;
      RECT 690 12460 3610 12740 ;
    LAYER M2 ;
      RECT 1120 17920 3180 18200 ;
    LAYER M2 ;
      RECT 1120 22120 3180 22400 ;
    LAYER M2 ;
      RECT 690 18340 3610 18620 ;
    LAYER M2 ;
      RECT 1120 23800 3180 24080 ;
    LAYER M2 ;
      RECT 1120 28000 3180 28280 ;
    LAYER M2 ;
      RECT 690 24220 3610 24500 ;
    LAYER M2 ;
      RECT 1120 29680 3180 29960 ;
    LAYER M2 ;
      RECT 1120 33880 3180 34160 ;
    LAYER M2 ;
      RECT 690 30100 3610 30380 ;
    LAYER M2 ;
      RECT 1120 35560 3180 35840 ;
    LAYER M2 ;
      RECT 1120 39760 3180 40040 ;
    LAYER M2 ;
      RECT 690 35980 3610 36260 ;
    LAYER M2 ;
      RECT 1120 41440 3180 41720 ;
    LAYER M2 ;
      RECT 1120 45640 3180 45920 ;
    LAYER M2 ;
      RECT 690 41860 3610 42140 ;
    LAYER M2 ;
      RECT 1120 47320 3180 47600 ;
    LAYER M2 ;
      RECT 1120 51520 3180 51800 ;
    LAYER M2 ;
      RECT 690 47740 3610 48020 ;
    LAYER M2 ;
      RECT 1120 53200 3180 53480 ;
    LAYER M2 ;
      RECT 1120 57400 3180 57680 ;
    LAYER M2 ;
      RECT 690 53620 3610 53900 ;
    LAYER M2 ;
      RECT 1120 59080 3180 59360 ;
    LAYER M2 ;
      RECT 1120 63280 3180 63560 ;
    LAYER M2 ;
      RECT 690 59500 3610 59780 ;
    LAYER M2 ;
      RECT 1120 64960 3180 65240 ;
    LAYER M2 ;
      RECT 1120 69160 3180 69440 ;
    LAYER M2 ;
      RECT 1120 71260 3180 71540 ;
    LAYER M2 ;
      RECT 690 65380 3610 65660 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 35615 3095 35785 ;
    LAYER V1 ;
      RECT 2925 39815 3095 39985 ;
    LAYER V1 ;
      RECT 2925 41495 3095 41665 ;
    LAYER V1 ;
      RECT 2925 45695 3095 45865 ;
    LAYER V1 ;
      RECT 2925 47375 3095 47545 ;
    LAYER V1 ;
      RECT 2925 51575 3095 51745 ;
    LAYER V1 ;
      RECT 2925 53255 3095 53425 ;
    LAYER V1 ;
      RECT 2925 57455 3095 57625 ;
    LAYER V1 ;
      RECT 2925 59135 3095 59305 ;
    LAYER V1 ;
      RECT 2925 63335 3095 63505 ;
    LAYER V1 ;
      RECT 2925 65015 3095 65185 ;
    LAYER V1 ;
      RECT 2925 69215 3095 69385 ;
    LAYER V1 ;
      RECT 2925 71315 3095 71485 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 71315 1375 71485 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59135 2235 59305 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65015 2235 65185 ;
    LAYER V1 ;
      RECT 2065 69215 2235 69385 ;
    LAYER V1 ;
      RECT 2065 71315 2235 71485 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 41915 3525 42085 ;
    LAYER V1 ;
      RECT 3355 47795 3525 47965 ;
    LAYER V1 ;
      RECT 3355 53675 3525 53845 ;
    LAYER V1 ;
      RECT 3355 59555 3525 59725 ;
    LAYER V1 ;
      RECT 3355 65435 3525 65605 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 2495 59555 2665 59725 ;
    LAYER V1 ;
      RECT 2495 65435 2665 65605 ;
    LAYER V2 ;
      RECT 1645 345 1795 495 ;
    LAYER V2 ;
      RECT 1645 6225 1795 6375 ;
    LAYER V2 ;
      RECT 1645 12105 1795 12255 ;
    LAYER V2 ;
      RECT 1645 17985 1795 18135 ;
    LAYER V2 ;
      RECT 1645 23865 1795 24015 ;
    LAYER V2 ;
      RECT 1645 29745 1795 29895 ;
    LAYER V2 ;
      RECT 1645 35625 1795 35775 ;
    LAYER V2 ;
      RECT 1645 41505 1795 41655 ;
    LAYER V2 ;
      RECT 1645 47385 1795 47535 ;
    LAYER V2 ;
      RECT 1645 53265 1795 53415 ;
    LAYER V2 ;
      RECT 1645 59145 1795 59295 ;
    LAYER V2 ;
      RECT 1645 65025 1795 65175 ;
    LAYER V2 ;
      RECT 2075 4545 2225 4695 ;
    LAYER V2 ;
      RECT 2075 10425 2225 10575 ;
    LAYER V2 ;
      RECT 2075 16305 2225 16455 ;
    LAYER V2 ;
      RECT 2075 22185 2225 22335 ;
    LAYER V2 ;
      RECT 2075 28065 2225 28215 ;
    LAYER V2 ;
      RECT 2075 33945 2225 34095 ;
    LAYER V2 ;
      RECT 2075 39825 2225 39975 ;
    LAYER V2 ;
      RECT 2075 45705 2225 45855 ;
    LAYER V2 ;
      RECT 2075 51585 2225 51735 ;
    LAYER V2 ;
      RECT 2075 57465 2225 57615 ;
    LAYER V2 ;
      RECT 2075 63345 2225 63495 ;
    LAYER V2 ;
      RECT 2075 69225 2225 69375 ;
    LAYER V2 ;
      RECT 2505 765 2655 915 ;
    LAYER V2 ;
      RECT 2505 6645 2655 6795 ;
    LAYER V2 ;
      RECT 2505 12525 2655 12675 ;
    LAYER V2 ;
      RECT 2505 18405 2655 18555 ;
    LAYER V2 ;
      RECT 2505 24285 2655 24435 ;
    LAYER V2 ;
      RECT 2505 30165 2655 30315 ;
    LAYER V2 ;
      RECT 2505 36045 2655 36195 ;
    LAYER V2 ;
      RECT 2505 41925 2655 42075 ;
    LAYER V2 ;
      RECT 2505 47805 2655 47955 ;
    LAYER V2 ;
      RECT 2505 53685 2655 53835 ;
    LAYER V2 ;
      RECT 2505 59565 2655 59715 ;
    LAYER V2 ;
      RECT 2505 65445 2655 65595 ;
    LAYER V2 ;
      RECT 2505 71325 2655 71475 ;
  END
END PMOS_S_24460802_X3_Y12
