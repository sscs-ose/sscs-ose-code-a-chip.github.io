# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50 ;
  ORIGIN -0.050000  0.000000 ;
  SIZE  9.700000 BY  3.930000 ;
  PIN DRAIN
    ANTENNADIFFAREA  4.214000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.090000 9.750000 3.370000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  15.049999 ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.100000 8.805000 0.270000 ;
        RECT 0.995000 3.660000 8.805000 3.830000 ;
      LAYER mcon ;
        RECT 1.035000 0.100000 1.205000 0.270000 ;
        RECT 1.035000 3.660000 1.205000 3.830000 ;
        RECT 1.395000 0.100000 1.565000 0.270000 ;
        RECT 1.395000 3.660000 1.565000 3.830000 ;
        RECT 1.755000 0.100000 1.925000 0.270000 ;
        RECT 1.755000 3.660000 1.925000 3.830000 ;
        RECT 2.115000 0.100000 2.285000 0.270000 ;
        RECT 2.115000 3.660000 2.285000 3.830000 ;
        RECT 2.475000 0.100000 2.645000 0.270000 ;
        RECT 2.475000 3.660000 2.645000 3.830000 ;
        RECT 2.835000 0.100000 3.005000 0.270000 ;
        RECT 2.835000 3.660000 3.005000 3.830000 ;
        RECT 3.195000 0.100000 3.365000 0.270000 ;
        RECT 3.195000 3.660000 3.365000 3.830000 ;
        RECT 3.555000 0.100000 3.725000 0.270000 ;
        RECT 3.555000 3.660000 3.725000 3.830000 ;
        RECT 3.915000 0.100000 4.085000 0.270000 ;
        RECT 3.915000 3.660000 4.085000 3.830000 ;
        RECT 4.275000 0.100000 4.445000 0.270000 ;
        RECT 4.275000 3.660000 4.445000 3.830000 ;
        RECT 4.635000 0.100000 4.805000 0.270000 ;
        RECT 4.635000 3.660000 4.805000 3.830000 ;
        RECT 4.995000 0.100000 5.165000 0.270000 ;
        RECT 4.995000 3.660000 5.165000 3.830000 ;
        RECT 5.355000 0.100000 5.525000 0.270000 ;
        RECT 5.355000 3.660000 5.525000 3.830000 ;
        RECT 5.715000 0.100000 5.885000 0.270000 ;
        RECT 5.715000 3.660000 5.885000 3.830000 ;
        RECT 6.075000 0.100000 6.245000 0.270000 ;
        RECT 6.075000 3.660000 6.245000 3.830000 ;
        RECT 6.435000 0.100000 6.605000 0.270000 ;
        RECT 6.435000 3.660000 6.605000 3.830000 ;
        RECT 6.795000 0.100000 6.965000 0.270000 ;
        RECT 6.795000 3.660000 6.965000 3.830000 ;
        RECT 7.155000 0.100000 7.325000 0.270000 ;
        RECT 7.155000 3.660000 7.325000 3.830000 ;
        RECT 7.515000 0.100000 7.685000 0.270000 ;
        RECT 7.515000 3.660000 7.685000 3.830000 ;
        RECT 7.875000 0.100000 8.045000 0.270000 ;
        RECT 7.875000 3.660000 8.045000 3.830000 ;
        RECT 8.235000 0.100000 8.405000 0.270000 ;
        RECT 8.235000 3.660000 8.405000 3.830000 ;
        RECT 8.595000 0.100000 8.765000 0.270000 ;
        RECT 8.595000 3.660000 8.765000 3.830000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.975000 0.000000 8.825000 0.330000 ;
        RECT 0.975000 3.600000 8.825000 3.930000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  5.056800 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.560000 9.750000 1.840000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.872900 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.560000 0.470000 3.370000 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.330000 0.560000 9.620000 3.370000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.610000 0.410000 3.320000 ;
      RECT 0.915000 0.440000 1.085000 3.490000 ;
      RECT 1.695000 0.440000 1.865000 3.490000 ;
      RECT 2.475000 0.440000 2.645000 3.490000 ;
      RECT 3.255000 0.440000 3.425000 3.490000 ;
      RECT 4.035000 0.440000 4.205000 3.490000 ;
      RECT 4.815000 0.440000 4.985000 3.490000 ;
      RECT 5.595000 0.440000 5.765000 3.490000 ;
      RECT 6.375000 0.440000 6.545000 3.490000 ;
      RECT 7.155000 0.440000 7.325000 3.490000 ;
      RECT 7.935000 0.440000 8.105000 3.490000 ;
      RECT 8.715000 0.440000 8.885000 3.490000 ;
      RECT 9.390000 0.610000 9.560000 3.320000 ;
    LAYER mcon ;
      RECT 0.240000 0.620000 0.410000 0.790000 ;
      RECT 0.240000 0.980000 0.410000 1.150000 ;
      RECT 0.240000 1.340000 0.410000 1.510000 ;
      RECT 0.240000 1.700000 0.410000 1.870000 ;
      RECT 0.240000 2.060000 0.410000 2.230000 ;
      RECT 0.240000 2.420000 0.410000 2.590000 ;
      RECT 0.240000 2.780000 0.410000 2.950000 ;
      RECT 0.240000 3.140000 0.410000 3.310000 ;
      RECT 0.915000 0.620000 1.085000 0.790000 ;
      RECT 0.915000 0.980000 1.085000 1.150000 ;
      RECT 0.915000 1.340000 1.085000 1.510000 ;
      RECT 0.915000 1.700000 1.085000 1.870000 ;
      RECT 0.915000 2.060000 1.085000 2.230000 ;
      RECT 0.915000 2.420000 1.085000 2.590000 ;
      RECT 0.915000 2.780000 1.085000 2.950000 ;
      RECT 0.915000 3.140000 1.085000 3.310000 ;
      RECT 1.695000 0.620000 1.865000 0.790000 ;
      RECT 1.695000 0.980000 1.865000 1.150000 ;
      RECT 1.695000 1.340000 1.865000 1.510000 ;
      RECT 1.695000 1.700000 1.865000 1.870000 ;
      RECT 1.695000 2.060000 1.865000 2.230000 ;
      RECT 1.695000 2.420000 1.865000 2.590000 ;
      RECT 1.695000 2.780000 1.865000 2.950000 ;
      RECT 1.695000 3.140000 1.865000 3.310000 ;
      RECT 2.475000 0.620000 2.645000 0.790000 ;
      RECT 2.475000 0.980000 2.645000 1.150000 ;
      RECT 2.475000 1.340000 2.645000 1.510000 ;
      RECT 2.475000 1.700000 2.645000 1.870000 ;
      RECT 2.475000 2.060000 2.645000 2.230000 ;
      RECT 2.475000 2.420000 2.645000 2.590000 ;
      RECT 2.475000 2.780000 2.645000 2.950000 ;
      RECT 2.475000 3.140000 2.645000 3.310000 ;
      RECT 3.255000 0.620000 3.425000 0.790000 ;
      RECT 3.255000 0.980000 3.425000 1.150000 ;
      RECT 3.255000 1.340000 3.425000 1.510000 ;
      RECT 3.255000 1.700000 3.425000 1.870000 ;
      RECT 3.255000 2.060000 3.425000 2.230000 ;
      RECT 3.255000 2.420000 3.425000 2.590000 ;
      RECT 3.255000 2.780000 3.425000 2.950000 ;
      RECT 3.255000 3.140000 3.425000 3.310000 ;
      RECT 4.035000 0.620000 4.205000 0.790000 ;
      RECT 4.035000 0.980000 4.205000 1.150000 ;
      RECT 4.035000 1.340000 4.205000 1.510000 ;
      RECT 4.035000 1.700000 4.205000 1.870000 ;
      RECT 4.035000 2.060000 4.205000 2.230000 ;
      RECT 4.035000 2.420000 4.205000 2.590000 ;
      RECT 4.035000 2.780000 4.205000 2.950000 ;
      RECT 4.035000 3.140000 4.205000 3.310000 ;
      RECT 4.815000 0.620000 4.985000 0.790000 ;
      RECT 4.815000 0.980000 4.985000 1.150000 ;
      RECT 4.815000 1.340000 4.985000 1.510000 ;
      RECT 4.815000 1.700000 4.985000 1.870000 ;
      RECT 4.815000 2.060000 4.985000 2.230000 ;
      RECT 4.815000 2.420000 4.985000 2.590000 ;
      RECT 4.815000 2.780000 4.985000 2.950000 ;
      RECT 4.815000 3.140000 4.985000 3.310000 ;
      RECT 5.595000 0.620000 5.765000 0.790000 ;
      RECT 5.595000 0.980000 5.765000 1.150000 ;
      RECT 5.595000 1.340000 5.765000 1.510000 ;
      RECT 5.595000 1.700000 5.765000 1.870000 ;
      RECT 5.595000 2.060000 5.765000 2.230000 ;
      RECT 5.595000 2.420000 5.765000 2.590000 ;
      RECT 5.595000 2.780000 5.765000 2.950000 ;
      RECT 5.595000 3.140000 5.765000 3.310000 ;
      RECT 6.375000 0.620000 6.545000 0.790000 ;
      RECT 6.375000 0.980000 6.545000 1.150000 ;
      RECT 6.375000 1.340000 6.545000 1.510000 ;
      RECT 6.375000 1.700000 6.545000 1.870000 ;
      RECT 6.375000 2.060000 6.545000 2.230000 ;
      RECT 6.375000 2.420000 6.545000 2.590000 ;
      RECT 6.375000 2.780000 6.545000 2.950000 ;
      RECT 6.375000 3.140000 6.545000 3.310000 ;
      RECT 7.155000 0.620000 7.325000 0.790000 ;
      RECT 7.155000 0.980000 7.325000 1.150000 ;
      RECT 7.155000 1.340000 7.325000 1.510000 ;
      RECT 7.155000 1.700000 7.325000 1.870000 ;
      RECT 7.155000 2.060000 7.325000 2.230000 ;
      RECT 7.155000 2.420000 7.325000 2.590000 ;
      RECT 7.155000 2.780000 7.325000 2.950000 ;
      RECT 7.155000 3.140000 7.325000 3.310000 ;
      RECT 7.935000 0.620000 8.105000 0.790000 ;
      RECT 7.935000 0.980000 8.105000 1.150000 ;
      RECT 7.935000 1.340000 8.105000 1.510000 ;
      RECT 7.935000 1.700000 8.105000 1.870000 ;
      RECT 7.935000 2.060000 8.105000 2.230000 ;
      RECT 7.935000 2.420000 8.105000 2.590000 ;
      RECT 7.935000 2.780000 8.105000 2.950000 ;
      RECT 7.935000 3.140000 8.105000 3.310000 ;
      RECT 8.715000 0.620000 8.885000 0.790000 ;
      RECT 8.715000 0.980000 8.885000 1.150000 ;
      RECT 8.715000 1.340000 8.885000 1.510000 ;
      RECT 8.715000 1.700000 8.885000 1.870000 ;
      RECT 8.715000 2.060000 8.885000 2.230000 ;
      RECT 8.715000 2.420000 8.885000 2.590000 ;
      RECT 8.715000 2.780000 8.885000 2.950000 ;
      RECT 8.715000 3.140000 8.885000 3.310000 ;
      RECT 9.390000 0.620000 9.560000 0.790000 ;
      RECT 9.390000 0.980000 9.560000 1.150000 ;
      RECT 9.390000 1.340000 9.560000 1.510000 ;
      RECT 9.390000 1.700000 9.560000 1.870000 ;
      RECT 9.390000 2.060000 9.560000 2.230000 ;
      RECT 9.390000 2.420000 9.560000 2.590000 ;
      RECT 9.390000 2.780000 9.560000 2.950000 ;
      RECT 9.390000 3.140000 9.560000 3.310000 ;
    LAYER met1 ;
      RECT 0.870000 0.560000 1.130000 3.370000 ;
      RECT 1.650000 0.560000 1.910000 3.370000 ;
      RECT 2.430000 0.560000 2.690000 3.370000 ;
      RECT 3.210000 0.560000 3.470000 3.370000 ;
      RECT 3.990000 0.560000 4.250000 3.370000 ;
      RECT 4.770000 0.560000 5.030000 3.370000 ;
      RECT 5.550000 0.560000 5.810000 3.370000 ;
      RECT 6.330000 0.560000 6.590000 3.370000 ;
      RECT 7.110000 0.560000 7.370000 3.370000 ;
      RECT 7.890000 0.560000 8.150000 3.370000 ;
      RECT 8.670000 0.560000 8.930000 3.370000 ;
    LAYER via ;
      RECT 0.870000 0.590000 1.130000 0.850000 ;
      RECT 0.870000 0.910000 1.130000 1.170000 ;
      RECT 0.870000 1.230000 1.130000 1.490000 ;
      RECT 0.870000 1.550000 1.130000 1.810000 ;
      RECT 1.650000 2.120000 1.910000 2.380000 ;
      RECT 1.650000 2.440000 1.910000 2.700000 ;
      RECT 1.650000 2.760000 1.910000 3.020000 ;
      RECT 1.650000 3.080000 1.910000 3.340000 ;
      RECT 2.430000 0.590000 2.690000 0.850000 ;
      RECT 2.430000 0.910000 2.690000 1.170000 ;
      RECT 2.430000 1.230000 2.690000 1.490000 ;
      RECT 2.430000 1.550000 2.690000 1.810000 ;
      RECT 3.210000 2.120000 3.470000 2.380000 ;
      RECT 3.210000 2.440000 3.470000 2.700000 ;
      RECT 3.210000 2.760000 3.470000 3.020000 ;
      RECT 3.210000 3.080000 3.470000 3.340000 ;
      RECT 3.990000 0.590000 4.250000 0.850000 ;
      RECT 3.990000 0.910000 4.250000 1.170000 ;
      RECT 3.990000 1.230000 4.250000 1.490000 ;
      RECT 3.990000 1.550000 4.250000 1.810000 ;
      RECT 4.770000 2.120000 5.030000 2.380000 ;
      RECT 4.770000 2.440000 5.030000 2.700000 ;
      RECT 4.770000 2.760000 5.030000 3.020000 ;
      RECT 4.770000 3.080000 5.030000 3.340000 ;
      RECT 5.550000 0.590000 5.810000 0.850000 ;
      RECT 5.550000 0.910000 5.810000 1.170000 ;
      RECT 5.550000 1.230000 5.810000 1.490000 ;
      RECT 5.550000 1.550000 5.810000 1.810000 ;
      RECT 6.330000 2.120000 6.590000 2.380000 ;
      RECT 6.330000 2.440000 6.590000 2.700000 ;
      RECT 6.330000 2.760000 6.590000 3.020000 ;
      RECT 6.330000 3.080000 6.590000 3.340000 ;
      RECT 7.110000 0.590000 7.370000 0.850000 ;
      RECT 7.110000 0.910000 7.370000 1.170000 ;
      RECT 7.110000 1.230000 7.370000 1.490000 ;
      RECT 7.110000 1.550000 7.370000 1.810000 ;
      RECT 7.890000 2.120000 8.150000 2.380000 ;
      RECT 7.890000 2.440000 8.150000 2.700000 ;
      RECT 7.890000 2.760000 8.150000 3.020000 ;
      RECT 7.890000 3.080000 8.150000 3.340000 ;
      RECT 8.670000 0.590000 8.930000 0.850000 ;
      RECT 8.670000 0.910000 8.930000 1.170000 ;
      RECT 8.670000 1.230000 8.930000 1.490000 ;
      RECT 8.670000 1.550000 8.930000 1.810000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50
END LIBRARY
