# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15 ;
  ORIGIN  0.000000  0.485000 ;
  SIZE  2.330000 BY  6.160000 ;
  PIN DRAIN
    ANTENNADIFFAREA  2.800000 ;
    PORT
      LAYER met3 ;
        RECT 0.570000 4.375000 0.900000 4.815000 ;
        RECT 0.570000 4.815000 1.760000 5.145000 ;
        RECT 1.430000 4.375000 1.760000 4.815000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.000000 ;
    PORT
      LAYER met1 ;
        RECT 0.480000 5.365000 1.850000 5.655000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.050000 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.485000 2.140000 -0.225000 ;
        RECT 0.190000 -0.225000 0.420000  5.105000 ;
        RECT 1.050000 -0.225000 1.280000  5.105000 ;
        RECT 1.910000 -0.225000 2.140000  5.105000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.255000 0.390000 5.105000 ;
      RECT 0.490000 5.335000 1.840000 5.675000 ;
      RECT 0.650000 0.255000 0.820000 5.105000 ;
      RECT 1.080000 0.255000 1.250000 5.105000 ;
      RECT 1.510000 0.255000 1.680000 5.105000 ;
      RECT 1.940000 0.255000 2.110000 5.105000 ;
    LAYER mcon ;
      RECT 0.220000 0.425000 0.390000 0.595000 ;
      RECT 0.220000 0.785000 0.390000 0.955000 ;
      RECT 0.220000 1.145000 0.390000 1.315000 ;
      RECT 0.220000 1.505000 0.390000 1.675000 ;
      RECT 0.220000 1.865000 0.390000 2.035000 ;
      RECT 0.220000 2.225000 0.390000 2.395000 ;
      RECT 0.220000 2.585000 0.390000 2.755000 ;
      RECT 0.220000 2.945000 0.390000 3.115000 ;
      RECT 0.220000 3.305000 0.390000 3.475000 ;
      RECT 0.220000 3.665000 0.390000 3.835000 ;
      RECT 0.220000 4.025000 0.390000 4.195000 ;
      RECT 0.220000 4.385000 0.390000 4.555000 ;
      RECT 0.220000 4.745000 0.390000 4.915000 ;
      RECT 0.540000 5.425000 0.710000 5.595000 ;
      RECT 0.650000 0.425000 0.820000 0.595000 ;
      RECT 0.650000 0.785000 0.820000 0.955000 ;
      RECT 0.650000 1.145000 0.820000 1.315000 ;
      RECT 0.650000 1.505000 0.820000 1.675000 ;
      RECT 0.650000 1.865000 0.820000 2.035000 ;
      RECT 0.650000 2.225000 0.820000 2.395000 ;
      RECT 0.650000 2.585000 0.820000 2.755000 ;
      RECT 0.650000 2.945000 0.820000 3.115000 ;
      RECT 0.650000 3.305000 0.820000 3.475000 ;
      RECT 0.650000 3.665000 0.820000 3.835000 ;
      RECT 0.650000 4.025000 0.820000 4.195000 ;
      RECT 0.650000 4.385000 0.820000 4.555000 ;
      RECT 0.650000 4.745000 0.820000 4.915000 ;
      RECT 0.900000 5.425000 1.070000 5.595000 ;
      RECT 1.080000 0.425000 1.250000 0.595000 ;
      RECT 1.080000 0.785000 1.250000 0.955000 ;
      RECT 1.080000 1.145000 1.250000 1.315000 ;
      RECT 1.080000 1.505000 1.250000 1.675000 ;
      RECT 1.080000 1.865000 1.250000 2.035000 ;
      RECT 1.080000 2.225000 1.250000 2.395000 ;
      RECT 1.080000 2.585000 1.250000 2.755000 ;
      RECT 1.080000 2.945000 1.250000 3.115000 ;
      RECT 1.080000 3.305000 1.250000 3.475000 ;
      RECT 1.080000 3.665000 1.250000 3.835000 ;
      RECT 1.080000 4.025000 1.250000 4.195000 ;
      RECT 1.080000 4.385000 1.250000 4.555000 ;
      RECT 1.080000 4.745000 1.250000 4.915000 ;
      RECT 1.260000 5.425000 1.430000 5.595000 ;
      RECT 1.510000 0.425000 1.680000 0.595000 ;
      RECT 1.510000 0.785000 1.680000 0.955000 ;
      RECT 1.510000 1.145000 1.680000 1.315000 ;
      RECT 1.510000 1.505000 1.680000 1.675000 ;
      RECT 1.510000 1.865000 1.680000 2.035000 ;
      RECT 1.510000 2.225000 1.680000 2.395000 ;
      RECT 1.510000 2.585000 1.680000 2.755000 ;
      RECT 1.510000 2.945000 1.680000 3.115000 ;
      RECT 1.510000 3.305000 1.680000 3.475000 ;
      RECT 1.510000 3.665000 1.680000 3.835000 ;
      RECT 1.510000 4.025000 1.680000 4.195000 ;
      RECT 1.510000 4.385000 1.680000 4.555000 ;
      RECT 1.510000 4.745000 1.680000 4.915000 ;
      RECT 1.620000 5.425000 1.790000 5.595000 ;
      RECT 1.940000 0.425000 2.110000 0.595000 ;
      RECT 1.940000 0.785000 2.110000 0.955000 ;
      RECT 1.940000 1.145000 2.110000 1.315000 ;
      RECT 1.940000 1.505000 2.110000 1.675000 ;
      RECT 1.940000 1.865000 2.110000 2.035000 ;
      RECT 1.940000 2.225000 2.110000 2.395000 ;
      RECT 1.940000 2.585000 2.110000 2.755000 ;
      RECT 1.940000 2.945000 2.110000 3.115000 ;
      RECT 1.940000 3.305000 2.110000 3.475000 ;
      RECT 1.940000 3.665000 2.110000 3.835000 ;
      RECT 1.940000 4.025000 2.110000 4.195000 ;
      RECT 1.940000 4.385000 2.110000 4.555000 ;
      RECT 1.940000 4.745000 2.110000 4.915000 ;
    LAYER met1 ;
      RECT 0.605000 0.255000 0.865000 5.105000 ;
      RECT 1.465000 0.255000 1.725000 5.105000 ;
    LAYER met2 ;
      RECT 0.570000 4.375000 0.900000 5.145000 ;
      RECT 1.430000 4.375000 1.760000 5.145000 ;
    LAYER via ;
      RECT 0.605000 4.470000 0.865000 4.730000 ;
      RECT 0.605000 4.790000 0.865000 5.050000 ;
      RECT 1.465000 4.470000 1.725000 4.730000 ;
      RECT 1.465000 4.790000 1.725000 5.050000 ;
    LAYER via2 ;
      RECT 0.595000 4.420000 0.875000 4.700000 ;
      RECT 0.595000 4.820000 0.875000 5.100000 ;
      RECT 1.455000 4.420000 1.735000 4.700000 ;
      RECT 1.455000 4.820000 1.735000 5.100000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15
END LIBRARY
