MACRO SCM_PMOS_85912433_X1_Y5
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_PMOS_85912433_X1_Y5 0 0 ;
  SIZE 5160 BY 31080 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 260 2290 28300 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 680 2720 24520 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 1100 3150 30400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 4115 1845 5125 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 9995 1845 11005 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 15875 1845 16885 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 21755 1845 22765 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 27635 1845 28645 ;
    LAYER M1 ;
      RECT 1595 29735 1845 30745 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 4115 3565 5125 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 9995 3565 11005 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 15875 3565 16885 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 21755 3565 22765 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 27635 3565 28645 ;
    LAYER M1 ;
      RECT 3315 29735 3565 30745 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 1550 4480 3610 4760 ;
    LAYER M2 ;
      RECT 2410 700 3610 980 ;
    LAYER M2 ;
      RECT 690 1120 4470 1400 ;
    LAYER M2 ;
      RECT 1980 6160 3610 6440 ;
    LAYER M2 ;
      RECT 1550 10360 3610 10640 ;
    LAYER M2 ;
      RECT 1550 6580 2750 6860 ;
    LAYER M2 ;
      RECT 690 7000 4470 7280 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 1550 16240 3610 16520 ;
    LAYER M2 ;
      RECT 2410 12460 3610 12740 ;
    LAYER M2 ;
      RECT 690 12880 4470 13160 ;
    LAYER M2 ;
      RECT 1980 17920 3610 18200 ;
    LAYER M2 ;
      RECT 1550 22120 3610 22400 ;
    LAYER M2 ;
      RECT 1550 18340 2750 18620 ;
    LAYER M2 ;
      RECT 690 18760 4470 19040 ;
    LAYER M2 ;
      RECT 1120 23800 2320 24080 ;
    LAYER M2 ;
      RECT 1550 28000 3610 28280 ;
    LAYER M2 ;
      RECT 2410 24220 3610 24500 ;
    LAYER M2 ;
      RECT 690 24640 4470 24920 ;
    LAYER M2 ;
      RECT 1550 30100 3610 30380 ;
    LAYER V1 ;
      RECT 1635 335 1805 505 ;
    LAYER V1 ;
      RECT 1635 4535 1805 4705 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 10415 1805 10585 ;
    LAYER V1 ;
      RECT 1635 12095 1805 12265 ;
    LAYER V1 ;
      RECT 1635 16295 1805 16465 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 22175 1805 22345 ;
    LAYER V1 ;
      RECT 1635 23855 1805 24025 ;
    LAYER V1 ;
      RECT 1635 28055 1805 28225 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 4535 3525 4705 ;
    LAYER V1 ;
      RECT 3355 6215 3525 6385 ;
    LAYER V1 ;
      RECT 3355 10415 3525 10585 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 16295 3525 16465 ;
    LAYER V1 ;
      RECT 3355 17975 3525 18145 ;
    LAYER V1 ;
      RECT 3355 22175 3525 22345 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 28055 3525 28225 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 775 7055 945 7225 ;
    LAYER V1 ;
      RECT 775 12935 945 13105 ;
    LAYER V1 ;
      RECT 775 18815 945 18985 ;
    LAYER V1 ;
      RECT 775 24695 945 24865 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 4215 7055 4385 7225 ;
    LAYER V1 ;
      RECT 4215 12935 4385 13105 ;
    LAYER V1 ;
      RECT 4215 18815 4385 18985 ;
    LAYER V1 ;
      RECT 4215 24695 4385 24865 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 2495 7055 2665 7225 ;
    LAYER V1 ;
      RECT 2495 12935 2665 13105 ;
    LAYER V1 ;
      RECT 2495 18815 2665 18985 ;
    LAYER V1 ;
      RECT 2495 24695 2665 24865 ;
    LAYER V2 ;
      RECT 2075 345 2225 495 ;
    LAYER V2 ;
      RECT 2075 4545 2225 4695 ;
    LAYER V2 ;
      RECT 2075 6225 2225 6375 ;
    LAYER V2 ;
      RECT 2075 10425 2225 10575 ;
    LAYER V2 ;
      RECT 2075 12105 2225 12255 ;
    LAYER V2 ;
      RECT 2075 16305 2225 16455 ;
    LAYER V2 ;
      RECT 2075 17985 2225 18135 ;
    LAYER V2 ;
      RECT 2075 22185 2225 22335 ;
    LAYER V2 ;
      RECT 2075 23865 2225 24015 ;
    LAYER V2 ;
      RECT 2075 28065 2225 28215 ;
    LAYER V2 ;
      RECT 2505 765 2655 915 ;
    LAYER V2 ;
      RECT 2505 6645 2655 6795 ;
    LAYER V2 ;
      RECT 2505 12525 2655 12675 ;
    LAYER V2 ;
      RECT 2505 18405 2655 18555 ;
    LAYER V2 ;
      RECT 2505 24285 2655 24435 ;
    LAYER V2 ;
      RECT 2935 1185 3085 1335 ;
    LAYER V2 ;
      RECT 2935 7065 3085 7215 ;
    LAYER V2 ;
      RECT 2935 12945 3085 13095 ;
    LAYER V2 ;
      RECT 2935 18825 3085 18975 ;
    LAYER V2 ;
      RECT 2935 24705 3085 24855 ;
    LAYER V2 ;
      RECT 2935 30165 3085 30315 ;
  END
END SCM_PMOS_85912433_X1_Y5
