magic
tech sky130A
magscale 1 2
timestamp 1762091453
<< locali >>
rect -4052 119728 -88 119742
rect -4052 118536 5082 119728
rect -4052 118144 -88 118536
rect -4024 7782 -106 118144
rect -4046 7200 -106 7782
rect 634 46536 5080 118536
rect 634 46140 5050 46536
rect -1366 3778 -884 3782
rect -1366 3722 -1252 3778
rect -972 3722 -884 3778
rect -1366 3720 -884 3722
rect -3288 1740 -2674 1876
rect -3288 -2712 -3128 1740
rect -2818 -2542 -2674 1740
rect 634 -1048 1500 46140
rect 1784 6980 5050 46140
rect 1784 6860 5064 6980
rect 634 -2090 854 -1048
rect 1256 -2090 1472 -1048
rect 634 -2104 1472 -2090
rect 1784 -2104 2174 6860
rect 156 -2158 506 -2142
rect 156 -2168 242 -2158
rect 156 -2202 192 -2168
rect 156 -2214 242 -2202
rect 418 -2168 506 -2158
rect 480 -2202 506 -2168
rect 418 -2214 506 -2202
rect 156 -2220 506 -2214
rect 634 -2150 2174 -2104
rect 2630 -2150 5064 6860
rect -658 -2542 -112 -2246
rect 634 -2470 5064 -2150
rect 634 -2542 2660 -2470
rect -2818 -2662 4540 -2542
rect -3282 -2994 -3128 -2712
rect 4380 -2994 4540 -2662
rect -3282 -3112 4540 -2994
<< viali >>
rect -1252 3722 -972 3778
rect -3128 -2662 -2818 1740
rect 242 -2214 418 -2158
rect -3128 -2994 4380 -2662
<< metal1 >>
rect -1846 20202 -1554 21016
rect -3202 17330 -3192 17652
rect -2902 17330 -2892 17652
rect 350 17346 360 17648
rect 416 17346 426 17648
rect -3192 16690 -2898 17330
rect -2470 16746 -2190 16752
rect -3190 15490 -2906 16690
rect -2470 16380 -2460 16746
rect -2200 16380 -2190 16746
rect 1654 16382 1664 16756
rect 1728 16382 1738 16756
rect -2470 15510 -2190 16380
rect -1012 6812 -282 7046
rect 2240 7022 3014 7028
rect -3076 6200 -2976 6708
rect -2388 6424 -2302 6766
rect -2388 6423 -1872 6424
rect -1779 6423 -1685 6797
rect -2388 6329 -1685 6423
rect 2240 6358 3976 7022
rect 2754 6354 3976 6358
rect -2388 6322 -1872 6329
rect -2254 6200 -2156 6202
rect -3076 6110 -2156 6200
rect -4038 6038 -3854 6050
rect -3200 6038 -3098 6040
rect -4038 6036 -3098 6038
rect -4060 5966 -3098 6036
rect -4060 1178 -3854 5966
rect -3200 5756 -3098 5966
rect -2254 5886 -2156 6110
rect -1980 5866 -1886 6322
rect -1286 3988 -1276 4270
rect -1220 3988 -1210 4270
rect -1692 3852 -1374 3876
rect -1692 3820 -1028 3852
rect -1692 3732 -1374 3820
rect -1264 3778 -960 3784
rect -1264 3722 -1252 3778
rect -972 3746 -960 3778
rect -972 3722 -900 3746
rect -1264 3716 -900 3722
rect -1246 3034 -900 3716
rect -1246 2900 -1236 3034
rect -1098 2900 -900 3034
rect -3134 1744 -2812 1752
rect -4038 -2114 -3854 1178
rect -4058 -2124 -3854 -2114
rect -3486 1740 -2672 1744
rect -4058 -3708 -3860 -2124
rect -3486 -2994 -3128 1740
rect -2818 -2594 -2672 1740
rect -1246 -2594 -900 2900
rect 3312 -1256 3960 6354
rect 218 -1650 268 -1638
rect 218 -2000 294 -1650
rect 1148 -1852 1372 -1790
rect 218 -2152 268 -2000
rect 984 -2058 1104 -1988
rect 1326 -1990 1372 -1852
rect 1534 -1906 1544 -1600
rect 1606 -1906 1616 -1600
rect 1326 -2006 1670 -1990
rect 3280 -1992 6426 -1256
rect 1326 -2050 2400 -2006
rect 1326 -2054 1372 -2050
rect 298 -2112 1104 -2058
rect 298 -2118 362 -2112
rect 984 -2118 1104 -2112
rect 218 -2158 430 -2152
rect 218 -2166 242 -2158
rect 418 -2166 430 -2158
rect 214 -2226 224 -2166
rect 426 -2226 436 -2166
rect -2818 -2606 5140 -2594
rect -2818 -2662 1486 -2606
rect 1606 -2662 5140 -2606
rect 4380 -2994 5140 -2662
rect -3486 -3258 5140 -2994
rect -2672 -3268 5140 -3258
rect 4448 -3696 5404 -3688
rect 5798 -3696 6426 -1992
rect 4448 -3708 6426 -3696
rect -4058 -3822 144 -3708
rect 508 -3710 6426 -3708
rect 510 -3758 6426 -3710
rect 510 -3822 6356 -3758
rect -4058 -4298 6356 -3822
rect -4058 -4306 -3860 -4298
rect 4448 -4338 6356 -4298
rect 5262 -4358 6356 -4338
<< via1 >>
rect -3192 17330 -2902 17652
rect 360 17346 416 17648
rect -2460 16380 -2200 16746
rect 1664 16382 1728 16756
rect -1276 3988 -1220 4270
rect -1236 2900 -1098 3034
rect 1544 -1906 1606 -1600
rect 224 -2214 242 -2166
rect 242 -2214 418 -2166
rect 418 -2214 426 -2166
rect 224 -2226 426 -2214
rect 1486 -2662 1606 -2606
rect 1486 -2740 1606 -2662
rect 144 -3822 510 -3710
<< metal2 >>
rect -3192 17654 -2902 17662
rect 360 17654 416 17658
rect -3234 17652 416 17654
rect -3234 17330 -3192 17652
rect -2902 17648 416 17652
rect -2902 17346 360 17648
rect -2902 17330 416 17346
rect -3234 17328 416 17330
rect -3192 17320 -2902 17328
rect 1664 16762 1728 16766
rect -2460 16756 1732 16762
rect -2460 16746 1664 16756
rect -2200 16382 1664 16746
rect 1728 16382 1732 16756
rect -2200 16380 1732 16382
rect -2460 16378 1732 16380
rect -2460 16370 -2200 16378
rect 1664 16372 1728 16378
rect -1296 4270 -1218 4280
rect -1296 3988 -1276 4270
rect -1220 3988 -1218 4270
rect -1296 3722 -1218 3988
rect -1296 3718 -1216 3722
rect -1294 3044 -1216 3718
rect -1294 3034 -1098 3044
rect -1294 2902 -1236 3034
rect -1236 2890 -1098 2900
rect 1544 -1594 1606 -1590
rect 1486 -1600 1606 -1594
rect 1486 -1906 1544 -1600
rect 1486 -1916 1606 -1906
rect 224 -2162 426 -2156
rect 202 -2166 438 -2162
rect 202 -2226 224 -2166
rect 426 -2226 438 -2166
rect 202 -3700 438 -2226
rect 1486 -2596 1604 -1916
rect 1486 -2606 1606 -2596
rect 1486 -2750 1606 -2740
rect 144 -3710 510 -3700
rect 144 -3832 510 -3822
use integration  integration_0 sky130-opamp/integration/mag
timestamp 1729420727
transform 1 0 -3826 0 1 3213
box 0 -1397 2410 2687
use sky130_fd_pr__nfet_01v8_DVKA3G  XM1
timestamp 1762084523
transform 1 0 1050 0 1 -1581
box -276 -579 276 579
use sky130_fd_pr__nfet_01v8_FAV24X  XM4
timestamp 1762084523
transform 1 0 1633 0 1 22011
box -211 -24179 211 24179
use sky130_fd_pr__pfet_01v8_U7EAHW  XM5
timestamp 1762087944
transform -1 0 331 0 -1 57946
box -211 -60184 211 60184
use sky130_fd_pr__nfet_01v8_G4U28Y  XM13
timestamp 1762072077
transform 1 0 -1126 0 -1 5461
box -276 -1779 276 1779
use sky130_fd_pr__res_high_po_1p41_8KNH8U  XR1
timestamp 1762072077
transform 1 0 -3041 0 1 11288
box -307 -4782 307 4782
use sky130_fd_pr__res_high_po_1p41_8KNH8U  XR3
timestamp 1762072077
transform 1 0 -385 0 1 2474
box -307 -4782 307 4782
use sky130_fd_pr__res_high_po_1p41_6QW2RV  XR4
timestamp 1762072077
transform 1 0 -1703 0 1 13498
box -307 -6982 307 6982
use sky130_fd_pr__res_high_po_1p41_8KNH8U  XR5
timestamp 1762072077
transform 1 0 -2339 0 1 11292
box -307 -4782 307 4782
use sky130_fd_pr__res_high_po_1p41_QAVZGT  XR7
timestamp 1762072077
transform 1 0 2383 0 1 2370
box -307 -4582 307 4582
<< labels >>
flabel metal1 1160 -4254 1796 -3904 0 FreeSans 1600 0 0 0 VCC
port 5 nsew
flabel metal1 -3158 16240 -2948 16544 0 FreeSans 1600 0 0 0 CAN+
port 3 nsew
flabel metal1 -2458 16228 -2220 16522 0 FreeSans 1600 0 0 0 CAN-
port 4 nsew
flabel metal1 -1824 20584 -1568 20862 0 FreeSans 1600 0 0 0 RX
port 7 nsew
flabel metal1 572 -2112 754 -2064 0 FreeSans 1600 0 0 0 TX
port 8 nsew
flabel locali 1156 -3040 1792 -2690 0 FreeSans 1600 0 0 0 GND
port 6 nsew
<< end >>
