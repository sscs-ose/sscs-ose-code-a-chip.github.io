* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p18 BULK DRAIN GATE SOURCE
X0 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 w=1.65e+06u l=180000u
X1 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 w=1.65e+06u l=180000u
X2 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 w=1.65e+06u l=180000u
X3 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 w=1.65e+06u l=180000u
.ends
