# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.580000 BY  7.840000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT 0.000000 0.000000 8.580000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 7.510000 ;
        RECT 0.000000 7.510000 8.580000 7.840000 ;
        RECT 1.320000 0.330000 1.710000 3.455000 ;
        RECT 1.320000 4.385000 1.710000 7.510000 ;
        RECT 2.700000 0.330000 3.090000 3.455000 ;
        RECT 2.700000 4.385000 3.090000 7.510000 ;
        RECT 4.095000 0.330000 4.485000 3.455000 ;
        RECT 4.095000 4.385000 4.485000 7.510000 ;
        RECT 5.490000 0.330000 5.880000 3.455000 ;
        RECT 5.490000 4.385000 5.880000 7.510000 ;
        RECT 6.870000 0.330000 7.260000 3.455000 ;
        RECT 6.870000 4.385000 7.260000 7.510000 ;
        RECT 8.250000 0.330000 8.580000 7.510000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT 0.630000 0.630000 1.020000 3.755000 ;
        RECT 0.630000 3.755000 7.950000 4.085000 ;
        RECT 0.630000 4.085000 1.020000 7.210000 ;
        RECT 2.010000 0.630000 2.400000 3.755000 ;
        RECT 2.010000 4.085000 2.400000 7.210000 ;
        RECT 3.390000 0.630000 3.780000 3.755000 ;
        RECT 3.390000 4.085000 3.780000 7.210000 ;
        RECT 4.800000 0.630000 5.190000 3.755000 ;
        RECT 4.800000 4.085000 5.190000 7.210000 ;
        RECT 6.180000 0.630000 6.570000 3.755000 ;
        RECT 6.180000 4.085000 6.570000 7.210000 ;
        RECT 7.560000 0.630000 7.950000 3.755000 ;
        RECT 7.560000 4.085000 7.950000 7.210000 ;
    END
  END C1
  PIN MET5
    PORT
      LAYER met5 ;
        RECT 0.000000 0.000000 8.580000 7.840000 ;
    END
  END MET5
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 4.470000 4.105000 4.590000 4.360000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 8.580000 7.840000 ;
    LAYER mcon ;
      RECT 0.080000 0.415000 0.250000 0.585000 ;
      RECT 0.080000 0.775000 0.250000 0.945000 ;
      RECT 0.080000 1.135000 0.250000 1.305000 ;
      RECT 0.080000 1.495000 0.250000 1.665000 ;
      RECT 0.080000 1.855000 0.250000 2.025000 ;
      RECT 0.080000 2.215000 0.250000 2.385000 ;
      RECT 0.080000 2.575000 0.250000 2.745000 ;
      RECT 0.080000 2.935000 0.250000 3.105000 ;
      RECT 0.080000 3.295000 0.250000 3.465000 ;
      RECT 0.080000 3.655000 0.250000 3.825000 ;
      RECT 0.080000 4.015000 0.250000 4.185000 ;
      RECT 0.080000 4.375000 0.250000 4.545000 ;
      RECT 0.080000 4.735000 0.250000 4.905000 ;
      RECT 0.080000 5.095000 0.250000 5.265000 ;
      RECT 0.080000 5.455000 0.250000 5.625000 ;
      RECT 0.080000 5.815000 0.250000 5.985000 ;
      RECT 0.080000 6.175000 0.250000 6.345000 ;
      RECT 0.080000 6.535000 0.250000 6.705000 ;
      RECT 0.080000 6.895000 0.250000 7.065000 ;
      RECT 0.080000 7.255000 0.250000 7.425000 ;
      RECT 0.425000 0.080000 0.595000 0.250000 ;
      RECT 0.425000 7.590000 0.595000 7.760000 ;
      RECT 0.785000 0.080000 0.955000 0.250000 ;
      RECT 0.785000 7.590000 0.955000 7.760000 ;
      RECT 1.145000 0.080000 1.315000 0.250000 ;
      RECT 1.145000 7.590000 1.315000 7.760000 ;
      RECT 1.505000 0.080000 1.675000 0.250000 ;
      RECT 1.505000 7.590000 1.675000 7.760000 ;
      RECT 1.865000 0.080000 2.035000 0.250000 ;
      RECT 1.865000 7.590000 2.035000 7.760000 ;
      RECT 2.225000 0.080000 2.395000 0.250000 ;
      RECT 2.225000 7.590000 2.395000 7.760000 ;
      RECT 2.585000 0.080000 2.755000 0.250000 ;
      RECT 2.585000 7.590000 2.755000 7.760000 ;
      RECT 2.945000 0.080000 3.115000 0.250000 ;
      RECT 2.945000 7.590000 3.115000 7.760000 ;
      RECT 3.305000 0.080000 3.475000 0.250000 ;
      RECT 3.305000 7.590000 3.475000 7.760000 ;
      RECT 3.665000 0.080000 3.835000 0.250000 ;
      RECT 3.665000 7.590000 3.835000 7.760000 ;
      RECT 4.025000 0.080000 4.195000 0.250000 ;
      RECT 4.025000 7.590000 4.195000 7.760000 ;
      RECT 4.385000 0.080000 4.555000 0.250000 ;
      RECT 4.385000 7.590000 4.555000 7.760000 ;
      RECT 4.745000 0.080000 4.915000 0.250000 ;
      RECT 4.745000 7.590000 4.915000 7.760000 ;
      RECT 5.105000 0.080000 5.275000 0.250000 ;
      RECT 5.105000 7.590000 5.275000 7.760000 ;
      RECT 5.465000 0.080000 5.635000 0.250000 ;
      RECT 5.465000 7.590000 5.635000 7.760000 ;
      RECT 5.825000 0.080000 5.995000 0.250000 ;
      RECT 5.825000 7.590000 5.995000 7.760000 ;
      RECT 6.185000 0.080000 6.355000 0.250000 ;
      RECT 6.185000 7.590000 6.355000 7.760000 ;
      RECT 6.545000 0.080000 6.715000 0.250000 ;
      RECT 6.545000 7.590000 6.715000 7.760000 ;
      RECT 6.905000 0.080000 7.075000 0.250000 ;
      RECT 6.905000 7.590000 7.075000 7.760000 ;
      RECT 7.265000 0.080000 7.435000 0.250000 ;
      RECT 7.265000 7.590000 7.435000 7.760000 ;
      RECT 7.625000 0.080000 7.795000 0.250000 ;
      RECT 7.625000 7.590000 7.795000 7.760000 ;
      RECT 7.985000 0.080000 8.155000 0.250000 ;
      RECT 7.985000 7.590000 8.155000 7.760000 ;
      RECT 8.330000 0.415000 8.500000 0.585000 ;
      RECT 8.330000 0.775000 8.500000 0.945000 ;
      RECT 8.330000 1.135000 8.500000 1.305000 ;
      RECT 8.330000 1.495000 8.500000 1.665000 ;
      RECT 8.330000 1.855000 8.500000 2.025000 ;
      RECT 8.330000 2.215000 8.500000 2.385000 ;
      RECT 8.330000 2.575000 8.500000 2.745000 ;
      RECT 8.330000 2.935000 8.500000 3.105000 ;
      RECT 8.330000 3.295000 8.500000 3.465000 ;
      RECT 8.330000 3.655000 8.500000 3.825000 ;
      RECT 8.330000 4.015000 8.500000 4.185000 ;
      RECT 8.330000 4.375000 8.500000 4.545000 ;
      RECT 8.330000 4.735000 8.500000 4.905000 ;
      RECT 8.330000 5.095000 8.500000 5.265000 ;
      RECT 8.330000 5.455000 8.500000 5.625000 ;
      RECT 8.330000 5.815000 8.500000 5.985000 ;
      RECT 8.330000 6.175000 8.500000 6.345000 ;
      RECT 8.330000 6.535000 8.500000 6.705000 ;
      RECT 8.330000 6.895000 8.500000 7.065000 ;
      RECT 8.330000 7.255000 8.500000 7.425000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 8.580000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 7.510000 ;
      RECT 0.000000 7.510000 8.580000 7.840000 ;
      RECT 0.495000 0.470000 0.635000 3.760000 ;
      RECT 0.495000 3.760000 8.085000 4.080000 ;
      RECT 0.495000 4.080000 0.635000 7.370000 ;
      RECT 0.775000 0.330000 0.915000 3.620000 ;
      RECT 0.775000 4.220000 0.915000 7.510000 ;
      RECT 1.055000 0.470000 1.195000 3.760000 ;
      RECT 1.055000 4.080000 1.195000 7.370000 ;
      RECT 1.335000 0.330000 1.475000 3.620000 ;
      RECT 1.335000 4.220000 1.475000 7.510000 ;
      RECT 1.615000 0.470000 1.755000 3.760000 ;
      RECT 1.615000 4.080000 1.755000 7.370000 ;
      RECT 1.895000 0.330000 2.035000 3.620000 ;
      RECT 1.895000 4.220000 2.035000 7.510000 ;
      RECT 2.175000 0.470000 2.315000 3.760000 ;
      RECT 2.175000 4.080000 2.315000 7.370000 ;
      RECT 2.455000 0.330000 2.595000 3.620000 ;
      RECT 2.455000 4.220000 2.595000 7.510000 ;
      RECT 2.735000 0.470000 2.875000 3.760000 ;
      RECT 2.735000 4.080000 2.875000 7.370000 ;
      RECT 3.015000 0.330000 3.155000 3.620000 ;
      RECT 3.015000 4.220000 3.155000 7.510000 ;
      RECT 3.295000 0.470000 3.435000 3.760000 ;
      RECT 3.295000 4.080000 3.435000 7.370000 ;
      RECT 3.575000 0.330000 3.715000 3.620000 ;
      RECT 3.575000 4.220000 3.715000 7.510000 ;
      RECT 3.855000 0.470000 3.995000 3.760000 ;
      RECT 3.855000 4.080000 3.995000 7.370000 ;
      RECT 4.155000 0.470000 4.425000 3.760000 ;
      RECT 4.155000 4.080000 4.425000 7.370000 ;
      RECT 4.585000 0.470000 4.725000 3.760000 ;
      RECT 4.585000 4.080000 4.725000 7.370000 ;
      RECT 4.865000 0.330000 5.005000 3.620000 ;
      RECT 4.865000 4.220000 5.005000 7.510000 ;
      RECT 5.145000 0.470000 5.285000 3.760000 ;
      RECT 5.145000 4.080000 5.285000 7.370000 ;
      RECT 5.425000 0.330000 5.565000 3.620000 ;
      RECT 5.425000 4.220000 5.565000 7.510000 ;
      RECT 5.705000 0.470000 5.845000 3.760000 ;
      RECT 5.705000 4.080000 5.845000 7.370000 ;
      RECT 5.985000 0.330000 6.125000 3.620000 ;
      RECT 5.985000 4.220000 6.125000 7.510000 ;
      RECT 6.265000 0.470000 6.405000 3.760000 ;
      RECT 6.265000 4.080000 6.405000 7.370000 ;
      RECT 6.545000 0.330000 6.685000 3.620000 ;
      RECT 6.545000 4.220000 6.685000 7.510000 ;
      RECT 6.825000 0.470000 6.965000 3.760000 ;
      RECT 6.825000 4.080000 6.965000 7.370000 ;
      RECT 7.105000 0.330000 7.245000 3.620000 ;
      RECT 7.105000 4.220000 7.245000 7.510000 ;
      RECT 7.385000 0.470000 7.525000 3.760000 ;
      RECT 7.385000 4.080000 7.525000 7.370000 ;
      RECT 7.665000 0.330000 7.805000 3.620000 ;
      RECT 7.665000 4.220000 7.805000 7.510000 ;
      RECT 7.945000 0.470000 8.085000 3.760000 ;
      RECT 7.945000 4.080000 8.085000 7.370000 ;
      RECT 8.250000 0.330000 8.580000 7.510000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 4.015000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 0.750000 ;
      RECT 0.000000 0.750000 4.010000 0.890000 ;
      RECT 0.000000 0.890000 0.330000 1.310000 ;
      RECT 0.000000 1.310000 4.010000 1.450000 ;
      RECT 0.000000 1.450000 0.330000 1.870000 ;
      RECT 0.000000 1.870000 4.010000 2.010000 ;
      RECT 0.000000 2.010000 0.330000 2.430000 ;
      RECT 0.000000 2.430000 4.010000 2.570000 ;
      RECT 0.000000 2.570000 0.330000 2.990000 ;
      RECT 0.000000 2.990000 4.010000 3.130000 ;
      RECT 0.000000 3.130000 0.330000 3.645000 ;
      RECT 0.000000 3.785000 8.580000 4.055000 ;
      RECT 0.000000 4.195000 0.330000 4.710000 ;
      RECT 0.000000 4.710000 4.010000 4.850000 ;
      RECT 0.000000 4.850000 0.330000 5.270000 ;
      RECT 0.000000 5.270000 4.010000 5.410000 ;
      RECT 0.000000 5.410000 0.330000 5.830000 ;
      RECT 0.000000 5.830000 4.010000 5.970000 ;
      RECT 0.000000 5.970000 0.330000 6.390000 ;
      RECT 0.000000 6.390000 4.010000 6.530000 ;
      RECT 0.000000 6.530000 0.330000 6.950000 ;
      RECT 0.000000 6.950000 4.010000 7.090000 ;
      RECT 0.000000 7.090000 0.330000 7.510000 ;
      RECT 0.000000 7.510000 4.015000 7.840000 ;
      RECT 0.370000 3.780000 8.210000 3.785000 ;
      RECT 0.370000 4.055000 8.210000 4.060000 ;
      RECT 0.470000 0.470000 8.110000 0.610000 ;
      RECT 0.470000 1.030000 8.110000 1.170000 ;
      RECT 0.470000 1.590000 8.110000 1.730000 ;
      RECT 0.470000 2.150000 8.110000 2.290000 ;
      RECT 0.470000 2.710000 8.110000 2.850000 ;
      RECT 0.470000 3.270000 8.110000 3.640000 ;
      RECT 0.470000 4.200000 8.110000 4.570000 ;
      RECT 0.470000 4.990000 8.110000 5.130000 ;
      RECT 0.470000 5.550000 8.110000 5.690000 ;
      RECT 0.470000 6.110000 8.110000 6.250000 ;
      RECT 0.470000 6.670000 8.110000 6.810000 ;
      RECT 0.470000 7.230000 8.110000 7.370000 ;
      RECT 4.150000 0.610000 4.430000 1.030000 ;
      RECT 4.150000 1.170000 4.430000 1.590000 ;
      RECT 4.150000 1.730000 4.430000 2.150000 ;
      RECT 4.150000 2.290000 4.430000 2.710000 ;
      RECT 4.150000 2.850000 4.430000 3.270000 ;
      RECT 4.150000 3.640000 4.430000 3.780000 ;
      RECT 4.150000 4.060000 4.430000 4.200000 ;
      RECT 4.150000 4.570000 4.430000 4.990000 ;
      RECT 4.150000 5.130000 4.430000 5.550000 ;
      RECT 4.150000 5.690000 4.430000 6.110000 ;
      RECT 4.150000 6.250000 4.430000 6.670000 ;
      RECT 4.150000 6.810000 4.430000 7.230000 ;
      RECT 4.155000 0.000000 4.425000 0.470000 ;
      RECT 4.155000 7.370000 4.425000 7.840000 ;
      RECT 4.565000 0.000000 8.580000 0.330000 ;
      RECT 4.565000 7.510000 8.580000 7.840000 ;
      RECT 4.570000 0.750000 8.580000 0.890000 ;
      RECT 4.570000 1.310000 8.580000 1.450000 ;
      RECT 4.570000 1.870000 8.580000 2.010000 ;
      RECT 4.570000 2.430000 8.580000 2.570000 ;
      RECT 4.570000 2.990000 8.580000 3.130000 ;
      RECT 4.570000 4.710000 8.580000 4.850000 ;
      RECT 4.570000 5.270000 8.580000 5.410000 ;
      RECT 4.570000 5.830000 8.580000 5.970000 ;
      RECT 4.570000 6.390000 8.580000 6.530000 ;
      RECT 4.570000 6.950000 8.580000 7.090000 ;
      RECT 8.250000 0.330000 8.580000 0.750000 ;
      RECT 8.250000 0.890000 8.580000 1.310000 ;
      RECT 8.250000 1.450000 8.580000 1.870000 ;
      RECT 8.250000 2.010000 8.580000 2.430000 ;
      RECT 8.250000 2.570000 8.580000 2.990000 ;
      RECT 8.250000 3.130000 8.580000 3.645000 ;
      RECT 8.250000 4.195000 8.580000 4.710000 ;
      RECT 8.250000 4.850000 8.580000 5.270000 ;
      RECT 8.250000 5.410000 8.580000 5.830000 ;
      RECT 8.250000 5.970000 8.580000 6.390000 ;
      RECT 8.250000 6.530000 8.580000 6.950000 ;
      RECT 8.250000 7.090000 8.580000 7.510000 ;
    LAYER met4 ;
      RECT 0.315000 0.315000 2.325000 2.325000 ;
      RECT 0.315000 2.920000 2.325000 4.930000 ;
      RECT 0.315000 5.515000 2.325000 7.525000 ;
      RECT 3.290000 0.315000 5.300000 2.325000 ;
      RECT 3.290000 2.920000 5.300000 4.930000 ;
      RECT 3.290000 5.515000 5.300000 7.525000 ;
      RECT 6.255000 0.315000 8.265000 2.325000 ;
      RECT 6.255000 2.920000 8.265000 4.930000 ;
      RECT 6.255000 5.515000 8.265000 7.525000 ;
    LAYER via ;
      RECT 0.035000 0.265000 0.295000 0.525000 ;
      RECT 0.035000 0.585000 0.295000 0.845000 ;
      RECT 0.035000 0.905000 0.295000 1.165000 ;
      RECT 0.035000 1.225000 0.295000 1.485000 ;
      RECT 0.035000 1.545000 0.295000 1.805000 ;
      RECT 0.035000 1.865000 0.295000 2.125000 ;
      RECT 0.035000 2.185000 0.295000 2.445000 ;
      RECT 0.035000 2.505000 0.295000 2.765000 ;
      RECT 0.035000 2.825000 0.295000 3.085000 ;
      RECT 0.035000 3.145000 0.295000 3.405000 ;
      RECT 0.035000 4.435000 0.295000 4.695000 ;
      RECT 0.035000 4.755000 0.295000 5.015000 ;
      RECT 0.035000 5.075000 0.295000 5.335000 ;
      RECT 0.035000 5.395000 0.295000 5.655000 ;
      RECT 0.035000 5.715000 0.295000 5.975000 ;
      RECT 0.035000 6.035000 0.295000 6.295000 ;
      RECT 0.035000 6.355000 0.295000 6.615000 ;
      RECT 0.035000 6.675000 0.295000 6.935000 ;
      RECT 0.035000 6.995000 0.295000 7.255000 ;
      RECT 0.035000 7.315000 0.295000 7.575000 ;
      RECT 0.440000 0.035000 0.700000 0.295000 ;
      RECT 0.440000 7.545000 0.700000 7.805000 ;
      RECT 0.525000 3.790000 0.785000 4.050000 ;
      RECT 0.760000 0.035000 1.020000 0.295000 ;
      RECT 0.760000 7.545000 1.020000 7.805000 ;
      RECT 0.845000 3.790000 1.105000 4.050000 ;
      RECT 1.080000 0.035000 1.340000 0.295000 ;
      RECT 1.080000 7.545000 1.340000 7.805000 ;
      RECT 1.165000 3.790000 1.425000 4.050000 ;
      RECT 1.400000 0.035000 1.660000 0.295000 ;
      RECT 1.400000 7.545000 1.660000 7.805000 ;
      RECT 1.485000 3.790000 1.745000 4.050000 ;
      RECT 1.720000 0.035000 1.980000 0.295000 ;
      RECT 1.720000 7.545000 1.980000 7.805000 ;
      RECT 1.805000 3.790000 2.065000 4.050000 ;
      RECT 2.040000 0.035000 2.300000 0.295000 ;
      RECT 2.040000 7.545000 2.300000 7.805000 ;
      RECT 2.125000 3.790000 2.385000 4.050000 ;
      RECT 2.360000 0.035000 2.620000 0.295000 ;
      RECT 2.360000 7.545000 2.620000 7.805000 ;
      RECT 2.445000 3.790000 2.705000 4.050000 ;
      RECT 2.680000 0.035000 2.940000 0.295000 ;
      RECT 2.680000 7.545000 2.940000 7.805000 ;
      RECT 2.765000 3.790000 3.025000 4.050000 ;
      RECT 3.000000 0.035000 3.260000 0.295000 ;
      RECT 3.000000 7.545000 3.260000 7.805000 ;
      RECT 3.085000 3.790000 3.345000 4.050000 ;
      RECT 3.320000 0.035000 3.580000 0.295000 ;
      RECT 3.320000 7.545000 3.580000 7.805000 ;
      RECT 3.405000 3.790000 3.665000 4.050000 ;
      RECT 3.640000 0.035000 3.900000 0.295000 ;
      RECT 3.640000 7.545000 3.900000 7.805000 ;
      RECT 3.725000 3.790000 3.985000 4.050000 ;
      RECT 4.160000 0.500000 4.420000 0.760000 ;
      RECT 4.160000 0.820000 4.420000 1.080000 ;
      RECT 4.160000 1.140000 4.420000 1.400000 ;
      RECT 4.160000 1.460000 4.420000 1.720000 ;
      RECT 4.160000 1.780000 4.420000 2.040000 ;
      RECT 4.160000 2.100000 4.420000 2.360000 ;
      RECT 4.160000 2.420000 4.420000 2.680000 ;
      RECT 4.160000 2.740000 4.420000 3.000000 ;
      RECT 4.160000 3.060000 4.420000 3.320000 ;
      RECT 4.160000 3.380000 4.420000 3.640000 ;
      RECT 4.160000 4.200000 4.420000 4.460000 ;
      RECT 4.160000 4.520000 4.420000 4.780000 ;
      RECT 4.160000 4.840000 4.420000 5.100000 ;
      RECT 4.160000 5.160000 4.420000 5.420000 ;
      RECT 4.160000 5.480000 4.420000 5.740000 ;
      RECT 4.160000 5.800000 4.420000 6.060000 ;
      RECT 4.160000 6.120000 4.420000 6.380000 ;
      RECT 4.160000 6.440000 4.420000 6.700000 ;
      RECT 4.160000 6.760000 4.420000 7.020000 ;
      RECT 4.160000 7.080000 4.420000 7.340000 ;
      RECT 4.595000 3.790000 4.855000 4.050000 ;
      RECT 4.710000 0.035000 4.970000 0.295000 ;
      RECT 4.710000 7.545000 4.970000 7.805000 ;
      RECT 4.915000 3.790000 5.175000 4.050000 ;
      RECT 5.030000 0.035000 5.290000 0.295000 ;
      RECT 5.030000 7.545000 5.290000 7.805000 ;
      RECT 5.235000 3.790000 5.495000 4.050000 ;
      RECT 5.350000 0.035000 5.610000 0.295000 ;
      RECT 5.350000 7.545000 5.610000 7.805000 ;
      RECT 5.555000 3.790000 5.815000 4.050000 ;
      RECT 5.670000 0.035000 5.930000 0.295000 ;
      RECT 5.670000 7.545000 5.930000 7.805000 ;
      RECT 5.875000 3.790000 6.135000 4.050000 ;
      RECT 5.990000 0.035000 6.250000 0.295000 ;
      RECT 5.990000 7.545000 6.250000 7.805000 ;
      RECT 6.195000 3.790000 6.455000 4.050000 ;
      RECT 6.310000 0.035000 6.570000 0.295000 ;
      RECT 6.310000 7.545000 6.570000 7.805000 ;
      RECT 6.515000 3.790000 6.775000 4.050000 ;
      RECT 6.630000 0.035000 6.890000 0.295000 ;
      RECT 6.630000 7.545000 6.890000 7.805000 ;
      RECT 6.835000 3.790000 7.095000 4.050000 ;
      RECT 6.950000 0.035000 7.210000 0.295000 ;
      RECT 6.950000 7.545000 7.210000 7.805000 ;
      RECT 7.155000 3.790000 7.415000 4.050000 ;
      RECT 7.270000 0.035000 7.530000 0.295000 ;
      RECT 7.270000 7.545000 7.530000 7.805000 ;
      RECT 7.475000 3.790000 7.735000 4.050000 ;
      RECT 7.590000 0.035000 7.850000 0.295000 ;
      RECT 7.590000 7.545000 7.850000 7.805000 ;
      RECT 7.795000 3.790000 8.055000 4.050000 ;
      RECT 7.910000 0.035000 8.170000 0.295000 ;
      RECT 7.910000 7.545000 8.170000 7.805000 ;
      RECT 8.285000 0.265000 8.545000 0.525000 ;
      RECT 8.285000 0.585000 8.545000 0.845000 ;
      RECT 8.285000 0.905000 8.545000 1.165000 ;
      RECT 8.285000 1.225000 8.545000 1.485000 ;
      RECT 8.285000 1.545000 8.545000 1.805000 ;
      RECT 8.285000 1.865000 8.545000 2.125000 ;
      RECT 8.285000 2.185000 8.545000 2.445000 ;
      RECT 8.285000 2.505000 8.545000 2.765000 ;
      RECT 8.285000 2.825000 8.545000 3.085000 ;
      RECT 8.285000 3.145000 8.545000 3.405000 ;
      RECT 8.285000 4.435000 8.545000 4.695000 ;
      RECT 8.285000 4.755000 8.545000 5.015000 ;
      RECT 8.285000 5.075000 8.545000 5.335000 ;
      RECT 8.285000 5.395000 8.545000 5.655000 ;
      RECT 8.285000 5.715000 8.545000 5.975000 ;
      RECT 8.285000 6.035000 8.545000 6.295000 ;
      RECT 8.285000 6.355000 8.545000 6.615000 ;
      RECT 8.285000 6.675000 8.545000 6.935000 ;
      RECT 8.285000 6.995000 8.545000 7.255000 ;
      RECT 8.285000 7.315000 8.545000 7.575000 ;
    LAYER via2 ;
      RECT 0.025000 0.520000 0.305000 0.800000 ;
      RECT 0.025000 0.920000 0.305000 1.200000 ;
      RECT 0.025000 1.320000 0.305000 1.600000 ;
      RECT 0.025000 1.720000 0.305000 2.000000 ;
      RECT 0.025000 2.120000 0.305000 2.400000 ;
      RECT 0.025000 2.520000 0.305000 2.800000 ;
      RECT 0.025000 2.920000 0.305000 3.200000 ;
      RECT 0.025000 3.320000 0.305000 3.600000 ;
      RECT 0.025000 4.240000 0.305000 4.520000 ;
      RECT 0.025000 4.640000 0.305000 4.920000 ;
      RECT 0.025000 5.040000 0.305000 5.320000 ;
      RECT 0.025000 5.440000 0.305000 5.720000 ;
      RECT 0.025000 5.840000 0.305000 6.120000 ;
      RECT 0.025000 6.240000 0.305000 6.520000 ;
      RECT 0.025000 6.640000 0.305000 6.920000 ;
      RECT 0.025000 7.040000 0.305000 7.320000 ;
      RECT 0.490000 0.025000 0.770000 0.305000 ;
      RECT 0.490000 7.535000 0.770000 7.815000 ;
      RECT 0.890000 0.025000 1.170000 0.305000 ;
      RECT 0.890000 7.535000 1.170000 7.815000 ;
      RECT 0.950000 3.780000 1.230000 4.060000 ;
      RECT 1.290000 0.025000 1.570000 0.305000 ;
      RECT 1.290000 7.535000 1.570000 7.815000 ;
      RECT 1.350000 3.780000 1.630000 4.060000 ;
      RECT 1.690000 0.025000 1.970000 0.305000 ;
      RECT 1.690000 7.535000 1.970000 7.815000 ;
      RECT 1.750000 3.780000 2.030000 4.060000 ;
      RECT 2.090000 0.025000 2.370000 0.305000 ;
      RECT 2.090000 7.535000 2.370000 7.815000 ;
      RECT 2.150000 3.780000 2.430000 4.060000 ;
      RECT 2.490000 0.025000 2.770000 0.305000 ;
      RECT 2.490000 7.535000 2.770000 7.815000 ;
      RECT 2.550000 3.780000 2.830000 4.060000 ;
      RECT 2.890000 0.025000 3.170000 0.305000 ;
      RECT 2.890000 7.535000 3.170000 7.815000 ;
      RECT 2.950000 3.780000 3.230000 4.060000 ;
      RECT 3.290000 0.025000 3.570000 0.305000 ;
      RECT 3.290000 7.535000 3.570000 7.815000 ;
      RECT 3.350000 3.780000 3.630000 4.060000 ;
      RECT 3.690000 0.025000 3.970000 0.305000 ;
      RECT 3.690000 7.535000 3.970000 7.815000 ;
      RECT 3.750000 3.780000 4.030000 4.060000 ;
      RECT 4.150000 3.780000 4.430000 4.060000 ;
      RECT 4.550000 3.780000 4.830000 4.060000 ;
      RECT 4.610000 0.025000 4.890000 0.305000 ;
      RECT 4.610000 7.535000 4.890000 7.815000 ;
      RECT 4.950000 3.780000 5.230000 4.060000 ;
      RECT 5.010000 0.025000 5.290000 0.305000 ;
      RECT 5.010000 7.535000 5.290000 7.815000 ;
      RECT 5.350000 3.780000 5.630000 4.060000 ;
      RECT 5.410000 0.025000 5.690000 0.305000 ;
      RECT 5.410000 7.535000 5.690000 7.815000 ;
      RECT 5.750000 3.780000 6.030000 4.060000 ;
      RECT 5.810000 0.025000 6.090000 0.305000 ;
      RECT 5.810000 7.535000 6.090000 7.815000 ;
      RECT 6.150000 3.780000 6.430000 4.060000 ;
      RECT 6.210000 0.025000 6.490000 0.305000 ;
      RECT 6.210000 7.535000 6.490000 7.815000 ;
      RECT 6.550000 3.780000 6.830000 4.060000 ;
      RECT 6.610000 0.025000 6.890000 0.305000 ;
      RECT 6.610000 7.535000 6.890000 7.815000 ;
      RECT 6.950000 3.780000 7.230000 4.060000 ;
      RECT 7.010000 0.025000 7.290000 0.305000 ;
      RECT 7.010000 7.535000 7.290000 7.815000 ;
      RECT 7.350000 3.780000 7.630000 4.060000 ;
      RECT 7.410000 0.025000 7.690000 0.305000 ;
      RECT 7.410000 7.535000 7.690000 7.815000 ;
      RECT 7.810000 0.025000 8.090000 0.305000 ;
      RECT 7.810000 7.535000 8.090000 7.815000 ;
      RECT 8.275000 0.520000 8.555000 0.800000 ;
      RECT 8.275000 0.920000 8.555000 1.200000 ;
      RECT 8.275000 1.320000 8.555000 1.600000 ;
      RECT 8.275000 1.720000 8.555000 2.000000 ;
      RECT 8.275000 2.120000 8.555000 2.400000 ;
      RECT 8.275000 2.520000 8.555000 2.800000 ;
      RECT 8.275000 2.920000 8.555000 3.200000 ;
      RECT 8.275000 3.320000 8.555000 3.600000 ;
      RECT 8.275000 4.240000 8.555000 4.520000 ;
      RECT 8.275000 4.640000 8.555000 4.920000 ;
      RECT 8.275000 5.040000 8.555000 5.320000 ;
      RECT 8.275000 5.440000 8.555000 5.720000 ;
      RECT 8.275000 5.840000 8.555000 6.120000 ;
      RECT 8.275000 6.240000 8.555000 6.520000 ;
      RECT 8.275000 6.640000 8.555000 6.920000 ;
      RECT 8.275000 7.040000 8.555000 7.320000 ;
  END
END sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4
END LIBRARY
