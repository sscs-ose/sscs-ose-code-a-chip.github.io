# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield ;
  ORIGIN  0.440000  0.000000 ;
  SIZE  2.420000 BY  4.590000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT 0.000000 0.000000 1.540000 0.320000 ;
        RECT 0.280000 0.320000 0.420000 4.130000 ;
        RECT 0.840000 0.320000 0.980000 4.130000 ;
        RECT 1.400000 0.320000 1.540000 4.130000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT -0.440000 0.460000 -0.170000 4.270000 ;
        RECT -0.440000 4.270000  1.980000 4.590000 ;
        RECT  0.000000 0.460000  0.140000 4.270000 ;
        RECT  0.560000 0.460000  0.700000 4.270000 ;
        RECT  1.120000 0.460000  1.260000 4.270000 ;
        RECT  1.710000 0.460000  1.980000 4.270000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 0.450000 2.430000 0.530000 2.515000 ;
    END
  END SUB
  OBS
    LAYER met1 ;
      RECT -0.440000 0.460000 -0.170000 4.270000 ;
      RECT -0.440000 4.270000  1.980000 4.590000 ;
      RECT  0.000000 0.000000  1.540000 0.320000 ;
      RECT  0.000000 0.320000  0.140000 4.130000 ;
      RECT  0.280000 0.460000  0.420000 4.270000 ;
      RECT  0.560000 0.320000  0.700000 4.130000 ;
      RECT  0.840000 0.460000  0.980000 4.270000 ;
      RECT  1.120000 0.320000  1.260000 4.130000 ;
      RECT  1.400000 0.460000  1.540000 4.270000 ;
      RECT  1.710000 0.460000  1.980000 4.270000 ;
    LAYER via ;
      RECT -0.435000 0.585000 -0.175000 0.845000 ;
      RECT -0.435000 0.905000 -0.175000 1.165000 ;
      RECT -0.435000 1.225000 -0.175000 1.485000 ;
      RECT -0.435000 1.545000 -0.175000 1.805000 ;
      RECT -0.435000 1.865000 -0.175000 2.125000 ;
      RECT -0.435000 2.185000 -0.175000 2.445000 ;
      RECT -0.435000 2.505000 -0.175000 2.765000 ;
      RECT -0.435000 2.825000 -0.175000 3.085000 ;
      RECT -0.435000 3.145000 -0.175000 3.405000 ;
      RECT -0.435000 3.465000 -0.175000 3.725000 ;
      RECT -0.435000 3.785000 -0.175000 4.045000 ;
      RECT -0.180000 4.300000  0.080000 4.560000 ;
      RECT  0.140000 0.030000  0.400000 0.290000 ;
      RECT  0.140000 4.300000  0.400000 4.560000 ;
      RECT  0.460000 0.030000  0.720000 0.290000 ;
      RECT  0.460000 4.300000  0.720000 4.560000 ;
      RECT  0.780000 0.030000  1.040000 0.290000 ;
      RECT  0.780000 4.300000  1.040000 4.560000 ;
      RECT  1.100000 0.030000  1.360000 0.290000 ;
      RECT  1.100000 4.300000  1.360000 4.560000 ;
      RECT  1.420000 4.300000  1.680000 4.560000 ;
      RECT  1.715000 0.585000  1.975000 0.845000 ;
      RECT  1.715000 0.905000  1.975000 1.165000 ;
      RECT  1.715000 1.225000  1.975000 1.485000 ;
      RECT  1.715000 1.545000  1.975000 1.805000 ;
      RECT  1.715000 1.865000  1.975000 2.125000 ;
      RECT  1.715000 2.185000  1.975000 2.445000 ;
      RECT  1.715000 2.505000  1.975000 2.765000 ;
      RECT  1.715000 2.825000  1.975000 3.085000 ;
      RECT  1.715000 3.145000  1.975000 3.405000 ;
      RECT  1.715000 3.465000  1.975000 3.725000 ;
      RECT  1.715000 3.785000  1.975000 4.045000 ;
  END
END sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield
END LIBRARY
