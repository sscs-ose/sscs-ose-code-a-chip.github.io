magic
tech sky130A
magscale 1 2
timestamp 1762084523
<< pwell >>
rect -276 -579 276 579
<< nmos >>
rect -80 -369 80 431
<< ndiff >>
rect -138 419 -80 431
rect -138 -357 -126 419
rect -92 -357 -80 419
rect -138 -369 -80 -357
rect 80 419 138 431
rect 80 -357 92 419
rect 126 -357 138 419
rect 80 -369 138 -357
<< ndiffc >>
rect -126 -357 -92 419
rect 92 -357 126 419
<< psubdiff >>
rect -240 509 -144 543
rect 144 509 240 543
rect -240 447 -206 509
rect 206 447 240 509
rect -240 -509 -206 -447
rect 206 -509 240 -447
rect -240 -543 -144 -509
rect 144 -543 240 -509
<< psubdiffcont >>
rect -144 509 144 543
rect -240 -447 -206 447
rect 206 -447 240 447
rect -144 -543 144 -509
<< poly >>
rect -80 431 80 457
rect -80 -407 80 -369
rect -80 -441 -64 -407
rect 64 -441 80 -407
rect -80 -457 80 -441
<< polycont >>
rect -64 -441 64 -407
<< locali >>
rect -240 509 -144 543
rect 144 509 240 543
rect -240 447 -206 509
rect 206 447 240 509
rect -126 419 -92 435
rect -126 -373 -92 -357
rect 92 419 126 435
rect 92 -373 126 -357
rect -80 -441 -64 -407
rect 64 -441 80 -407
rect -240 -509 -206 -447
rect 206 -509 240 -447
rect -240 -543 -144 -509
rect 144 -543 240 -509
<< viali >>
rect -126 -357 -92 419
rect 92 -357 126 419
rect -64 -441 64 -407
<< metal1 >>
rect -132 419 -86 431
rect -132 -357 -126 419
rect -92 -357 -86 419
rect -132 -369 -86 -357
rect 86 419 132 431
rect 86 -357 92 419
rect 126 -357 132 419
rect 86 -369 132 -357
rect -76 -407 76 -401
rect -76 -441 -64 -407
rect 64 -441 76 -407
rect -76 -447 76 -441
<< labels >>
rlabel psubdiffcont 0 -526 0 -526 0 B
port 1 nsew
rlabel ndiffc -109 31 -109 31 0 D
port 2 nsew
rlabel ndiffc 109 31 109 31 0 S
port 3 nsew
rlabel polycont 0 -424 0 -424 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -223 -526 223 526
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
