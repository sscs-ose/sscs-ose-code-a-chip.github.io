# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15 ;
  ORIGIN  0.050000  0.000000 ;
  SIZE  4.500000 BY  7.590000 ;
  PIN BULK
    ANTENNADIFFAREA  1.618200 ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.995000 0.440000 5.595000 ;
        RECT 3.960000 1.995000 4.290000 5.595000 ;
      LAYER mcon ;
        RECT 0.190000 2.630000 0.360000 2.800000 ;
        RECT 0.190000 2.990000 0.360000 3.160000 ;
        RECT 0.190000 3.350000 0.360000 3.520000 ;
        RECT 0.190000 3.710000 0.360000 3.880000 ;
        RECT 0.190000 4.070000 0.360000 4.240000 ;
        RECT 0.190000 4.430000 0.360000 4.600000 ;
        RECT 0.190000 4.790000 0.360000 4.960000 ;
        RECT 4.040000 2.630000 4.210000 2.800000 ;
        RECT 4.040000 2.990000 4.210000 3.160000 ;
        RECT 4.040000 3.350000 4.210000 3.520000 ;
        RECT 4.040000 3.710000 4.210000 3.880000 ;
        RECT 4.040000 4.070000 4.210000 4.240000 ;
        RECT 4.040000 4.430000 4.210000 4.600000 ;
        RECT 4.040000 4.790000 4.210000 4.960000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.130000 2.600000 0.420000 4.990000 ;
        RECT 3.980000 2.600000 4.270000 4.990000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  3.732400 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3.980000 4.400000 5.260000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.806000 ;
    PORT
      LAYER li1 ;
        RECT 0.840000 1.880000 3.550000 2.050000 ;
        RECT 0.840000 5.540000 3.550000 5.710000 ;
      LAYER mcon ;
        RECT 0.850000 1.880000 1.020000 2.050000 ;
        RECT 0.850000 5.540000 1.020000 5.710000 ;
        RECT 1.330000 1.880000 1.500000 2.050000 ;
        RECT 1.330000 5.540000 1.500000 5.710000 ;
        RECT 1.810000 1.880000 1.980000 2.050000 ;
        RECT 1.810000 5.540000 1.980000 5.710000 ;
        RECT 2.290000 1.880000 2.460000 2.050000 ;
        RECT 2.290000 5.540000 2.460000 5.710000 ;
        RECT 2.770000 1.880000 2.940000 2.050000 ;
        RECT 2.770000 5.540000 2.940000 5.710000 ;
        RECT 3.250000 1.880000 3.420000 2.050000 ;
        RECT 3.250000 5.540000 3.420000 5.710000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.820000 1.820000 3.450000 2.110000 ;
        RECT 0.820000 5.480000 3.450000 5.770000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  3.551800 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2.330000 4.400000 3.610000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.690000 2.270000 0.915000 5.320000 ;
      RECT 1.165000 2.270000 1.695000 5.320000 ;
      RECT 1.935000 2.270000 2.465000 5.320000 ;
      RECT 2.705000 2.270000 3.235000 5.320000 ;
      RECT 3.485000 2.270000 3.710000 5.320000 ;
    LAYER mcon ;
      RECT 0.735000 2.475000 0.905000 2.645000 ;
      RECT 0.735000 2.835000 0.905000 3.005000 ;
      RECT 0.735000 3.195000 0.905000 3.365000 ;
      RECT 0.735000 3.555000 0.905000 3.725000 ;
      RECT 0.735000 3.915000 0.905000 4.085000 ;
      RECT 0.735000 4.275000 0.905000 4.445000 ;
      RECT 0.735000 4.635000 0.905000 4.805000 ;
      RECT 0.735000 4.995000 0.905000 5.165000 ;
      RECT 1.165000 2.475000 1.695000 5.165000 ;
      RECT 1.935000 2.425000 2.465000 5.115000 ;
      RECT 2.705000 2.475000 3.235000 5.165000 ;
      RECT 3.495000 2.475000 3.665000 2.645000 ;
      RECT 3.495000 2.835000 3.665000 3.005000 ;
      RECT 3.495000 3.195000 3.665000 3.365000 ;
      RECT 3.495000 3.555000 3.665000 3.725000 ;
      RECT 3.495000 3.915000 3.665000 4.085000 ;
      RECT 3.495000 4.275000 3.665000 4.445000 ;
      RECT 3.495000 4.635000 3.665000 4.805000 ;
      RECT 3.495000 4.995000 3.665000 5.165000 ;
    LAYER met1 ;
      RECT 0.650000 2.330000 0.970000 3.610000 ;
      RECT 0.690000 2.290000 0.970000 2.330000 ;
      RECT 0.690000 3.610000 0.970000 5.300000 ;
      RECT 1.115000 2.290000 1.745000 5.300000 ;
      RECT 1.885000 2.290000 2.515000 5.300000 ;
      RECT 2.655000 2.290000 3.285000 5.300000 ;
      RECT 3.430000 2.290000 3.710000 2.330000 ;
      RECT 3.430000 2.330000 3.750000 3.610000 ;
      RECT 3.430000 3.610000 3.710000 5.300000 ;
    LAYER via ;
      RECT 0.680000 2.330000 0.940000 2.590000 ;
      RECT 0.680000 2.670000 0.940000 2.930000 ;
      RECT 0.680000 3.010000 0.940000 3.270000 ;
      RECT 0.680000 3.350000 0.940000 3.610000 ;
      RECT 1.130000 3.980000 1.390000 4.240000 ;
      RECT 1.130000 4.320000 1.390000 4.580000 ;
      RECT 1.130000 4.660000 1.390000 4.920000 ;
      RECT 1.130000 5.000000 1.390000 5.260000 ;
      RECT 1.450000 3.980000 1.710000 4.240000 ;
      RECT 1.450000 4.320000 1.710000 4.580000 ;
      RECT 1.450000 4.660000 1.710000 4.920000 ;
      RECT 1.450000 5.000000 1.710000 5.260000 ;
      RECT 1.920000 2.330000 2.180000 2.590000 ;
      RECT 1.920000 2.670000 2.180000 2.930000 ;
      RECT 1.920000 3.010000 2.180000 3.270000 ;
      RECT 1.920000 3.350000 2.180000 3.610000 ;
      RECT 2.240000 2.330000 2.500000 2.590000 ;
      RECT 2.240000 2.670000 2.500000 2.930000 ;
      RECT 2.240000 3.010000 2.500000 3.270000 ;
      RECT 2.240000 3.350000 2.500000 3.610000 ;
      RECT 2.670000 3.980000 2.930000 4.240000 ;
      RECT 2.670000 4.320000 2.930000 4.580000 ;
      RECT 2.670000 4.660000 2.930000 4.920000 ;
      RECT 2.670000 5.000000 2.930000 5.260000 ;
      RECT 2.990000 3.980000 3.250000 4.240000 ;
      RECT 2.990000 4.320000 3.250000 4.580000 ;
      RECT 2.990000 4.660000 3.250000 4.920000 ;
      RECT 2.990000 5.000000 3.250000 5.260000 ;
      RECT 3.460000 2.330000 3.720000 2.590000 ;
      RECT 3.460000 2.670000 3.720000 2.930000 ;
      RECT 3.460000 3.010000 3.720000 3.270000 ;
      RECT 3.460000 3.350000 3.720000 3.610000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15
END LIBRARY
