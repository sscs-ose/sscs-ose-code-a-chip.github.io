* SKY130 Spice File.
.include "../../sonos_see_p/begin_of_life.pm3.spice"
.include "../../sonos_see_e/begin_of_life.pm3.spice"
.include "../../sonos_see_e/end_of_life/ff.spice"
.include "../../sonos_see_p/end_of_life/ff.spice"
