* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.3015+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.64774
+ k2 = 0.002296
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00225441
+ a0 = 1.75737
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.283503
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.3015+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.64774
+ k2 = 0.002296
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00225441
+ a0 = 1.75737
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.283503
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.058359263e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.451288897e-8
+ k1 = 0.64774
+ k2 = -9.370912500e-05 lk2 = 1.902148721e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.063707319e-09 lua = 4.641116804e-16
+ ub = 3.130202425e-18 lub = -7.028652274e-25
+ uc = 3.789249356e-11 luc = 9.122276612e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.176779101e-03 lu0 = 6.179225463e-10
+ a0 = 1.849196603e+00 la0 = -7.309167992e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.705724364e-01 lags = 1.029240538e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 9.025288750e-05 lpdiblc2 = 1.398008393e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.927296312e-03 ldelta = 6.131159568e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 2.990532506e+05 lat = -1.070845117e-1
+ ute = -3.115370919e-01 lute = 7.070414446e-7
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.751307275e-19 lub1 = 2.108595682e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.628429926e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.357283800e-7
+ k1 = 0.64774
+ k2 = -1.128156000e-02 lk2 = 6.332257971e-08 pk2 = 2.524354897e-29
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.561076335e+05 lvsat = -1.280885418e-1
+ ua = -3.110237112e-09 lua = 6.483580312e-16
+ ub = 3.171996025e-18 lub = -8.683574350e-25
+ uc = 4.861983037e-11 luc = 4.874519417e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.036878354e-03 lu0 = 1.171894531e-9
+ a0 = 2.218745970e+00 la0 = -2.194239909e-6
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.422712694e-01 lags = -1.809854002e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.221488000e-04 lpdiblc2 = 1.306183409e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.970993700e-02 ldelta = 6.735784214e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.761903100e+05 lat = -4.125279825e-1
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.565136819e-19 lub1 = 1.371407218e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.398697895e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.522488522e-8
+ k1 = 0.64774
+ k2 = 1.089799375e-01 lk2 = -1.723598900e-7
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 90748.0
+ ua = -2.247467100e-09 lua = -1.042455501e-15
+ ub = 1.852758050e-18 lub = 1.717019187e-24
+ uc = 7.920646150e-11 luc = -1.119695617e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.930255010e-03 lu0 = -5.789003708e-10
+ a0 = 9.687460835e-01 la0 = 2.554473696e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.459449270e-01 lags = 2.037651493e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.040698600e-03 lpdiblc2 = 1.965217428e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.711239350e-02 ldelta = 1.182632009e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.048988850e+05 lat = -7.683961238e-2
+ ute = -0.13298
+ ua1 = 7.976886000e-10 lua1 = -1.991078563e-16
+ ub1 = -3.072346025e-19 lub1 = 4.325160460e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.094349710e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.920234108e-8
+ k1 = 0.64774
+ k2 = -4.248662200e-02 lk2 = 4.874342021e-08 pk2 = -2.524354897e-29
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.005122150e+04 lvsat = 1.017122415e-3
+ ua = -3.146447850e-09 lua = 2.698316490e-16
+ ub = 3.137067850e-18 lub = -1.577520440e-25
+ uc = 5.217208400e-11 luc = 2.826647638e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.824002460e-03 lu0 = 1.035951789e-9
+ a0 = 1.056633090e+00 la0 = 1.271543119e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -2.318686300e-02 lags = 4.506552798e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.539712750e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.076895632e-8
+ nfactor = {2.595652800e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.518049980e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 9.396700000e-04 lpdiblc2 = 1.384183122e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.075824550e-02 ldelta = 2.110178763e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.489350000e-01 lkt1 = 8.405970375e-8
+ kt2 = -9.202608700e-02 lkt2 = 5.398314175e-8
+ at = 2.025317050e+05 lat = -7.338412137e-2
+ ute = 4.956445000e-02 lute = -2.664692609e-7
+ ua1 = 6.6129e-10
+ ub1 = -1.051962950e-20 lub1 = -6.136358374e-28
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.362382505e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.477893583e-9
+ k1 = 0.64774
+ k2 = 2.549013300e-02 lk2 = -1.649727040e-08 wk2 = -2.646977960e-23 pk2 = -6.310887242e-30
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.467314300e+04 lvsat = -3.418766744e-3
+ ua = -2.795142150e-09 lua = -6.733399654e-17
+ ub = 2.835418650e-18 lub = 1.317557757e-25
+ uc = 9.281615400e-11 luc = -1.074166980e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.917118940e-03 lu0 = -1.316675266e-11
+ a0 = 1.274688670e+00 la0 = -8.212453103e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.698134110e-01 lags = -2.250173321e-8
+ b0 = 7.194076050e-08 lb0 = -6.904514489e-14
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.098287250e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.284023132e-8
+ nfactor = {2.478947200e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.682769980e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.007644950e-02 lpdiblc2 = 3.401205191e-08 ppdiblc2 = -1.262177448e-29
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.216615250e-02 ldelta = 1.015304889e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.964241050e-01 lkt1 = -6.231262773e-8
+ kt2 = -1.717199800e-02 lkt2 = -1.785807017e-8
+ at = 1.874319130e+05 lat = -5.889209600e-2
+ ute = -7.139720000e-02 lute = -1.503763173e-7
+ ua1 = 4.451523300e-10 lua1 = 2.074381288e-16
+ ub1 = 5.295630895e-19 lub1 = -5.189580254e-25 wub1 = 4.591774808e-41 pub1 = 3.503246161e-46
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.620328200e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 8.381159745e-9
+ k1 = 0.64774
+ k2 = -3.375434500e-02 lk2 = 1.074037836e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.428050850e+04 lvsat = -3.238253033e-3
+ ua = -3.060750500e-09 lua = 5.477944238e-17
+ ub = 3.039400000e-18 lub = 3.797535000e-26
+ uc = 8.249041000e-11 luc = -5.994408998e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.319304050e-03 lu0 = 2.616786430e-10
+ a0 = 1.294423900e+00 la0 = -9.119780303e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.120937500e-01 lags = 4.034880938e-9
+ b0 = -2.398025350e-07 lb0 = 7.427883522e-14
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.416210500e-02 lpdiblc2 = 5.887793202e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.684411500e-02 ldelta = 8.002355629e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.526100000e-01 lkt1 = 9.493837500e-9
+ kt2 = -0.056015
+ at = 1.297958650e+05 lat = -3.239392293e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.178348025e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.151505243e-7
+ k1 = 0.64774
+ k2 = 2.535185090e-04 wk2 = 1.439826494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.123303443e-09 wua = 8.311482974e-16
+ ub = 3.234534534e-18 wub = -1.357957497e-24
+ uc = 5.089054169e-11 wuc = -1.083874332e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.277990689e-03 wu0 = -1.662296595e-10
+ a0 = 1.762570880e+00 wa0 = -3.666307265e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.111731961e-01 wags = -1.950582250e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.357346608e-03 wpdiblc2 = -3.600456115e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.354475070e-03 wdelta = 7.243626489e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.178348025e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.151505243e-7
+ k1 = 0.64774
+ k2 = 2.535185090e-04 wk2 = 1.439826494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.123303443e-09 wua = 8.311482974e-16
+ ub = 3.234534534e-18 wub = -1.357957497e-24
+ uc = 5.089054169e-11 wuc = -1.083874332e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.277990689e-03 wu0 = -1.662296595e-10
+ a0 = 1.762570880e+00 wa0 = -3.666307265e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.111731961e-01 wags = -1.950582250e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.357346608e-03 wpdiblc2 = -3.600456115e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.354475070e-03 wdelta = 7.243626489e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.900797910e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.209229527e-07 wvth0 = -1.110712680e-07 pvth0 = 1.800668911e-12
+ k1 = 0.64774
+ k2 = 1.834052690e-02 lk2 = -1.439680650e-07 wk2 = -1.299502666e-07 pk2 = 1.148978224e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.328819191e-09 lua = 1.635853976e-15 wua = 1.868879105e-15 pua = -8.260077794e-21
+ ub = 3.545774003e-18 lub = -2.477388364e-24 wub = -2.929529449e-24 pub = 1.250931985e-29
+ uc = 1.049570611e-11 luc = 3.215327925e-16 wuc = 1.931308587e-16 puc = -1.623547039e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.017186517e-03 lu0 = 2.075936007e-09 wu0 = 1.125031646e-09 pu0 = -1.027811717e-14
+ a0 = 2.092105355e+00 la0 = -2.623012041e-06 wa0 = -1.712360477e-06 pa0 = 1.333813241e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.540913612e-01 lags = -3.416178644e-07 wags = -5.887581414e-07 pags = 3.133752910e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.080502740e-04 lpdiblc2 = 1.962394283e-08 wpdiblc2 = 1.397917910e-09 ppdiblc2 = -3.978580764e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.202606045e-02 ldelta = 1.224252176e-07 wdelta = 1.265603573e-07 pdelta = -4.308142442e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 2.990532506e+05 lat = -1.070845117e-1
+ ute = -3.115370919e-01 lute = 7.070414446e-7
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.751307275e-19 lub1 = 2.108595682e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.473509370e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.860935325e-07 wvth0 = -8.141494660e-07 pvth0 = 4.584682806e-12
+ k1 = 0.64774
+ k2 = -7.395726696e-02 lk2 = 2.215081242e-07 wk2 = 4.418260033e-07 pk2 = -1.115112861e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.377756714e+05 lvsat = -4.514735550e-01 wvsat = -5.757105034e-01 pvsat = 2.279669666e-6
+ ua = -3.639276963e-09 lua = 2.865189138e-15 wua = 3.729412466e-15 pua = -1.562732477e-20
+ ub = 3.986487150e-18 lub = -4.222502247e-24 wub = -5.741672105e-24 pub = 2.364470173e-29
+ uc = 6.639541898e-11 luc = 1.001839045e-16 wuc = -1.253071987e-16 puc = -3.626119416e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.284907704e-03 lu0 = 4.975577035e-09 wu0 = 5.300940392e-09 pu0 = -2.681367183e-14
+ a0 = 3.424311646e+00 la0 = -7.898215898e-06 wa0 = -8.498512260e-06 pa0 = 4.020959693e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.892182002e-01 lags = -8.766863652e-07 wags = -1.035887400e-06 pags = 4.904272991e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.444947878e-03 lpdiblc2 = 9.514708398e-09 wpdiblc2 = -1.496445557e-08 ppdiblc2 = 2.500510075e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.338684151e-02 ldelta = -5.739852094e-08 wdelta = -9.641394332e-08 pdelta = 4.521082425e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 5.786534212e+05 lat = -1.214231287e+00 wat = -1.427243051e+00 pat = 5.651525671e-6
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -2.439533039e-19 lub1 = 4.833797650e-25 wub1 = 6.163966964e-25 pub1 = -2.440776819e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-8.952321824e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.795667381e-07 wvth0 = 3.914970542e-06 pvth0 = -4.683210129e-12
+ k1 = 0.64774
+ k2 = 2.815367481e-01 lk2 = -4.751712719e-07 wk2 = -1.216421636e-06 pk2 = 2.134637950e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.845648890e+05 lvsat = 7.681583582e-01 wvsat = 3.350669729e+00 pvsat = -5.415053994e-6
+ ua = -5.072658005e-10 lua = -3.272769738e-15 wua = -1.226737156e-14 pua = 1.572237272e-20
+ ub = -7.882126803e-19 lub = 5.134715744e-24 wub = 1.861725378e-23 pub = -2.409270328e-29
+ uc = 2.333871217e-10 luc = -2.270780849e-16 wuc = -1.086880838e-15 puc = 1.521831997e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 6.095460906e-03 lu0 = -4.451904602e-09 wu0 = -2.231279611e-08 pu0 = 2.730234828e-14
+ a0 = -1.379631464e+00 la0 = 1.516311611e-06 wa0 = 1.655464799e-05 pa0 = -8.888333860e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.500989599e-01 lags = -1.191972434e-06 wags = -3.553982431e-06 pags = 9.839109728e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -6.473021715e-03 lpdiblc2 = 2.699169931e-08 wpdiblc2 = 2.419581170e-08 ppdiblc2 = -5.173923304e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.447425998e-03 ldelta = 2.066668481e-08 wdelta = 1.660825445e-07 pdelta = -6.231924940e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.124757619e-01 lkt1 = 4.333512119e-07 wkt1 = 1.558803504e-06 pkt1 = -3.054865167e-12
+ kt2 = -2.051672798e-01 lkt2 = 2.942021378e-07 wkt2 = 1.058271699e-06 pkt2 = -2.073947962e-12
+ at = -8.405999133e+05 lat = 1.567150435e+00 wat = 7.370137138e+00 pat = -1.158914015e-5
+ ute = -0.13298
+ ua1 = 8.435353413e-10 lua1 = -2.889560076e-16 wua1 = -3.231919265e-16 pua1 = 6.333753779e-22
+ ub1 = 4.252388548e-20 lub1 = -7.804390684e-26 wub1 = -2.465586786e-24 pub1 = 3.599140310e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.951140259e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.549425915e-08 wvth0 = 1.308925558e-06 pvth0 = -8.790359643e-13
+ k1 = 0.64774
+ k2 = -1.828955162e-01 lk2 = 2.027837260e-07 wk2 = 9.897981781e-07 pk2 = -1.085891424e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.190611777e+05 lvsat = -4.049347925e-01 wvsat = -2.319322127e+00 pvsat = 2.861716617e-6
+ ua = -3.206959457e-09 lua = 6.681080769e-16 wua = 4.265704008e-16 pua = -2.807609054e-21
+ ub = 3.110224872e-18 lub = -5.560284719e-25 wub = 1.892268388e-25 pub = 2.807609054e-30
+ uc = 4.266515319e-11 luc = 5.132830861e-17 wuc = 6.701813906e-17 puc = -1.625720340e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.775068428e-03 lu0 = 1.854788317e-09 wu0 = 3.449554645e-10 pu0 = -5.772304582e-15
+ a0 = -1.497635286e+00 la0 = 1.688567689e-06 wa0 = 1.800605438e-05 pa0 = -1.100702434e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.423560121e+00 lags = 1.835051409e-06 wags = 9.871788445e-06 pags = -9.759159307e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.345965092e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.436982996e-07 wvoff = -4.970645018e-07 pvoff = 7.255899064e-13
+ nfactor = {2.742976056e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.002356225e-07 wnfactor = -1.038540265e-06 pnfactor = 1.516009152e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.741299014e-02 lpdiblc2 = -7.875906499e-09 wpdiblc2 = -1.161269901e-07 ppdiblc2 = 1.530969768e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.520137611e-03 ldelta = 3.197033833e-09 wdelta = 3.692550728e-08 pdelta = 1.262177356e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.216556273e-01 lkt1 = 1.548015204e-07 wkt1 = -1.923031553e-07 pkt1 = -4.986872209e-13
+ kt2 = 5.809619276e-02 lkt2 = -9.009671626e-08 wkt2 = -1.058271699e-06 pkt2 = 1.015676263e-12
+ at = 9.217763381e+05 lat = -1.005478298e+00 wat = -5.070241678e+00 pat = 6.570702823e-6
+ ute = 3.300117136e-01 lute = -6.758521539e-07 wute = -1.976984379e-06 pute = 2.885902947e-12
+ ua1 = 5.192954496e-10 lua1 = 1.843531742e-16 wua1 = 1.000976099e-15 pua1 = -1.299578898e-21
+ ub1 = -9.458320519e-21 lub1 = -2.162881622e-27 wub1 = -7.481589408e-27 pub1 = 1.092125014e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.436049725e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.991655480e-08 wvth0 = 5.193095541e-08 pvth0 = 3.273646055e-13
+ k1 = 0.64774
+ k2 = 5.859115358e-02 lk2 = -2.898310533e-08 wk2 = -2.333422682e-07 pk2 = 8.801761978e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.729136042e+04 lvsat = -7.692121042e-02 wvsat = 1.225311034e-01 pvsat = 5.181479794e-7
+ ua = -1.814808597e-09 lua = -6.680087105e-16 wua = -6.910761385e-15 pua = 4.234395127e-21
+ ub = 1.545566720e-18 lub = 9.456521889e-25 wub = 9.092679615e-24 pub = -5.737479748e-30
+ uc = 9.889274851e-11 luc = -2.636125998e-18 wuc = -4.283633319e-17 puc = -5.713920428e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.490833180e-03 lu0 = -7.516669036e-10 wu0 = -1.109373802e-08 pu0 = 5.205981487e-15
+ a0 = 1.049581319e+00 la0 = -7.561234469e-07 wa0 = 1.586871311e-06 pa0 = 4.751286610e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.647098407e-01 lags = 1.187593136e-07 wags = 7.409168983e-07 pags = -9.958053407e-13
+ b0 = 1.276335481e-06 lb0 = -1.224962978e-12 wb0 = -8.490257731e-12 pb0 = 8.148524858e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.803403491e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.525795049e-08 wvoff = 4.970645018e-07 pvoff = -2.285254047e-13
+ nfactor = {2.331623944e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.455956666e-08 wnfactor = 1.038540265e-06 pnfactor = -4.774688868e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.820576011e-02 lpdiblc2 = 4.550418905e-08 wpdiblc2 = 1.278007260e-07 ppdiblc2 = -8.101264862e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.231590859e-03 ldelta = 4.433716578e-09 wdelta = 1.264278630e-07 pdelta = 4.031784975e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.172493476e-01 lkt1 = -1.373524065e-07 wkt1 = -1.263074176e-06 pkt1 = 5.289852666e-13
+ kt2 = -1.717199800e-02 lkt2 = -1.785807017e-8
+ at = -2.961663665e+05 lat = 1.634422130e-01 wat = 3.409076744e+00 pat = -1.567323033e-6
+ ute = -3.518444636e-01 lute = -2.144068786e-08 wute = 1.976984379e-06 pute = -9.089185683e-13
+ ua1 = 5.413001391e-10 lua1 = 1.632341736e-16 wua1 = -6.777841728e-16 pua1 = 3.116112735e-22
+ ub1 = 5.285017805e-19 lub1 = -5.184700886e-25 wub1 = 7.481589408e-27 pub1 = -3.439660730e-33
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.351597619e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.815075964e-08 wvth0 = 1.220440718e-06 pvth0 = -2.098577580e-13
+ k1 = 0.64774
+ k2 = 2.265497763e-03 lk2 = -3.087385067e-09 wk2 = -2.539182075e-07 pk2 = 9.747740787e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.859804205e+05 lvsat = 1.820429908e-01 wvsat = 4.090490232e+00 pvsat = -1.306121230e-6
+ ua = -4.060526255e-09 lua = 3.644599824e-16 wua = 7.047817205e-15 pua = -2.183061379e-21
+ ub = 4.511979923e-18 lub = -4.181562813e-25 wub = -1.038080197e-23 pub = 3.215453409e-30
+ uc = 1.551521309e-10 luc = -2.850137704e-17 wuc = -5.122213897e-16 puc = 1.586605755e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.117949080e-03 lu0 = 3.392665616e-10 wu0 = 1.419431325e-09 pu0 = -5.469481180e-16
+ a0 = -3.888856237e+00 la0 = 1.514323219e-06 wa0 = 3.653900463e-05 pa0 = -1.131795668e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.054057549e+00 lags = -1.981682952e-07 wags = -4.525458319e-06 pags = 1.425410665e-12
+ b0 = -4.254451602e-06 lb0 = 1.317816384e-12 wb0 = 2.830085910e-11 pb0 = -8.766191108e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.364520468e-01 lpdiblc2 = 9.067291935e-08 wpdiblc2 = 4.391065910e-07 ppdiblc2 = -2.241355201e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.407641743e-03 ldelta = 5.272277184e-09 wdelta = 1.722624257e-07 pdelta = 1.924540953e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.037045606e-01 lkt1 = -5.654622351e-09 wkt1 = -3.447539066e-07 pkt1 = 1.067875226e-13
+ kt2 = -0.056015
+ at = 1.297958650e+05 lat = -3.239392293e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.933528311e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -8.468693289e-9
+ k1 = 0.64774
+ k2 = 1.012318950e-02 wk2 = -3.543763201e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.111169900e-09 wua = 7.698812081e-16
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.905656756e-03 wu0 = 1.713832557e-9
+ a0 = 1.759731627e+00 wa0 = -2.232655504e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.900699199e-01 wags = -8.849938464e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.244490933e-04 wpdiblc2 = 4.644693329e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.317621807e-02 wdelta = 2.284237544e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899606391e+05 wat = -2.201860255e-2
+ ute = -1.174447810e-01 wute = -5.315259861e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463681985e-19 wub1 = -1.147123000e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.933528311e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -8.468693289e-9
+ k1 = 0.64774
+ k2 = 1.012318950e-02 wk2 = -3.543763201e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.111169900e-09 wua = 7.698812081e-16
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.905656756e-03 wu0 = 1.713832557e-9
+ a0 = 1.759731627e+00 wa0 = -2.232655504e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.900699199e-01 wags = -8.849938464e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.244490933e-04 wpdiblc2 = 4.644693329e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.317621807e-02 wdelta = 2.284237544e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899606391e+05 wat = -2.201860255e-2
+ ute = -1.174447810e-01 wute = -5.315259861e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463681985e-19 wub1 = -1.147123000e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.958342625e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.975157389e-08 wvth0 = -8.201465116e-08 pvth0 = 5.854074382e-13
+ k1 = 0.64774
+ k2 = -9.778015386e-04 lk2 = 8.836111340e-08 wk2 = -3.240433758e-08 pk2 = -2.414426533e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.156450601e-09 lua = 3.604230637e-16 wua = 9.985214917e-16 pua = -1.819919497e-21
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.723062933e-03 lu0 = 1.453401181e-09 wu0 = 2.610178682e-09 pu0 = -7.134691068e-15
+ a0 = 1.839346741e+00 la0 = -6.337164009e-07 wa0 = -4.360816335e-07 pa0 = 3.293386986e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.364234381e-01 lags = 4.270125842e-07 wags = 5.394034202e-09 pags = -7.473681406e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.513579764e-03 lpdiblc2 = 1.781415019e-08 wpdiblc2 = 8.494995703e-09 ppdiblc2 = -3.064744433e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.180500002e-02 ldelta = 1.091455284e-08 wdelta = 6.227848174e-09 pdelta = 1.322474834e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 3.077306500e+05 lat = -1.414448437e-01 wat = -4.381564292e-02 pat = 1.734989920e-7
+ ute = -1.020658852e-01 lute = -1.224121660e-07 wute = -1.057703492e-06 pute = 4.188241402e-12
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.706099845e-19 lub1 = 1.929585561e-25 wub1 = -2.282703075e-26 pub1 = 9.038933501e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.562254245e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.588854773e-07 wvth0 = 2.405409533e-07 pvth0 = -6.918321165e-13
+ k1 = 0.64774
+ k2 = 1.761123283e-02 lk2 = 1.475318454e-08 wk2 = -2.053979644e-08 pk2 = -7.112488210e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.918974676e-09 lua = -5.799222339e-16 wua = 9.231953519e-17 pua = 1.768413700e-21
+ ub = 2.778925643e-18 lub = 1.161803665e-24 wub = 3.557865500e-25 pub = -3.542801771e-30
+ uc = -2.490208249e-12 luc = 1.293025723e-16 wuc = 2.225237496e-16 puc = -5.096436848e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.270770451e-03 lu0 = -7.153836651e-10 wu0 = 3.229270096e-10 pu0 = 1.922253743e-15
+ a0 = 1.334565902e+00 la0 = 1.365089524e-06 wa0 = 2.053445716e-06 pa0 = -6.564518938e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.780976250e-01 lags = 2.619932225e-07 wags = 3.014441000e-08 pags = -8.453734412e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.408670462e-03 lpdiblc2 = 1.739873559e-08 wpdiblc2 = 4.493997166e-09 ppdiblc2 = -1.480449037e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.266166368e-02 ldelta = 7.522378933e-09 wdelta = 8.235728198e-09 pdelta = 1.242967805e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.848968128e+05 lat = -5.102855685e-02 wat = 5.605098002e-02 pat = -2.219478681e-7
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.678553806e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.063318401e-07 wvth0 = -5.206561873e-07 pvth0 = 7.999239797e-13
+ k1 = 0.64774
+ k2 = 5.025413836e-02 lk2 = -4.921874958e-08 wk2 = -4.858368854e-08 pk2 = -1.616586457e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.157275256e+05 lvsat = -7.681583582e-01 wvsat = -1.195264989e+00 pvsat = 2.342420561e-6
+ ua = -3.009981238e-09 lua = -4.015721230e-16 wua = 3.698347649e-16 pua = 1.224553229e-21
+ ub = 2.903708702e-18 lub = 9.172600652e-25 wub = -2.472665970e-26 pub = -2.797091008e-30
+ uc = -3.224380557e-11 luc = 1.876121847e-16 wuc = 2.543954352e-16 puc = -5.721042207e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 9.146796540e-04 lu0 = 1.942215275e-09 wu0 = 3.847030380e-09 pu0 = -4.984107836e-15
+ a0 = 2.005699166e+00 la0 = 4.983611068e-08 wa0 = -5.392337249e-07 pa0 = -1.483515403e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -3.616324866e-01 lags = 1.515704309e-06 wags = 1.554652311e-06 pags = -3.833027801e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.195305916e-03 lpdiblc2 = 2.873909442e-08 wpdiblc2 = 2.784291210e-08 ppdiblc2 = -6.056252642e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.454495035e-02 ldelta = 6.084054077e-08 wdelta = 2.069701677e-07 pdelta = -2.651730373e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.702242381e-01 lkt1 = -4.333512119e-07 wkt1 = -6.743004561e-07 pkt1 = 1.321460319e-12
+ kt2 = 9.507727976e-02 lkt2 = -2.942021378e-07 wkt2 = -4.577825797e-07 pkt2 = 8.971394105e-13
+ at = 1.100532716e+06 lat = -1.649471019e+00 wat = -2.431414080e+00 pat = 4.652861783e-6
+ ute = -0.13298
+ ua1 = 9.067491425e-10 lua1 = -4.128392545e-16 wua1 = -6.423835679e-16 pua1 = 1.258911197e-21
+ ub1 = -9.396030676e-19 lub1 = 1.602532782e-24 wub1 = 2.493563087e-24 pub1 = -4.886760259e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.400441623e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.043006338e-08 wvth0 = 2.097629888e-08 pvth0 = 9.275958033e-15
+ k1 = 0.64774
+ k2 = 1.178609028e-01 lk2 = -1.479077240e-07 wk2 = -5.288406828e-07 pk2 = 6.848892828e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.903544755e+05 lvsat = 4.085198429e-01 wvsat = 1.262799853e+00 pvsat = -1.245739592e-6
+ ua = -3.166649539e-09 lua = -1.728755708e-16 wua = 2.230295818e-16 pua = 1.438852095e-21
+ ub = 3.637729034e-18 lub = -1.542261147e-25 wub = -2.474351625e-24 pub = 7.787490349e-31
+ uc = 1.880736170e-10 luc = -1.339961729e-16 wuc = -6.672070671e-16 puc = 7.732050320e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.010540999e-03 lu0 = -1.117218323e-09 wu0 = -5.893437261e-09 pu0 = 9.234539802e-15
+ a0 = 2.394186849e+00 la0 = -5.172587843e-07 wa0 = -1.645304523e-06 pa0 = 1.310714442e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 9.797326015e-01 lags = -4.423533787e-07 wags = -2.263393022e-06 pags = 1.740363875e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {6.714228767e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.097271768e-06 wnfactor = -2.109097576e-05 pnfactor = 3.078755187e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.406441466e-02 lpdiblc2 = 3.876627591e-08 wpdiblc2 = 4.281495479e-08 ppdiblc2 = -8.241796572e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.790876938e-02 ldelta = -1.572877660e-08 wdelta = -1.266175852e-07 pdelta = 2.217816850e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.518139565e-01 lkt1 = 2.696493796e-07 wkt1 = 9.698578519e-07 pkt1 = -1.078599771e-12
+ kt2 = -2.421483668e-01 lkt2 = 1.980629998e-07 wkt2 = 4.577825797e-07 pkt2 = -4.393568308e-13
+ at = -6.358975664e+05 lat = 8.852830864e-01 wat = 2.795073820e+00 pat = -2.976503929e-6
+ ute = -6.632089890e-01 lute = 7.740017667e-07 wute = 3.038182250e-06 pute = -4.434986540e-12
+ ua1 = 5.903123375e-10 lua1 = 4.907937160e-17 wua1 = 6.423835679e-16 pua1 = -6.165276293e-22
+ ub1 = 4.828937376e-19 lub1 = -4.739569296e-25 wub1 = -2.493563087e-24 pub1 = 2.393197173e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.275042699e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.509774930e-09 wvth0 = -2.936790011e-08 pvth0 = 5.759380302e-14
+ k1 = 0.64774
+ k2 = -5.698295111e-02 lk2 = 1.989866482e-08 wk2 = 3.502373848e-07 pk2 = -1.588058926e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.909500921e+04 lvsat = 9.233069989e-02 wvsat = 3.153996828e-01 pvsat = -3.364722780e-7
+ ua = -3.837572347e-09 lua = 4.710425946e-16 wua = 3.302977849e-15 pua = -1.517128254e-21
+ ub = 3.978470502e-18 lub = -4.812527382e-25 wub = -3.192019875e-24 pub = 1.467531137e-30
+ uc = 4.437997240e-11 luc = 3.913802512e-18 wuc = 2.324203695e-16 puc = -9.021240019e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 7.616481119e-04 lu0 = 1.041156625e-09 wu0 = 7.736401608e-09 pu0 = -3.846698053e-15
+ a0 = 1.689496340e+00 la0 = 1.590679314e-07 wa0 = -1.644314317e-06 pa0 = 1.301210942e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.335959417e-01 lags = -1.101487195e-07 wags = -6.167960424e-07 pags = 1.600424235e-13
+ b0 = -1.318902119e-06 lb0 = 1.265816309e-12 wb0 = 4.614129815e-12 pb0 = -4.428411089e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.612495872e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.098774460e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.163536690e-03 lpdiblc2 = 3.214315827e-08 wpdiblc2 = -2.894381490e-08 ppdiblc2 = -1.354748652e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.747194670e-03 ldelta = 1.705779472e-08 wdelta = 1.288737721e-07 pdelta = -2.342614519e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.368988850e-01 lkt1 = -3.259036032e-08 wkt1 = -1.539762416e-07 pkt1 = -1.615587134e-27
+ kt2 = -1.010471396e-02 lkt2 = -2.464089603e-08 wkt2 = -3.568552991e-08 pkt2 = 3.424918733e-14
+ at = 5.003923223e+05 lat = -2.052711343e-01 wat = -6.130651057e-01 pat = 2.944574051e-7
+ ute = 5.911019272e-01 lute = -4.298231351e-07 wute = -2.784327241e-06 pute = 1.153166944e-12
+ ua1 = 4.070694500e-10 lua1 = 2.249467329e-16
+ ub1 = 4.795829717e-19 lub1 = -4.707794221e-25 wub1 = 2.544921246e-25 pub1 = -2.442488166e-31
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.985272472e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.578741128e-08 wvth0 = -4.793508287e-07 pvth0 = 2.644734544e-13
+ k1 = 0.64774
+ k2 = -3.423243876e-03 lk2 = -4.725410586e-09 wk2 = -2.251934869e-07 pk2 = 1.057484507e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.335596538e+05 lvsat = -1.809744204e-01 wvsat = -1.562513180e+00 pvsat = 5.268981605e-7
+ ua = -2.881034865e-09 lua = 3.127448699e-17 wua = 1.092095741e-15 pua = -5.006752053e-22
+ ub = 2.752719524e-18 lub = 8.228627404e-26 wub = -1.497596022e-24 pub = 6.885197713e-31
+ uc = -8.003748206e-12 luc = 2.799721806e-17 wuc = 3.116175797e-16 puc = -1.266233176e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.523871802e-03 lu0 = 6.907242834e-10 wu0 = 4.419163943e-09 pu0 = -2.321598036e-15
+ a0 = 5.729119855e+00 la0 = -1.698148980e-06 wa0 = -1.202598461e-05 pa0 = 4.903094012e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -6.795654428e-02 lags = 2.123900360e-07 wags = 1.140037398e-06 pags = -6.476617509e-13
+ b0 = 4.396340397e-06 lb0 = -1.361766438e-12 wb0 = -1.538043272e-11 pb0 = 4.764089033e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.612495872e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.098774460e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.097044619e-02 lpdiblc2 = 3.849088492e-08 wpdiblc2 = -1.440059720e-07 ppdiblc2 = 3.935234022e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.786927005e-02 ldelta = -7.824829430e-09 wdelta = -1.077854093e-07 pdelta = 8.537791347e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.729718544e-01 lkt1 = 2.996918734e-08 wkt1 = 5.004227853e-09 pkt1 = -7.309127084e-14
+ kt2 = -7.957261347e-02 lkt2 = 7.296970774e-09 wkt2 = 1.189517664e-07 pkt2 = -3.684530963e-14
+ at = 1.131592643e+05 lat = -2.724073588e-02 wat = 8.400481814e-02 pat = -2.602049242e-8
+ ute = -2.308989607e-01 lute = -5.190822693e-08 wute = -8.461833648e-07 pute = 2.621052972e-13
+ ua1 = 8.9635e-10
+ ub1 = -4.312183725e-19 lub1 = -5.203850413e-26 wub1 = -8.483070821e-25 pub1 = 2.627631187e-31
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.114931867e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.684847086e-8
+ k1 = 0.64774
+ k2 = -1.062828730e-02 wk2 = 2.784187983e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844218308e-09 wua = -4.416044384e-17
+ ub = 2.872303364e-18 wub = 7.104071401e-26
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.489161177e-03 wu0 = -6.550465836e-11
+ a0 = 1.872875643e+00 wa0 = -3.673476921e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.448266893e-01 wags = -2.554745677e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.696427525e-03 wpdiblc2 = -1.368653756e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.473866424e-02 wdelta = -1.241612479e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.908560200e-01 wkt1 = -3.200032162e-8
+ kt2 = -0.055045
+ at = 2.871894475e+05 wat = -1.356813637e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.114931867e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.684847086e-8
+ k1 = 0.64774
+ k2 = -1.062828730e-02 wk2 = 2.784187983e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844218308e-09 wua = -4.416044384e-17
+ ub = 2.872303364e-18 wub = 7.104071401e-26
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.489161177e-03 wu0 = -6.550465836e-11
+ a0 = 1.872875643e+00 wa0 = -3.673476921e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.448266893e-01 wags = -2.554745677e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.696427525e-03 wpdiblc2 = -1.368653756e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.473866424e-02 wdelta = -1.241612479e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.908560200e-01 wkt1 = -3.200032162e-8
+ kt2 = -0.055045
+ at = 2.871894475e+05 wat = -1.356813637e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.489798341e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.983843416e-07 wvth0 = 8.004734853e-08 pvth0 = -2.642547665e-13
+ k1 = 0.64774
+ k2 = -2.910344165e-02 lk2 = 1.470576098e-07 wk2 = 5.336193312e-08 pk2 = -2.031332442e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.824908567e-09 lua = -1.537007083e-16 wua = -1.248212545e-17 pua = -2.521514948e-22
+ ub = 2.915415159e-18 lub = -3.431591099e-25 wub = -6.042430730e-26 pub = 1.046428703e-30
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.667052143e-03 lu0 = -1.415967615e-09 wu0 = -2.684201268e-10 pu0 = 1.615156400e-15
+ a0 = 1.832789622e+00 la0 = 3.190747085e-07 wa0 = -4.160863688e-07 pa0 = 3.879476823e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.384334850e-01 lags = 5.088830839e-08 wags = -3.056751988e-07 pags = 3.995844738e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.864751278e-03 lpdiblc2 = -1.339814998e-09 wpdiblc2 = -4.856278219e-09 ppdiblc2 = 2.776061882e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.940244608e-02 ldelta = 4.247496246e-08 wdelta = -1.693978866e-08 pdelta = 3.600723346e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.903670107e-01 lkt1 = -3.892391985e-09 wkt1 = -6.367864001e-08 pkt1 = 2.521514948e-13
+ kt2 = -0.055045
+ at = 3.022161518e+05 lat = -1.196088098e-01 wat = -2.699974336e-02 pat = 1.069122338e-7
+ ute = -4.489223769e-01 lute = 1.251052827e-6
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.521398367e-19 lub1 = 1.599779781e-26 wub1 = -7.914986241e-26 pub1 = 6.300131173e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.901567753e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.545973451e-08 wvth0 = 3.907134669e-08 pvth0 = -1.020000433e-13
+ k1 = 0.64774
+ k2 = 9.356532334e-03 lk2 = -5.234272139e-09 wk2 = 4.632070755e-09 pk2 = -1.017517169e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.838017356e-09 lua = -1.017931809e-16 wua = -1.545515533e-16 pua = 3.104079223e-22
+ ub = 2.797647912e-18 lub = 1.231697489e-25 wub = 2.986949021e-25 pub = -3.755935860e-31
+ uc = 7.357684716e-11 luc = -5.767433966e-17 wuc = -9.434977028e-18 puc = 6.052333669e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.390057084e-03 lu0 = -3.191364314e-10 wu0 = -4.082541032e-11 pu0 = 7.139382213e-16
+ a0 = 2.161300974e+00 la0 = -9.817481187e-07 wa0 = -4.675985585e-07 pa0 = 5.919230752e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.010784530e-01 lags = -1.971701038e-07 wags = -3.448730810e-07 pags = 5.547982877e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 5.084365503e-05 lpdiblc2 = 9.802555713e-09 wpdiblc2 = 4.335773577e-11 ppdiblc2 = 8.359285348e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.225946006e-02 ldelta = 7.075940138e-08 wdelta = 9.462207101e-09 pdelta = -6.853806924e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.032778113e+05 lat = -1.238127156e-1
+ ute = -1.439208871e-01 lute = 4.332317780e-08 wute = 3.336311932e-08 pute = -1.321096117e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.737917953e-19 lub1 = 1.017341409e-25 wub1 = 1.582997248e-25 pub1 = -3.102278857e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.447139919e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.195717603e-07 wvth0 = -1.305514161e-07 pvth0 = 2.304181662e-13
+ k1 = 0.64774
+ k2 = 4.910264199e-02 lk2 = -8.312671054e-08 wk2 = -4.507231781e-08 pk2 = 8.723300379e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.889959278e-09 wua = 3.840038595e-18
+ ub = 2.860497637e-18 wub = 1.070410758e-25
+ uc = 4.414740990e-11 wuc = 2.144821557e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.987773017e-03 lu0 = 4.692397691e-10 wu0 = 5.747416245e-10 pu0 = -4.924192753e-16
+ a0 = 2.000068427e+00 la0 = -6.657726332e-07 wa0 = -5.220633599e-07 pa0 = 6.986604698e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 9.917818660e-02 lags = 3.944789433e-07 wags = 1.494571661e-07 pags = -4.139654141e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.854832885e-03 lpdiblc2 = 1.353720531e-08 wpdiblc2 = 1.155768432e-08 ppdiblc2 = -1.420591618e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 6.868625346e-02 ldelta = -3.982300699e-08 wdelta = -4.683489872e-08 pdelta = 4.179018389e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.362938622e+05 lat = -1.885159214e-01 wat = -1.009456466e-01 pat = 1.978282309e-7
+ ute = -1.218144053e-01 wute = -3.404834221e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.592687422e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.983254636e-07 wvth0 = -2.253401056e-07 pvth0 = 3.687859556e-13
+ k1 = 0.64774
+ k2 = -5.912097746e-02 lk2 = 7.485271795e-08 wk2 = 1.084750902e-08 pk2 = 5.604036574e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.202233871e-09 lua = 4.558428375e-16 wua = 3.315403722e-16 pua = -4.783605620e-22
+ ub = 2.754845221e-18 lub = 1.542261147e-25 wub = 2.179125102e-25 pub = -1.618445763e-31
+ uc = -8.073608746e-11 luc = 1.822986853e-16 wuc = 1.525007079e-16 puc = -1.913038757e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.453452581e-04 lu0 = 3.012748690e-09 wu0 = 2.538745100e-09 pu0 = -3.359373349e-15
+ a0 = 2.021805015e+00 la0 = -6.975026184e-07 wa0 = -5.097641043e-07 pa0 = 6.807066314e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.228024469e-01 lags = 2.140184293e-07 wags = 4.478827735e-08 pags = -2.611750037e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {-1.639628767e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.097271768e-06 wnfactor = 4.383260695e-06 pnfactor = -6.398464799e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.828704778e-03 lpdiblc2 = 5.240661209e-09 wpdiblc2 = -1.174828784e-08 ppdiblc2 = 1.981497668e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.732044066e-03 ldelta = 5.353415017e-08 wdelta = -2.544854537e-08 pdelta = 1.057145459e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.296557883e-01 lkt1 = -9.005812553e-08 wkt1 = -1.253062194e-08 pkt1 = 1.829157538e-14
+ kt2 = -9.202608700e-02 lkt2 = 5.398314175e-8
+ at = 2.257723765e+05 lat = -2.718218264e-02 wat = 1.674992195e-01 pat = -1.940341623e-7
+ ute = 5.842142473e-01 lute = -1.030625326e-06 wute = -7.657076719e-07 pute = 1.068039706e-12
+ ua1 = 8.009714800e-10 lua1 = -1.531007404e-16
+ ub1 = -3.348293300e-19 lub1 = 3.108527845e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.668850332e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.342716901e-10 wvth0 = 9.071972059e-08 pvth0 = 6.544753744e-14
+ k1 = 0.64774
+ k2 = 6.768922514e-02 lk2 = -4.685337399e-08 wk2 = -2.993770009e-08 pk2 = 4.474764103e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.375099767e+05 lvsat = -1.319654014e-02 wvsat = 1.529327771e-02 pvsat = -1.467772328e-8
+ ua = -2.704513502e-09 lua = -2.184428689e-17 wua = -1.521695294e-16 pua = -1.411998392e-23
+ ub = 2.954136129e-18 lub = -3.704333489e-26 wub = -6.841668763e-26 pub = 1.129598713e-31
+ uc = 1.462490040e-10 luc = -3.555025625e-17 wuc = -7.821885175e-17 puc = 3.012922168e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.645139086e-03 lu0 = -2.502034365e-10 wu0 = -1.056510003e-09 pu0 = 9.117273614e-17
+ a0 = 8.189900392e-01 la0 = 4.568990548e-07 wa0 = 1.010205856e-06 pa0 = -7.780845376e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 5.508194773e-01 lags = -1.007959156e-07 wags = -3.643776574e-07 pags = 1.315220022e-13
+ b0 = 5.068653630e-07 lb0 = -4.864640321e-13 wb0 = -9.533618939e-13 pb0 = 9.149890777e-19
+ b1 = 2.325991428e-07 lb1 = -2.232370273e-13 wb1 = -7.092873608e-13 pb1 = 6.807385445e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.713350413e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.283542951e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.938584188e-02 lpdiblc2 = 2.752082236e-08 wpdiblc2 = 8.326858090e-09 ppdiblc2 = 5.478553759e-16
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.288997439e-02 ldelta = 7.314576543e-09 wdelta = -2.098212208e-08 pdelta = 6.284804841e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.818528621e-01 lkt1 = -3.996198396e-08 wkt1 = -1.689367379e-08 pkt1 = 2.247901439e-14
+ kt2 = -2.180719750e-02 lkt2 = -1.340943745e-8
+ at = 3.201167328e+05 lat = -1.177291786e-01 wat = -6.333308374e-02 pat = 2.750714066e-8
+ ute = -4.440801196e-01 lute = -4.371980700e-08 wute = 3.723548224e-07 pute = -2.421577241e-14
+ ua1 = 4.070694500e-10 lua1 = 2.249467329e-16
+ ub1 = 5.630394850e-19 lub1 = -5.508768107e-25 wub1 = -2.869859255e-41 pub1 = 2.736911063e-47
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.962467785e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.040833412e-08 wvth0 = 4.285145148e-07 pvth0 = -8.985361922e-14
+ k1 = 0.64774
+ k2 = -1.087877167e-01 lk2 = 3.428190003e-08 wk2 = 9.610472591e-08 pk2 = -1.320036433e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.181905300e+05 lvsat = -4.314424499e-03 wvsat = 9.052395782e-03 pvsat = -1.180847781e-8
+ ua = -2.354576561e-09 lua = -1.827277954e-16 wua = -5.132851588e-16 pua = 1.519029267e-22
+ ub = 2.093061851e-18 lub = 3.588355646e-25 wub = 5.139627657e-25 pub = -1.547890823e-31
+ uc = 1.137836906e-10 luc = -2.062432842e-17 wuc = -5.976079263e-17 puc = 2.164312900e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.535319273e-03 lu0 = -1.997137772e-10 wu0 = -1.714539952e-09 pu0 = 3.937020055e-16
+ a0 = 2.112123481e+00 la0 = -1.376190449e-07 wa0 = -9.963231017e-07 pa0 = 1.444171505e-13
+ keta = -1.176195491e-02 lketa = -3.760962317e-10 wketa = -2.494545072e-09 pketa = 1.146867097e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.315787691e-01 wags = -7.830478701e-8
+ b0 = -1.642697271e-06 lb0 = 5.017973888e-13 wb0 = 3.034996672e-12 pb0 = -9.186587729e-19
+ b1 = -5.551192378e-07 lb1 = 1.389164982e-13 wb1 = 1.692779494e-12 pb1 = -4.236116918e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.713350413e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.283542951e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -8.380581845e-02 lpdiblc2 = 5.713790659e-08 wpdiblc2 = 4.760408645e-08 ppdiblc2 = -1.750985036e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -8.821774543e-03 ldelta = 3.568655312e-08 wdelta = 9.558212866e-08 pdelta = -4.730560944e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.770573649e-01 lkt1 = 3.808286201e-09 wkt1 = 1.746257551e-08 pkt1 = 6.683728776e-15
+ kt2 = -7.233698973e-02 lkt2 = 9.821634527e-09 wkt2 = 9.688746978e-08 pkt2 = -4.454401423e-14
+ at = 1.424300879e+05 lat = -3.603774366e-02 wat = -5.253572802e-03 pat = 8.050855116e-10
+ ute = -6.280372522e-01 lute = 4.085448470e-08 wute = 3.648493470e-07 pute = -2.076513008e-14
+ ua1 = 7.087088751e-10 lua1 = 8.626800716e-17 wua1 = 5.721924709e-16 pua1 = -2.630654885e-22
+ ub1 = -3.120318652e-19 lub1 = -1.485627575e-25 wub1 = -1.211754179e-24 pub1 = 5.571039838e-31
+ uc1 = 3.224846359e-11 luc1 = -1.341323549e-17 wuc1 = -8.896638057e-17 puc1 = 4.090229347e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.868565732e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.099485795e-8
+ k1 = 0.64774
+ k2 = 1.825397216e-02 wk2 = -2.467105478e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.694093041e-09 wua = -2.017015980e-16
+ ub = 2.757516609e-18 wub = 1.914977057e-25
+ uc = 7.060795191e-11 wuc = -6.319424287e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.964266806e-03 wu0 = -5.640795556e-10
+ a0 = 1.254982334e+00 wa0 = 2.810683114e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.160462985e-01 wags = 2.281646240e-7
+ b0 = -2.317672267e-07 wb0 = 2.432160641e-13
+ b1 = -2.826228170e-07 wb1 = 2.965838189e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.669956697e-03 wpdiblc2 = -1.340875322e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.201855896e-02 wdelta = 9.323282458e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.504878364e-01 wkt1 = -7.436261271e-8
+ kt2 = -0.055045
+ at = 2.636706353e+05 wat = 1.111245810e-2
+ ute = -2.995155341e-01 wute = 8.149135942e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.868565732e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 2.099485795e-8
+ k1 = 0.64774
+ k2 = 1.825397216e-02 wk2 = -2.467105478e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.694093041e-09 wua = -2.017015980e-16
+ ub = 2.757516609e-18 wub = 1.914977057e-25
+ uc = 7.060795191e-11 wuc = -6.319424287e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.964266806e-03 wu0 = -5.640795556e-10
+ a0 = 1.254982334e+00 wa0 = 2.810683114e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.160462985e-01 wags = 2.281646240e-7
+ b0 = -2.317672267e-07 wb0 = 2.432160641e-13
+ b1 = -2.826228170e-07 wb1 = 2.965838189e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.669956697e-03 wpdiblc2 = -1.340875322e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.201855896e-02 wdelta = 9.323282458e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.504878364e-01 wkt1 = -7.436261271e-8
+ kt2 = -0.055045
+ at = 2.636706353e+05 wat = 1.111245810e-2
+ ute = -2.995155341e-01 wute = 8.149135942e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.473870848e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.141672607e-07 wvth0 = -2.656387943e-08 pvth0 = 3.785556599e-13
+ k1 = 0.64774
+ k2 = 5.608266786e-02 lk2 = -3.011069606e-07 wk2 = -3.603219982e-08 pk2 = 2.671697597e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.631805821e-09 lua = -4.957907057e-16 wua = -2.151237613e-16 pua = 1.068370643e-22
+ ub = 2.606521276e-18 lub = 1.201885103e-24 wub = 2.637283164e-25 pub = -5.749376039e-31
+ uc = 6.347964166e-11 luc = 5.673956748e-17 wuc = 1.161010228e-18 puc = -5.954238863e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.826837477e-03 lu0 = 1.093903106e-09 wu0 = -4.360985367e-10 pu0 = -1.018696915e-15
+ a0 = 1.007702303e+00 la0 = 1.968287221e-06 wa0 = 4.497586132e-07 pa0 = -1.342732630e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -2.774021344e-01 lags = 1.284352114e-06 wags = 3.405814684e-07 pags = -8.948099773e-13
+ b0 = -1.632795400e-07 lb0 = -5.451448640e-13 wb0 = 1.713452227e-13 pb0 = 5.720739300e-19
+ b1 = -2.943582889e-07 lb1 = 9.341142260e-14 wb1 = 3.088989997e-13 pb1 = -9.802576005e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.201194122e-03 lpdiblc2 = 3.081339272e-08 wpdiblc2 = -5.894832481e-10 ppdiblc2 = -5.980893059e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -4.572089290e-03 ldelta = 1.320574124e-07 wdelta = 8.219040816e-09 pdelta = -5.800041038e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.802123333e-01 lkt1 = 2.365995638e-07 wkt1 = -7.433493815e-08 pkt1 = -2.202826068e-16
+ kt2 = -0.055045
+ at = 2.517890566e+05 lat = 9.457439664e-02 wat = 2.591834958e-02 pat = -1.178511947e-7
+ ute = -4.152788368e-01 lute = 9.214469487e-07 wute = -3.530546367e-08 pute = 3.458877493e-13
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -2.934552795e-19 lub1 = 1.140833394e-24 wub1 = 6.914628064e-26 pub1 = -5.503871073e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.936522514e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.309687672e-07 wvth0 = 4.273949232e-08 pvth0 = 1.041316336e-13
+ k1 = 0.64774
+ k2 = -1.750953645e-02 lk2 = -9.700229611e-09 wk2 = 3.282526961e-08 pk2 = -5.488604854e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.884318497e-09 lua = 5.040963646e-16 wua = -1.059632286e-16 pua = -3.254113550e-22
+ ub = 3.074396941e-18 lub = -6.507855606e-25 wub = 8.275024716e-27 pub = 4.365935679e-31
+ uc = 7.780871988e-11 wuc = -1.387589580e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.925877599e-03 lu0 = 7.017289831e-10 wu0 = -6.031143868e-10 pu0 = -3.573559030e-16
+ a0 = 1.750763067e+00 la0 = -9.740476378e-07 wa0 = -3.678089968e-08 pa0 = 5.838422060e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -4.260503108e-02 lags = 3.546142846e-07 wags = 1.207274798e-07 pags = -2.424314594e-14
+ b0 = -3.524277357e-07 lb0 = 2.038347040e-13 wb0 = 3.698369610e-13 pb0 = -2.139037307e-19
+ b1 = -2.619058222e-07 lb1 = -3.509223225e-14 wb1 = 2.748434460e-13 pb1 = 3.682571834e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.447540278e-03 lpdiblc2 = 2.032506669e-08 wpdiblc2 = -1.422332907e-09 ppdiblc2 = -2.683016622e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.405204175e-02 ldelta = -2.088449046e-08 wdelta = -1.340688454e-08 pdelta = 2.763284756e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.204611965e-01 wkt1 = -7.439056858e-8
+ kt2 = -0.055045
+ at = 3.001146598e+05 lat = -9.678291079e-02 wat = 3.319404806e-03 pat = -2.836502311e-8
+ ute = -1.339493575e-01 lute = -1.925474569e-07 wute = 2.289901608e-08 pute = 1.154125606e-13
+ ua1 = 6.9609e-10
+ ub1 = 1.088390903e-19 lub1 = -4.521517372e-25 wub1 = -1.382925613e-25 pub1 = 2.710188470e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.604815752e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 9.587465425e-8
+ k1 = 0.64774
+ k2 = -2.245926453e-02 wk2 = 3.002460378e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.627093665e-09 wua = -2.720106097e-16
+ ub = 2.742321135e-18 wub = 2.310552609e-25
+ uc = 7.780871988e-11 wuc = -1.387589580e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.283948263e-03 wu0 = -7.854620857e-10
+ a0 = 1.253736590e+00 wa0 = 2.611357764e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.383437045e-01 wags = 1.083569500e-7
+ b0 = -2.484171711e-07 wb0 = 2.606884825e-13
+ b1 = -2.798123064e-07 wb1 = 2.936344747e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.181879512e-02 wpdiblc2 = -2.791393564e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.339533020e-02 wdelta = 6.933055621e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.204611965e-01 wkt1 = -7.439056858e-8
+ kt2 = -0.055045
+ at = 2.507293245e+05 wat = -1.115439191e-2
+ ute = -2.322003879e-01 wute = 8.179048722e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-6.192292011e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.777068469e-07 wvth0 = 2.573414800e-07 pvth0 = -2.357011990e-13
+ k1 = 0.64774
+ k2 = -1.237086042e-01 lk2 = 1.477987236e-07 wk2 = 7.862563539e-08 pk2 = -7.094535590e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.632068748e+04 lvsat = 1.130420365e-01 wvsat = 8.126465968e-02 pvsat = -1.186260870e-7
+ ua = -1.827593103e-09 lua = -1.167070946e-15 wua = -1.111004901e-15 pua = 1.224721916e-21
+ ub = 1.881969554e-18 lub = 1.255898219e-24 wub = 1.133906489e-24 pub = -1.317937080e-30
+ uc = 1.248148530e-10 luc = -6.861720286e-17 wuc = -6.320403791e-17 puc = 7.200675545e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.276213592e-03 lu0 = -2.908209315e-09 wu0 = -2.740638068e-09 pu0 = 2.854068140e-15
+ a0 = 3.834535850e-01 la0 = 1.270395617e-06 wa0 = 1.209518610e-06 pa0 = -1.384401841e-12
+ keta = -1.064964207e-02 lketa = -2.817839987e-09 wketa = -2.025713750e-09 pketa = 2.957035647e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 5.798021734e-01 lags = -6.444190000e-07 wags = -3.298465217e-07 pags = 6.396675177e-13
+ b0 = 2.265659339e-07 lb0 = -6.933565875e-13 wb0 = -2.377578379e-13 pb0 = 7.276070162e-19
+ b1 = 4.614707060e-07 lb1 = -1.082087877e-12 wb1 = -4.842664360e-13 pb1 = 1.135540854e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 6.589225566e-03 lpdiblc2 = 7.633864163e-09 wpdiblc2 = -1.464517283e-08 ppdiblc2 = 1.730355429e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.080112907e-02 ldelta = 1.229057814e-07 wdelta = 4.332183544e-08 pdelta = -6.222699649e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -2.347183038e-01 lkt1 = -4.171131877e-07 wkt1 = -3.220374283e-07 pkt1 = 3.615025035e-13
+ kt2 = -2.187393836e-01 lkt2 = 2.389528765e-07 wkt2 = 1.329726801e-07 pkt2 = -1.941068697e-13
+ at = 2.789164211e+05 lat = -4.114611415e-02 wat = 1.117299654e-01 pat = -1.793804405e-7
+ ute = -2.225308097e-01 lute = -1.411516677e-08 wute = 8.088897753e-08 pute = 1.315978778e-15
+ ua1 = 1.009910354e-09 lua1 = -4.580992619e-16 wua1 = -2.192600366e-16 pua1 = 3.200648385e-22
+ ub1 = -5.470613180e-19 lub1 = 6.206584290e-25 wub1 = 2.227158238e-25 pub1 = -3.251094238e-31
+ uc1 = 9.220990490e-11 luc1 = -1.491439784e-16 wuc1 = -1.072179433e-16 puc1 = 1.565113927e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.576541407e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.266601828e-07 wvth0 = 8.103284053e-08 pvth0 = -6.648898218e-14
+ k1 = 0.64774
+ k2 = 3.043344871e-02 lk2 = -1.391116839e-10 wk2 = 9.158437180e-09 pk2 = -4.274212413e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.998624180e+05 lvsat = -3.431963944e-02 wvsat = -5.013924951e-02 pvsat = 7.488814879e-9
+ ua = -3.126366219e-09 lua = 7.942655241e-17 wua = 2.905218682e-16 pua = -1.203934001e-22
+ ub = 3.371974735e-18 lub = -1.741342528e-25 wub = -5.068956849e-25 pub = 2.568228064e-31
+ uc = 6.331084342e-11 luc = -9.588729639e-18 wuc = 8.816288089e-18 puc = 2.885247571e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.434693424e-03 lu0 = -1.810603339e-10 wu0 = 2.137292544e-10 pu0 = 1.861410254e-17
+ a0 = 2.207727740e+00 la0 = -4.804515036e-07 wa0 = -4.471327105e-07 pa0 = 2.055692637e-13
+ keta = -1.358565664e-02 wketa = 1.055334071e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.145143683e-01 lags = 2.195130097e-08 wags = 3.338223495e-07 pags = 2.711318581e-15
+ b0 = -1.596017004e-06 lb0 = 1.055867387e-12 wb0 = 1.253398656e-12 pb0 = -7.035304290e-19
+ b1 = -1.842898358e-06 lb1 = 1.129530332e-12 wb1 = 1.468735565e-12 pb1 = -7.388528164e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.609295702e-02 lpdiblc2 = -1.487342103e-09 wpdiblc2 = -2.890452252e-08 ppdiblc2 = 3.098896515e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.875671355e-02 ldelta = 2.735514197e-08 wdelta = -6.150706422e-09 pdelta = -1.474572444e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.659154525e-01 lkt1 = -3.271724239e-09 wkt1 = 7.132144044e-08 pkt1 = -1.602367078e-14
+ kt2 = 6.281688107e-02 lkt2 = -3.127074853e-08 wkt2 = -8.880433880e-08 pkt2 = 1.874362413e-14
+ at = 4.456865844e+05 lat = -2.012037784e-01 wat = -1.951058348e-01 pat = 1.151052187e-7
+ ute = -7.493814870e-02 lute = -1.557672232e-07 wute = -1.502202354e-08 pute = 9.336656205e-14
+ ua1 = -1.397507771e-11 lua1 = 5.245747813e-16 wua1 = 4.418432853e-16 pua1 = -3.144290747e-22
+ ub1 = 1.211546764e-18 lub1 = -1.067165678e-24 wub1 = -6.805422414e-25 pub1 = 5.417925043e-31
+ uc1 = -9.113814615e-11 luc1 = 2.682431357e-17 wuc1 = 7.260996253e-17 puc1 = -1.607843991e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.200118850e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.765626203e-08 wvth0 = -6.915785883e-08 pvth0 = 2.561191848e-15
+ k1 = 0.64774
+ k2 = -5.242811922e-02 lk2 = 3.795649417e-08 wk2 = 3.696107700e-08 pk2 = -1.705647607e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.904192465e+05 lvsat = -2.997814131e-02 wvsat = -6.674427486e-02 pvsat = 1.512297528e-8
+ ua = -3.090501461e-09 lua = 6.293772985e-17 wua = 2.589929590e-16 pua = -1.058979842e-22
+ ub = 2.660073422e-18 lub = 1.531623757e-25 wub = -8.105804344e-26 pub = 6.104395078e-32
+ uc = 1.431885505e-11 luc = 1.293533702e-17 wuc = 4.461740688e-17 puc = -1.357431679e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.383850168e-03 lu0 = 3.020648534e-10 wu0 = 5.432074239e-10 pu0 = -1.328634859e-16
+ a0 = 1.1627
+ keta = -1.722141262e-02 lketa = 1.671538808e-09 wketa = 3.234598929e-09 pketa = -1.001917018e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -7.847497015e-01 lags = 3.300919954e-07 wags = 1.093168077e-06 pags = -3.463978798e-13
+ b0 = 1.939084068e-06 lb0 = -5.693953306e-13 wb0 = -7.237175015e-13 pb0 = 2.054487245e-19
+ b1 = 9.030021305e-07 lb1 = -1.328974178e-13 wb1 = 1.626298459e-13 pb1 = -1.383707119e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.792390015e-03 lpdiblc2 = 4.167843579e-09 wpdiblc2 = -4.432129831e-08 ppdiblc2 = 3.807682782e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.528726402e-01 ldelta = -2.510965531e-08 wdelta = -7.409966679e-08 pdelta = 1.649381009e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.944366650e-01 lkt1 = 5.581590322e-08 wkt1 = 1.406401783e-07 pkt1 = -4.789296051e-14
+ kt2 = 1.602871186e-01 lkt2 = -7.608269023e-08 wkt2 = -1.472278042e-07 pkt2 = 4.560381236e-14
+ at = -5.965818746e+04 lat = 3.112848044e-02 wat = 2.068174592e-01 pat = -6.967901573e-8
+ ute = -8.296308305e-01 lute = 1.912027372e-07 wute = 5.764012449e-07 pute = -1.785402856e-13
+ ua1 = 1.960985545e-09 lua1 = -3.834133652e-16 wua1 = -7.419441622e-16 pua1 = 2.298172042e-22
+ ub1 = -2.920996469e-18 lub1 = 8.327710739e-25 wub1 = 1.526088059e-24 pub1 = -4.727057762e-31
+ uc1 = -1.624596608e-10 luc1 = 5.961437994e-17 wuc1 = 1.153599358e-16 puc1 = -3.573274011e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-9.079398922e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -9.652466279e-8
+ k1 = 0.64774
+ k2 = 5.984653294e-02 wk2 = -2.739760323e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.406118400e-09 wua = 2.250849779e-16
+ ub = 3.775680869e-18 wub = -4.187879157e-25
+ uc = 5.984835477e-11 wuc = 1.298567180e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.614885955e-03 wu0 = 2.447366279e-10
+ a0 = 2.092557968e+00 wa0 = -2.209728485e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.697004740e-01 wags = -2.428104199e-7
+ b0 = 7.434122708e-07 wb0 = -3.413045763e-13
+ b1 = 4.554371000e-08 wb1 = 9.988145895e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.516110046e-03 wpdiblc2 = -6.492619474e-10
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.797151477e-03 wdelta = 2.263835451e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.911952308e-01 wkt1 = 1.298567180e-7
+ kt2 = -0.055045
+ at = 2.535045069e+05 wat = 1.720601514e-2
+ ute = -6.782284054e-01 wute = 2.351488736e-7
+ ua1 = 6.8217e-10
+ ub1 = -5.798356185e-20 wub1 = -5.523239074e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {7.436682648e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.296568591e-06 wvth0 = -1.955217254e-07 pvth0 = 1.975956620e-12
+ k1 = 0.64774
+ k2 = 1.146047477e-01 lk2 = -1.092960276e-06 wk2 = -6.021956762e-08 pk2 = 6.551182037e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.406118400e-09 wua = 2.250849779e-16
+ ub = 3.775680869e-18 wub = -4.187879157e-25
+ uc = 5.984835477e-11 wuc = 1.298567180e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.502653530e-03 lu0 = 2.240131153e-09 wu0 = 3.120085192e-10 pu0 = -1.342730133e-15
+ a0 = 1.688032644e+00 la0 = 8.074224322e-06 wa0 = 2.149882123e-08 pa0 = -4.839673910e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.697004740e-01 wags = -2.428104199e-7
+ b0 = 1.055893114e-06 lb0 = -6.237039509e-12 wb0 = -5.286049687e-13 pb0 = 3.738469008e-18
+ b1 = -1.314989892e-07 lb1 = 3.533728016e-12 wb1 = 2.060004988e-13 pb1 = -2.118109505e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 4.126891095e-03 lpdiblc2 = -5.211053704e-08 wpdiblc2 = -2.214158887e-09 ppdiblc2 = 3.123495168e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.316397107e-02 ldelta = -2.667983774e-07 wdelta = -5.748209480e-09 pdelta = 1.599184138e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.911952308e-01 wkt1 = 1.298567180e-7
+ kt2 = -0.055045
+ at = 2.141776519e+05 lat = 7.849541940e-01 wat = 4.077845337e-02 pat = -4.704999740e-7
+ ute = -6.782284054e-01 wute = 2.351488736e-7
+ ua1 = 6.8217e-10
+ ub1 = 3.138322412e-21 lub1 = -1.219977529e-24 wub1 = -9.186872592e-26 pub1 = 7.312520911e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.904819753e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.995461659e-06 wvth0 = 1.790865117e-07 pvth0 = -1.005831295e-12
+ k1 = 0.64774
+ k2 = -1.182723751e-01 lk2 = 7.606834019e-07 wk2 = 6.847586424e-08 pk2 = -3.692652600e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.472384212e-09 lua = 5.274592941e-16 wua = 2.887172452e-16 pua = -5.064969391e-22
+ ub = 4.176623365e-18 lub = -3.191402030e-24 wub = -6.773877357e-25 pub = 2.058389917e-30
+ uc = 1.060162661e-10 luc = -3.674850325e-16 wuc = -2.433535741e-17 puc = 1.947369881e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.379464306e-03 lu0 = -4.739063428e-09 wu0 = -1.679439531e-10 pu0 = 2.477571559e-15
+ a0 = 3.101515483e+00 la0 = -3.176745702e-06 wa0 = -8.052688190e-07 pa0 = 1.741189814e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.904733903e-01 lags = -9.613222203e-07 wags = -2.995009853e-07 pags = 4.512427275e-13
+ b0 = -2.577757892e-07 lb0 = 4.219436543e-12 wb0 = 2.279860855e-13 pb0 = -2.283806636e-18
+ b1 = 4.960502471e-07 lb1 = -1.461407018e-12 wb1 = -1.648702960e-13 pb1 = 8.339293037e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 2.122913568e-03 lpdiblc2 = -3.615937692e-08 wpdiblc2 = -2.581946749e-09 ppdiblc2 = 3.416245112e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.249104903e-03 ldelta = -3.267764591e-08 wdelta = 9.224240621e-09 pdelta = 4.074145412e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.028106176e+00 lkt1 = 1.089776897e-06 wkt1 = 1.941317354e-07 pkt1 = -5.116130698e-13
+ kt2 = -0.055045
+ at = 3.558881185e+05 lat = -3.430256922e-01 wat = -3.647841994e-02 pat = 1.444454234e-7
+ ute = -1.254849582e+00 lute = 4.589760407e-06 wute = 4.679315616e-07 pute = -1.852892001e-12
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.780957344e-19 lub1 = 2.226002542e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-7.710606428e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.737860487e-08 wvth0 = -8.705785916e-08 pvth0 = 4.803387746e-14
+ k1 = 0.64774
+ k2 = 8.473937114e-02 lk2 = -4.319236045e-08 wk2 = -2.846252111e-08 pk2 = 1.458651139e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.293999387e-09 lua = -1.789000171e-16 wua = 1.395986772e-16 pua = 8.397531024e-23
+ ub = 3.280303632e-18 lub = 3.578000342e-25 wub = -1.151450340e-25 pub = -1.679506205e-31
+ uc = 1.321115660e-11 wuc = 2.484375444e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.384669552e-03 lu0 = -7.999248980e-10 wu0 = 3.206826342e-10 pu0 = 5.427324301e-16
+ a0 = 2.060081615e+00 la0 = 9.470720576e-07 wa0 = -2.221858185e-07 pa0 = -5.676730972e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.760153667e-01 lags = 6.798279386e-07 wags = -1.301927493e-07 pags = -2.191755597e-13
+ b0 = 1.163634492e-06 lb0 = -1.408992819e-12 wb0 = -5.388877063e-13 pb0 = 7.528218612e-19
+ b1 = 7.628223154e-08 lb1 = 2.007693815e-13 wb1 = 7.213420299e-14 pb1 = -1.045492612e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -1.923241407e-02 lpdiblc2 = 4.840238170e-08 wpdiblc2 = 1.097319037e-08 ppdiblc2 = -1.951250309e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -5.727314582e-02 ldelta = 1.693648001e-07 wdelta = 4.133325024e-08 pdelta = -8.640219670e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.013426816e-01 lkt1 = -2.041248503e-07 wkt1 = 3.402943181e-08 pkt1 = 1.223520270e-13
+ kt2 = -0.055045
+ at = 3.056525575e+05 lat = -1.441054296e-1
+ ute = -1.499636517e-01 lute = 2.146883463e-07 wute = 3.249795199e-08 pute = -1.286837654e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-9.617921385e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -6.254765252e-8
+ k1 = 0.64774
+ k2 = 6.269964135e-02 wk2 = -2.101947409e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.385286549e-09 wua = 1.824486888e-16
+ ub = 3.462877957e-18 wub = -2.008450572e-25
+ uc = 1.321115660e-11 wuc = 2.484375444e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 9.764925405e-04 wu0 = 5.976222592e-10
+ a0 = 2.543343285e+00 wa0 = -5.118518969e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.229106026e-01 wags = -2.420312796e-7
+ b0 = 4.446689000e-07 wb0 = -1.547459223e-13
+ b1 = 1.787286566e-07 wb1 = 1.878593854e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 5.465828918e-03 wpdiblc2 = 1.016561674e-9
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.914848965e-02 wdelta = -2.755126701e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.055012989e-01 wkt1 = 9.646189871e-8
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -4.041480806e-02 wute = -3.316540579e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.140769277e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.069214026e-07 wvth0 = -1.822007469e-07 pvth0 = 1.746636045e-13
+ k1 = 0.64774
+ k2 = 1.289124583e-01 lk2 = -9.665415953e-08 wk2 = -7.279492425e-08 pk2 = 7.557921337e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.918191587e+05 lvsat = -3.912993570e-01 wvsat = -1.258264330e-01 pvsat = 1.836751356e-7
+ ua = -4.576715022e-09 lua = 1.739187714e-15 wua = 5.368132799e-16 pua = -5.172837118e-22
+ ub = 5.345945005e-18 lub = -2.748807124e-24 wub = -9.423934688e-25 pub = 1.082475294e-30
+ uc = -8.966149132e-11 luc = 1.501683478e-16 wuc = 6.535265394e-17 puc = -5.913286605e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = -2.925385563e-04 lu0 = 1.852468143e-09 wu0 = 5.972608322e-10 pu0 = 5.275930003e-19
+ a0 = 4.686504709e+00 la0 = -3.128479890e-06 wa0 = -1.369721628e-06 pa0 = 1.252275340e-12
+ keta = -7.470874428e-02 lketa = 9.069243446e-08 wketa = 3.637118399e-08 pketa = -5.309283584e-14
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -9.927243005e-01 lags = 2.504398050e-06 wags = 6.127227017e-07 pags = -1.247727124e-12
+ b0 = -8.884610589e-07 lb0 = 1.946036457e-12 wb0 = 4.305871115e-13 pb0 = -8.544398961e-19
+ b1 = -7.779787959e-07 lb1 = 1.396553704e-12 wb1 = 2.586571166e-13 pb1 = -3.501519522e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -4.715720763e-02 lpdiblc2 = 7.681647760e-08 wpdiblc2 = 1.757033173e-08 ppdiblc2 = -2.416436584e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.099183397e-02 ldelta = 1.190667812e-08 wdelta = -5.704703016e-09 pdelta = 4.305644026e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.219923876e+00 lkt1 = 6.049533576e-07 wkt1 = 2.684928215e-07 pkt1 = -2.511221396e-13
+ kt2 = 3.104333000e-03 lkt2 = -8.488348885e-8
+ at = 1.027896501e+06 lat = -1.161634747e+00 wat = -3.372071964e-01 pat = 4.922382050e-7
+ ute = -1.894130284e-01 lute = 2.175001522e-07 wute = 6.103824564e-08 pute = -1.375137802e-13
+ ua1 = 3.433807053e-10 lua1 = 5.148673930e-16 wua1 = 1.802565018e-16 pua1 = -2.631294285e-22
+ ub1 = -4.880210018e-19 lub1 = 5.344743274e-25 wub1 = 1.873271763e-25 pub1 = -2.734508456e-31
+ uc1 = -8.666613950e-11 luc1 = 1.119703274e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.591643602e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = -4.467807657e-08 wvth0 = -3.794153696e-08 pvth0 = 3.621082779e-14
+ k1 = 0.64774
+ k2 = 4.277508293e-02 lk2 = -1.398381352e-08 wk2 = 1.760886314e-09 pk2 = 4.024274178e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.645547492e+05 lvsat = -1.731823399e-01 wvsat = -2.897590342e-02 pvsat = 9.072283980e-8
+ ua = -2.778837784e-09 lua = 1.367503439e-17 wua = 8.221401961e-17 pua = -8.098207174e-23
+ ub = 2.092687198e-18 lub = 3.735070566e-25 wub = 2.599067061e-25 pub = -7.143229913e-32
+ uc = 8.813146605e-11 luc = -2.046844304e-17 wuc = -6.061143475e-18 puc = 9.406526022e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.036812071e-03 lu0 = 5.766238791e-10 wu0 = 1.051616542e-09 pu0 = -4.355402994e-16
+ a0 = 3.418373795e+00 la0 = -1.911391245e-06 wa0 = -1.172791534e-06 pa0 = 1.063271682e-12
+ keta = 4.634785522e-02 lketa = -2.549163690e-08 wketa = -3.486869307e-08 pketa = 1.527963618e-14
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.489515562e+00 lags = 1.220683421e-07 wags = -6.276299824e-07 pags = -5.729863566e-14
+ b0 = 1.664343631e-06 lb0 = -5.040178438e-13 wb0 = -7.008549878e-13 pb0 = 2.314616587e-19
+ b1 = 3.726066137e-07 lb1 = 2.922793569e-13 wb1 = 1.407663164e-13 pb1 = -2.370062567e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -9.344276432e-01 lpclm = 3.890023792e-07 wpclm = 5.781341421e-07 ppclm = -2.331672481e-13
+ pdiblc1 = 0.0
+ pdiblc2 = -1.273572964e-01 lpdiblc2 = 1.537885128e-07 wpdiblc2 = 5.707927250e-08 ppdiblc2 = -6.208307174e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.972205229e-02 ldelta = -6.365464891e-08 wdelta = -4.269320853e-08 pdelta = 3.980536220e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.563438738e-01 lkt1 = -1.278925500e-07 wkt1 = -5.429534466e-08 pkt1 = 5.867380292e-14
+ kt2 = -0.085339
+ at = -3.552405265e+05 lat = 1.658310149e-01 wat = 2.849682736e-01 pat = -1.048947024e-7
+ ute = 1.633719963e-01 lute = -1.210852753e-07 wute = -1.578646478e-07 pute = 7.257827184e-14
+ ua1 = 9.278490842e-10 lua1 = -4.607613370e-17 wua1 = -1.226842337e-16 pua1 = 2.761794239e-23
+ ub1 = 9.513846034e-19 lub1 = -8.469952022e-25 wub1 = -5.246015628e-25 pub1 = 4.098227617e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.690632801e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.054837069e-07 wvth0 = -6.621772801e-08 pvth0 = 4.921080662e-14
+ k1 = 0.64774
+ k2 = 6.313987534e-02 lk2 = -2.334652683e-08 wk2 = -3.231014780e-08 pk2 = 1.968843211e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -6.617423650e+05 lvsat = 2.067077584e-01 wvsat = 4.440396907e-01 pvsat = -1.267460796e-7
+ ua = -2.061790088e-09 lua = -3.159876438e-16 wua = -3.576145801e-16 pua = 1.212291270e-22
+ ub = 1.317011342e-18 lub = 7.301240316e-25 wub = 7.239706815e-25 pub = -2.847857118e-31
+ uc = 7.453845146e-11 luc = -1.421905458e-17 wuc = 8.521901228e-18 puc = 2.701971220e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.699113389e-03 lu0 = 2.721308479e-10 wu0 = 3.542392793e-10 pu0 = -1.149211029e-16
+ a0 = -7.390840508e-01 wa0 = 1.139925556e-6
+ keta = -9.098880846e-03 wketa = -1.634030369e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.240346405e+00 lags = -1.142626138e-06 wags = -1.918864479e-06 pags = 5.363464239e-13
+ b0 = 1.741094271e-06 lb0 = -5.393039504e-13 wb0 = -6.050428131e-13 pb0 = 1.874120114e-19
+ b1 = 3.090568317e-06 lb1 = -9.573035363e-13 wb1 = -1.148592951e-12 pb1 = 3.557766667e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.831045088e-02 wpclm = 7.097318924e-8
+ pdiblc1 = 0.0
+ pdiblc2 = -4.564133840e-02 lpdiblc2 = 1.162196011e-07 wpdiblc2 = -1.469082037e-08 ppdiblc2 = -2.908677155e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.249506561e-01 ldelta = -7.525349952e-08 wdelta = -5.736328537e-08 pdelta = 4.654993002e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.347495730e-01 lkt1 = 9.205447025e-08 wkt1 = 2.247434548e-07 pkt1 = -6.961428511e-14
+ kt2 = -0.085339
+ at = -5.123944135e+03 lat = 4.864916196e-03 wat = 1.741297428e-01 pat = -5.393668784e-8
+ ute = 1.320027500e-01 lute = -1.066632643e-07 pute = 2.524354897e-29
+ ua1 = 1.043337168e-09 lua1 = -9.917178040e-17 wua1 = -1.919075604e-16 pua1 = 5.944336683e-23
+ ub1 = -2.250590322e-18 lub1 = 6.251127698e-25 wub1 = 1.124247955e-24 pub1 = -3.482358040e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8_lvt
