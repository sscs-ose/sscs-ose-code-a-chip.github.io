# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p84L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p84L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  2.860000 BY  1.950000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.705600 ;
    PORT
      LAYER met3 ;
        RECT 0.585000 0.205000 0.915000 0.645000 ;
        RECT 0.585000 0.645000 2.635000 0.975000 ;
        RECT 1.445000 0.205000 1.775000 0.645000 ;
        RECT 2.305000 0.205000 2.635000 0.645000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.756000 ;
    PORT
      LAYER met1 ;
        RECT 0.565000 1.195000 2.655000 1.485000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.940800 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 3.015000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  0.945000 ;
        RECT 1.065000 -0.145000 1.295000  0.945000 ;
        RECT 1.925000 -0.145000 2.155000  0.945000 ;
        RECT 2.785000 -0.145000 3.015000  0.945000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.365000 1.050000 0.445000 1.125000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.255000 0.405000 0.945000 ;
      RECT 0.595000 1.175000 2.625000 1.505000 ;
      RECT 0.665000 0.255000 0.835000 0.945000 ;
      RECT 1.095000 0.255000 1.265000 0.945000 ;
      RECT 1.525000 0.255000 1.695000 0.945000 ;
      RECT 1.955000 0.255000 2.125000 0.945000 ;
      RECT 2.385000 0.255000 2.555000 0.945000 ;
      RECT 2.815000 0.255000 2.985000 0.945000 ;
    LAYER mcon ;
      RECT 0.235000 0.335000 0.405000 0.505000 ;
      RECT 0.235000 0.695000 0.405000 0.865000 ;
      RECT 0.625000 1.255000 0.795000 1.425000 ;
      RECT 0.665000 0.335000 0.835000 0.505000 ;
      RECT 0.665000 0.695000 0.835000 0.865000 ;
      RECT 0.985000 1.255000 1.155000 1.425000 ;
      RECT 1.095000 0.335000 1.265000 0.505000 ;
      RECT 1.095000 0.695000 1.265000 0.865000 ;
      RECT 1.345000 1.255000 1.515000 1.425000 ;
      RECT 1.525000 0.335000 1.695000 0.505000 ;
      RECT 1.525000 0.695000 1.695000 0.865000 ;
      RECT 1.705000 1.255000 1.875000 1.425000 ;
      RECT 1.955000 0.335000 2.125000 0.505000 ;
      RECT 1.955000 0.695000 2.125000 0.865000 ;
      RECT 2.065000 1.255000 2.235000 1.425000 ;
      RECT 2.385000 0.335000 2.555000 0.505000 ;
      RECT 2.385000 0.695000 2.555000 0.865000 ;
      RECT 2.425000 1.255000 2.595000 1.425000 ;
      RECT 2.815000 0.335000 2.985000 0.505000 ;
      RECT 2.815000 0.695000 2.985000 0.865000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 0.945000 ;
      RECT 1.480000 0.255000 1.740000 0.945000 ;
      RECT 2.340000 0.255000 2.600000 0.945000 ;
    LAYER met2 ;
      RECT 0.585000 0.205000 0.915000 0.975000 ;
      RECT 1.445000 0.205000 1.775000 0.975000 ;
      RECT 2.305000 0.205000 2.635000 0.975000 ;
    LAYER via ;
      RECT 0.620000 0.300000 0.880000 0.560000 ;
      RECT 0.620000 0.620000 0.880000 0.880000 ;
      RECT 1.480000 0.300000 1.740000 0.560000 ;
      RECT 1.480000 0.620000 1.740000 0.880000 ;
      RECT 2.340000 0.300000 2.600000 0.560000 ;
      RECT 2.340000 0.620000 2.600000 0.880000 ;
    LAYER via2 ;
      RECT 0.610000 0.250000 0.890000 0.530000 ;
      RECT 0.610000 0.650000 0.890000 0.930000 ;
      RECT 1.470000 0.250000 1.750000 0.530000 ;
      RECT 1.470000 0.650000 1.750000 0.930000 ;
      RECT 2.330000 0.250000 2.610000 0.530000 ;
      RECT 2.330000 0.650000 2.610000 0.930000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p84L0p15
END LIBRARY
