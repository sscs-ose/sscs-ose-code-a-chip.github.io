# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_20v0_zvt_withptap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_20v0_zvt_withptap ;
  ORIGIN  9.200000  4.910000 ;
  SIZE  19.15000 BY  39.82000 ;
  PIN D
    ANTENNADIFFAREA  22.50000 ;
    PORT
      LAYER met1 ;
        RECT -1.375000 -1.000000 2.125000 31.000000 ;
    END
  END D
  PIN PSUB
    ANTENNADIFFAREA  47.682999 ;
    PORT
      LAYER li1 ;
        RECT -9.200000 -4.910000  9.950000 -4.500000 ;
        RECT -9.200000 -4.500000 -8.790000 34.500000 ;
        RECT -9.200000 34.500000  9.950000 34.910000 ;
        RECT  9.540000 -4.500000  9.950000 34.500000 ;
    END
  END PSUB
  PIN S
    ANTENNADIFFAREA  8.700000 ;
    PORT
      LAYER met1 ;
        RECT -8.560000 -1.000000 -5.560000 31.000000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.310000 -1.000000 9.310000 31.000000 ;
    END
  END S
  OBS
    LAYER li1 ;
      RECT -8.310000  0.045000 -7.980000 29.955000 ;
      RECT -1.480000 -3.285000  2.300000 -2.215000 ;
      RECT -0.125000 -0.250000  0.875000 30.250000 ;
      RECT  8.730000  0.045000  9.060000 29.955000 ;
    LAYER mcon ;
      RECT -8.230000  0.155000 -8.060000  0.325000 ;
      RECT -8.230000  0.515000 -8.060000  0.685000 ;
      RECT -8.230000  0.875000 -8.060000  1.045000 ;
      RECT -8.230000  1.235000 -8.060000  1.405000 ;
      RECT -8.230000  1.595000 -8.060000  1.765000 ;
      RECT -8.230000  1.955000 -8.060000  2.125000 ;
      RECT -8.230000  2.315000 -8.060000  2.485000 ;
      RECT -8.230000  2.675000 -8.060000  2.845000 ;
      RECT -8.230000  3.035000 -8.060000  3.205000 ;
      RECT -8.230000  3.395000 -8.060000  3.565000 ;
      RECT -8.230000  3.755000 -8.060000  3.925000 ;
      RECT -8.230000  4.115000 -8.060000  4.285000 ;
      RECT -8.230000  4.475000 -8.060000  4.645000 ;
      RECT -8.230000  4.835000 -8.060000  5.005000 ;
      RECT -8.230000  5.195000 -8.060000  5.365000 ;
      RECT -8.230000  5.555000 -8.060000  5.725000 ;
      RECT -8.230000  5.915000 -8.060000  6.085000 ;
      RECT -8.230000  6.275000 -8.060000  6.445000 ;
      RECT -8.230000  6.635000 -8.060000  6.805000 ;
      RECT -8.230000  6.995000 -8.060000  7.165000 ;
      RECT -8.230000  7.355000 -8.060000  7.525000 ;
      RECT -8.230000  7.715000 -8.060000  7.885000 ;
      RECT -8.230000  8.075000 -8.060000  8.245000 ;
      RECT -8.230000  8.435000 -8.060000  8.605000 ;
      RECT -8.230000  8.795000 -8.060000  8.965000 ;
      RECT -8.230000  9.155000 -8.060000  9.325000 ;
      RECT -8.230000  9.515000 -8.060000  9.685000 ;
      RECT -8.230000  9.875000 -8.060000 10.045000 ;
      RECT -8.230000 10.235000 -8.060000 10.405000 ;
      RECT -8.230000 10.595000 -8.060000 10.765000 ;
      RECT -8.230000 10.955000 -8.060000 11.125000 ;
      RECT -8.230000 11.315000 -8.060000 11.485000 ;
      RECT -8.230000 11.675000 -8.060000 11.845000 ;
      RECT -8.230000 12.035000 -8.060000 12.205000 ;
      RECT -8.230000 12.395000 -8.060000 12.565000 ;
      RECT -8.230000 12.755000 -8.060000 12.925000 ;
      RECT -8.230000 13.115000 -8.060000 13.285000 ;
      RECT -8.230000 13.475000 -8.060000 13.645000 ;
      RECT -8.230000 13.835000 -8.060000 14.005000 ;
      RECT -8.230000 14.195000 -8.060000 14.365000 ;
      RECT -8.230000 14.555000 -8.060000 14.725000 ;
      RECT -8.230000 14.915000 -8.060000 15.085000 ;
      RECT -8.230000 15.275000 -8.060000 15.445000 ;
      RECT -8.230000 15.635000 -8.060000 15.805000 ;
      RECT -8.230000 15.995000 -8.060000 16.165000 ;
      RECT -8.230000 16.355000 -8.060000 16.525000 ;
      RECT -8.230000 16.715000 -8.060000 16.885000 ;
      RECT -8.230000 17.075000 -8.060000 17.245000 ;
      RECT -8.230000 17.435000 -8.060000 17.605000 ;
      RECT -8.230000 17.795000 -8.060000 17.965000 ;
      RECT -8.230000 18.155000 -8.060000 18.325000 ;
      RECT -8.230000 18.515000 -8.060000 18.685000 ;
      RECT -8.230000 18.875000 -8.060000 19.045000 ;
      RECT -8.230000 19.235000 -8.060000 19.405000 ;
      RECT -8.230000 19.595000 -8.060000 19.765000 ;
      RECT -8.230000 19.955000 -8.060000 20.125000 ;
      RECT -8.230000 20.315000 -8.060000 20.485000 ;
      RECT -8.230000 20.675000 -8.060000 20.845000 ;
      RECT -8.230000 21.035000 -8.060000 21.205000 ;
      RECT -8.230000 21.395000 -8.060000 21.565000 ;
      RECT -8.230000 21.755000 -8.060000 21.925000 ;
      RECT -8.230000 22.115000 -8.060000 22.285000 ;
      RECT -8.230000 22.475000 -8.060000 22.645000 ;
      RECT -8.230000 22.835000 -8.060000 23.005000 ;
      RECT -8.230000 23.195000 -8.060000 23.365000 ;
      RECT -8.230000 23.555000 -8.060000 23.725000 ;
      RECT -8.230000 23.915000 -8.060000 24.085000 ;
      RECT -8.230000 24.275000 -8.060000 24.445000 ;
      RECT -8.230000 24.635000 -8.060000 24.805000 ;
      RECT -8.230000 24.995000 -8.060000 25.165000 ;
      RECT -8.230000 25.355000 -8.060000 25.525000 ;
      RECT -8.230000 25.715000 -8.060000 25.885000 ;
      RECT -8.230000 26.075000 -8.060000 26.245000 ;
      RECT -8.230000 26.435000 -8.060000 26.605000 ;
      RECT -8.230000 26.795000 -8.060000 26.965000 ;
      RECT -8.230000 27.155000 -8.060000 27.325000 ;
      RECT -8.230000 27.515000 -8.060000 27.685000 ;
      RECT -8.230000 27.875000 -8.060000 28.045000 ;
      RECT -8.230000 28.235000 -8.060000 28.405000 ;
      RECT -8.230000 28.595000 -8.060000 28.765000 ;
      RECT -8.230000 28.955000 -8.060000 29.125000 ;
      RECT -8.230000 29.315000 -8.060000 29.485000 ;
      RECT -8.230000 29.675000 -8.060000 29.845000 ;
      RECT -1.400000 -3.205000 -1.230000 -3.035000 ;
      RECT -1.400000 -2.835000 -1.230000 -2.665000 ;
      RECT -1.400000 -2.465000 -1.230000 -2.295000 ;
      RECT -1.030000 -3.205000 -0.860000 -3.035000 ;
      RECT -1.030000 -2.835000 -0.860000 -2.665000 ;
      RECT -1.030000 -2.465000 -0.860000 -2.295000 ;
      RECT -0.660000 -3.205000 -0.490000 -3.035000 ;
      RECT -0.660000 -2.835000 -0.490000 -2.665000 ;
      RECT -0.660000 -2.465000 -0.490000 -2.295000 ;
      RECT -0.290000 -3.205000 -0.120000 -3.035000 ;
      RECT -0.290000 -2.835000 -0.120000 -2.665000 ;
      RECT -0.290000 -2.465000 -0.120000 -2.295000 ;
      RECT  0.080000 -3.205000  0.250000 -3.035000 ;
      RECT  0.080000 -2.835000  0.250000 -2.665000 ;
      RECT  0.080000 -2.465000  0.250000 -2.295000 ;
      RECT  0.110000  0.155000  0.640000 29.845000 ;
      RECT  0.450000 -3.205000  0.620000 -3.035000 ;
      RECT  0.450000 -2.835000  0.620000 -2.665000 ;
      RECT  0.450000 -2.465000  0.620000 -2.295000 ;
      RECT  0.820000 -3.205000  0.990000 -3.035000 ;
      RECT  0.820000 -2.835000  0.990000 -2.665000 ;
      RECT  0.820000 -2.465000  0.990000 -2.295000 ;
      RECT  1.190000 -3.205000  1.360000 -3.035000 ;
      RECT  1.190000 -2.835000  1.360000 -2.665000 ;
      RECT  1.190000 -2.465000  1.360000 -2.295000 ;
      RECT  1.560000 -3.205000  1.730000 -3.035000 ;
      RECT  1.560000 -2.835000  1.730000 -2.665000 ;
      RECT  1.560000 -2.465000  1.730000 -2.295000 ;
      RECT  1.930000 -3.205000  2.100000 -3.035000 ;
      RECT  1.930000 -2.835000  2.100000 -2.665000 ;
      RECT  1.930000 -2.465000  2.100000 -2.295000 ;
      RECT  8.810000  0.155000  8.980000  0.325000 ;
      RECT  8.810000  0.515000  8.980000  0.685000 ;
      RECT  8.810000  0.875000  8.980000  1.045000 ;
      RECT  8.810000  1.235000  8.980000  1.405000 ;
      RECT  8.810000  1.595000  8.980000  1.765000 ;
      RECT  8.810000  1.955000  8.980000  2.125000 ;
      RECT  8.810000  2.315000  8.980000  2.485000 ;
      RECT  8.810000  2.675000  8.980000  2.845000 ;
      RECT  8.810000  3.035000  8.980000  3.205000 ;
      RECT  8.810000  3.395000  8.980000  3.565000 ;
      RECT  8.810000  3.755000  8.980000  3.925000 ;
      RECT  8.810000  4.115000  8.980000  4.285000 ;
      RECT  8.810000  4.475000  8.980000  4.645000 ;
      RECT  8.810000  4.835000  8.980000  5.005000 ;
      RECT  8.810000  5.195000  8.980000  5.365000 ;
      RECT  8.810000  5.555000  8.980000  5.725000 ;
      RECT  8.810000  5.915000  8.980000  6.085000 ;
      RECT  8.810000  6.275000  8.980000  6.445000 ;
      RECT  8.810000  6.635000  8.980000  6.805000 ;
      RECT  8.810000  6.995000  8.980000  7.165000 ;
      RECT  8.810000  7.355000  8.980000  7.525000 ;
      RECT  8.810000  7.715000  8.980000  7.885000 ;
      RECT  8.810000  8.075000  8.980000  8.245000 ;
      RECT  8.810000  8.435000  8.980000  8.605000 ;
      RECT  8.810000  8.795000  8.980000  8.965000 ;
      RECT  8.810000  9.155000  8.980000  9.325000 ;
      RECT  8.810000  9.515000  8.980000  9.685000 ;
      RECT  8.810000  9.875000  8.980000 10.045000 ;
      RECT  8.810000 10.235000  8.980000 10.405000 ;
      RECT  8.810000 10.595000  8.980000 10.765000 ;
      RECT  8.810000 10.955000  8.980000 11.125000 ;
      RECT  8.810000 11.315000  8.980000 11.485000 ;
      RECT  8.810000 11.675000  8.980000 11.845000 ;
      RECT  8.810000 12.035000  8.980000 12.205000 ;
      RECT  8.810000 12.395000  8.980000 12.565000 ;
      RECT  8.810000 12.755000  8.980000 12.925000 ;
      RECT  8.810000 13.115000  8.980000 13.285000 ;
      RECT  8.810000 13.475000  8.980000 13.645000 ;
      RECT  8.810000 13.835000  8.980000 14.005000 ;
      RECT  8.810000 14.195000  8.980000 14.365000 ;
      RECT  8.810000 14.555000  8.980000 14.725000 ;
      RECT  8.810000 14.915000  8.980000 15.085000 ;
      RECT  8.810000 15.275000  8.980000 15.445000 ;
      RECT  8.810000 15.635000  8.980000 15.805000 ;
      RECT  8.810000 15.995000  8.980000 16.165000 ;
      RECT  8.810000 16.355000  8.980000 16.525000 ;
      RECT  8.810000 16.715000  8.980000 16.885000 ;
      RECT  8.810000 17.075000  8.980000 17.245000 ;
      RECT  8.810000 17.435000  8.980000 17.605000 ;
      RECT  8.810000 17.795000  8.980000 17.965000 ;
      RECT  8.810000 18.155000  8.980000 18.325000 ;
      RECT  8.810000 18.515000  8.980000 18.685000 ;
      RECT  8.810000 18.875000  8.980000 19.045000 ;
      RECT  8.810000 19.235000  8.980000 19.405000 ;
      RECT  8.810000 19.595000  8.980000 19.765000 ;
      RECT  8.810000 19.955000  8.980000 20.125000 ;
      RECT  8.810000 20.315000  8.980000 20.485000 ;
      RECT  8.810000 20.675000  8.980000 20.845000 ;
      RECT  8.810000 21.035000  8.980000 21.205000 ;
      RECT  8.810000 21.395000  8.980000 21.565000 ;
      RECT  8.810000 21.755000  8.980000 21.925000 ;
      RECT  8.810000 22.115000  8.980000 22.285000 ;
      RECT  8.810000 22.475000  8.980000 22.645000 ;
      RECT  8.810000 22.835000  8.980000 23.005000 ;
      RECT  8.810000 23.195000  8.980000 23.365000 ;
      RECT  8.810000 23.555000  8.980000 23.725000 ;
      RECT  8.810000 23.915000  8.980000 24.085000 ;
      RECT  8.810000 24.275000  8.980000 24.445000 ;
      RECT  8.810000 24.635000  8.980000 24.805000 ;
      RECT  8.810000 24.995000  8.980000 25.165000 ;
      RECT  8.810000 25.355000  8.980000 25.525000 ;
      RECT  8.810000 25.715000  8.980000 25.885000 ;
      RECT  8.810000 26.075000  8.980000 26.245000 ;
      RECT  8.810000 26.435000  8.980000 26.605000 ;
      RECT  8.810000 26.795000  8.980000 26.965000 ;
      RECT  8.810000 27.155000  8.980000 27.325000 ;
      RECT  8.810000 27.515000  8.980000 27.685000 ;
      RECT  8.810000 27.875000  8.980000 28.045000 ;
      RECT  8.810000 28.235000  8.980000 28.405000 ;
      RECT  8.810000 28.595000  8.980000 28.765000 ;
      RECT  8.810000 28.955000  8.980000 29.125000 ;
      RECT  8.810000 29.315000  8.980000 29.485000 ;
      RECT  8.810000 29.675000  8.980000 29.845000 ;
    LAYER met1 ;
      RECT -1.480000 -3.285000 2.300000 -2.215000 ;
    LAYER met2 ;
      RECT -1.480000 -3.285000 2.300000 -2.215000 ;
    LAYER via ;
      RECT -1.445000 -3.250000 -1.185000 -2.990000 ;
      RECT -1.445000 -2.880000 -1.185000 -2.620000 ;
      RECT -1.445000 -2.510000 -1.185000 -2.250000 ;
      RECT -1.075000 -3.250000 -0.815000 -2.990000 ;
      RECT -1.075000 -2.880000 -0.815000 -2.620000 ;
      RECT -1.075000 -2.510000 -0.815000 -2.250000 ;
      RECT -0.705000 -3.250000 -0.445000 -2.990000 ;
      RECT -0.705000 -2.880000 -0.445000 -2.620000 ;
      RECT -0.705000 -2.510000 -0.445000 -2.250000 ;
      RECT -0.335000 -3.250000 -0.075000 -2.990000 ;
      RECT -0.335000 -2.880000 -0.075000 -2.620000 ;
      RECT -0.335000 -2.510000 -0.075000 -2.250000 ;
      RECT  0.035000 -3.250000  0.295000 -2.990000 ;
      RECT  0.035000 -2.880000  0.295000 -2.620000 ;
      RECT  0.035000 -2.510000  0.295000 -2.250000 ;
      RECT  0.405000 -3.250000  0.665000 -2.990000 ;
      RECT  0.405000 -2.880000  0.665000 -2.620000 ;
      RECT  0.405000 -2.510000  0.665000 -2.250000 ;
      RECT  0.775000 -3.250000  1.035000 -2.990000 ;
      RECT  0.775000 -2.880000  1.035000 -2.620000 ;
      RECT  0.775000 -2.510000  1.035000 -2.250000 ;
      RECT  1.145000 -3.250000  1.405000 -2.990000 ;
      RECT  1.145000 -2.880000  1.405000 -2.620000 ;
      RECT  1.145000 -2.510000  1.405000 -2.250000 ;
      RECT  1.515000 -3.250000  1.775000 -2.990000 ;
      RECT  1.515000 -2.880000  1.775000 -2.620000 ;
      RECT  1.515000 -2.510000  1.775000 -2.250000 ;
      RECT  1.885000 -3.250000  2.145000 -2.990000 ;
      RECT  1.885000 -2.880000  2.145000 -2.620000 ;
      RECT  1.885000 -2.510000  2.145000 -2.250000 ;
  END
END sky130_fd_pr__rf_nfet_20v0_zvt_withptap
END LIBRARY
