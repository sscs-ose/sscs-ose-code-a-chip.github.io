# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18 ;
  ORIGIN -0.050000 -0.050000 ;
  SIZE  3.500000 BY  2.570000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 1.460000 3.550000 2.100000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.188000 ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.150000 2.645000 0.320000 ;
        RECT 0.955000 2.350000 2.645000 2.520000 ;
      LAYER mcon ;
        RECT 0.995000 0.150000 1.165000 0.320000 ;
        RECT 0.995000 2.350000 1.165000 2.520000 ;
        RECT 1.355000 0.150000 1.525000 0.320000 ;
        RECT 1.355000 2.350000 1.525000 2.520000 ;
        RECT 1.715000 0.150000 1.885000 0.320000 ;
        RECT 1.715000 2.350000 1.885000 2.520000 ;
        RECT 2.075000 0.150000 2.245000 0.320000 ;
        RECT 2.075000 2.350000 2.245000 2.520000 ;
        RECT 2.435000 0.150000 2.605000 0.320000 ;
        RECT 2.435000 2.350000 2.605000 2.520000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.935000 0.050000 2.665000 0.380000 ;
        RECT 0.935000 2.290000 2.665000 2.620000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.570000 3.550000 1.210000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.478500 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.570000 0.470000 2.100000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.130000 0.570000 3.420000 2.100000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.660000 0.410000 2.010000 ;
      RECT 0.795000 0.490000 0.965000 2.180000 ;
      RECT 1.255000 0.490000 1.425000 2.180000 ;
      RECT 1.715000 0.490000 1.885000 2.180000 ;
      RECT 2.175000 0.490000 2.345000 2.180000 ;
      RECT 2.635000 0.490000 2.805000 2.180000 ;
      RECT 3.190000 0.660000 3.360000 2.010000 ;
    LAYER mcon ;
      RECT 0.240000 0.710000 0.410000 0.880000 ;
      RECT 0.240000 1.070000 0.410000 1.240000 ;
      RECT 0.240000 1.430000 0.410000 1.600000 ;
      RECT 0.240000 1.790000 0.410000 1.960000 ;
      RECT 0.795000 0.710000 0.965000 0.880000 ;
      RECT 0.795000 1.070000 0.965000 1.240000 ;
      RECT 0.795000 1.430000 0.965000 1.600000 ;
      RECT 0.795000 1.790000 0.965000 1.960000 ;
      RECT 1.255000 0.710000 1.425000 0.880000 ;
      RECT 1.255000 1.070000 1.425000 1.240000 ;
      RECT 1.255000 1.430000 1.425000 1.600000 ;
      RECT 1.255000 1.790000 1.425000 1.960000 ;
      RECT 1.715000 0.710000 1.885000 0.880000 ;
      RECT 1.715000 1.070000 1.885000 1.240000 ;
      RECT 1.715000 1.430000 1.885000 1.600000 ;
      RECT 1.715000 1.790000 1.885000 1.960000 ;
      RECT 2.175000 0.710000 2.345000 0.880000 ;
      RECT 2.175000 1.070000 2.345000 1.240000 ;
      RECT 2.175000 1.430000 2.345000 1.600000 ;
      RECT 2.175000 1.790000 2.345000 1.960000 ;
      RECT 2.635000 0.710000 2.805000 0.880000 ;
      RECT 2.635000 1.070000 2.805000 1.240000 ;
      RECT 2.635000 1.430000 2.805000 1.600000 ;
      RECT 2.635000 1.790000 2.805000 1.960000 ;
      RECT 3.190000 0.710000 3.360000 0.880000 ;
      RECT 3.190000 1.070000 3.360000 1.240000 ;
      RECT 3.190000 1.430000 3.360000 1.600000 ;
      RECT 3.190000 1.790000 3.360000 1.960000 ;
    LAYER met1 ;
      RECT 0.750000 0.570000 1.010000 2.100000 ;
      RECT 1.210000 0.570000 1.470000 2.100000 ;
      RECT 1.670000 0.570000 1.930000 2.100000 ;
      RECT 2.130000 0.570000 2.390000 2.100000 ;
      RECT 2.590000 0.570000 2.850000 2.100000 ;
    LAYER via ;
      RECT 0.750000 0.600000 1.010000 0.860000 ;
      RECT 0.750000 0.920000 1.010000 1.180000 ;
      RECT 1.210000 1.490000 1.470000 1.750000 ;
      RECT 1.210000 1.810000 1.470000 2.070000 ;
      RECT 1.670000 0.600000 1.930000 0.860000 ;
      RECT 1.670000 0.920000 1.930000 1.180000 ;
      RECT 2.130000 1.490000 2.390000 1.750000 ;
      RECT 2.130000 1.810000 2.390000 2.070000 ;
      RECT 2.590000 0.600000 2.850000 0.860000 ;
      RECT 2.590000 0.920000 2.850000 1.180000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18
END LIBRARY
