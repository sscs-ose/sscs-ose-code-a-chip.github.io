magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -276 -2137 276 2137
<< nmos >>
rect -80 1127 80 1927
rect -80 109 80 909
rect -80 -909 80 -109
rect -80 -1927 80 -1127
<< ndiff >>
rect -138 1915 -80 1927
rect -138 1139 -126 1915
rect -92 1139 -80 1915
rect -138 1127 -80 1139
rect 80 1915 138 1927
rect 80 1139 92 1915
rect 126 1139 138 1915
rect 80 1127 138 1139
rect -138 897 -80 909
rect -138 121 -126 897
rect -92 121 -80 897
rect -138 109 -80 121
rect 80 897 138 909
rect 80 121 92 897
rect 126 121 138 897
rect 80 109 138 121
rect -138 -121 -80 -109
rect -138 -897 -126 -121
rect -92 -897 -80 -121
rect -138 -909 -80 -897
rect 80 -121 138 -109
rect 80 -897 92 -121
rect 126 -897 138 -121
rect 80 -909 138 -897
rect -138 -1139 -80 -1127
rect -138 -1915 -126 -1139
rect -92 -1915 -80 -1139
rect -138 -1927 -80 -1915
rect 80 -1139 138 -1127
rect 80 -1915 92 -1139
rect 126 -1915 138 -1139
rect 80 -1927 138 -1915
<< ndiffc >>
rect -126 1139 -92 1915
rect 92 1139 126 1915
rect -126 121 -92 897
rect 92 121 126 897
rect -126 -897 -92 -121
rect 92 -897 126 -121
rect -126 -1915 -92 -1139
rect 92 -1915 126 -1139
<< psubdiff >>
rect -240 2067 -144 2101
rect 144 2067 240 2101
rect -240 2005 -206 2067
rect 206 2005 240 2067
rect -240 -2067 -206 -2005
rect 206 -2067 240 -2005
rect -240 -2101 -144 -2067
rect 144 -2101 240 -2067
<< psubdiffcont >>
rect -144 2067 144 2101
rect -240 -2005 -206 2005
rect 206 -2005 240 2005
rect -144 -2101 144 -2067
<< poly >>
rect -80 1999 80 2015
rect -80 1965 -64 1999
rect 64 1965 80 1999
rect -80 1927 80 1965
rect -80 1089 80 1127
rect -80 1055 -64 1089
rect 64 1055 80 1089
rect -80 1039 80 1055
rect -80 981 80 997
rect -80 947 -64 981
rect 64 947 80 981
rect -80 909 80 947
rect -80 71 80 109
rect -80 37 -64 71
rect 64 37 80 71
rect -80 21 80 37
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -109 80 -71
rect -80 -947 80 -909
rect -80 -981 -64 -947
rect 64 -981 80 -947
rect -80 -997 80 -981
rect -80 -1055 80 -1039
rect -80 -1089 -64 -1055
rect 64 -1089 80 -1055
rect -80 -1127 80 -1089
rect -80 -1965 80 -1927
rect -80 -1999 -64 -1965
rect 64 -1999 80 -1965
rect -80 -2015 80 -1999
<< polycont >>
rect -64 1965 64 1999
rect -64 1055 64 1089
rect -64 947 64 981
rect -64 37 64 71
rect -64 -71 64 -37
rect -64 -981 64 -947
rect -64 -1089 64 -1055
rect -64 -1999 64 -1965
<< locali >>
rect -240 2067 -144 2101
rect 144 2067 240 2101
rect -240 2005 -206 2067
rect 206 2005 240 2067
rect -80 1965 -64 1999
rect 64 1965 80 1999
rect -126 1915 -92 1931
rect -126 1123 -92 1139
rect 92 1915 126 1931
rect 92 1123 126 1139
rect -80 1055 -64 1089
rect 64 1055 80 1089
rect -80 947 -64 981
rect 64 947 80 981
rect -126 897 -92 913
rect -126 105 -92 121
rect 92 897 126 913
rect 92 105 126 121
rect -80 37 -64 71
rect 64 37 80 71
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -121 -92 -105
rect -126 -913 -92 -897
rect 92 -121 126 -105
rect 92 -913 126 -897
rect -80 -981 -64 -947
rect 64 -981 80 -947
rect -80 -1089 -64 -1055
rect 64 -1089 80 -1055
rect -126 -1139 -92 -1123
rect -126 -1931 -92 -1915
rect 92 -1139 126 -1123
rect 92 -1931 126 -1915
rect -80 -1999 -64 -1965
rect 64 -1999 80 -1965
rect -240 -2067 -206 -2005
rect 206 -2067 240 -2005
rect -240 -2101 -144 -2067
rect 144 -2101 240 -2067
<< viali >>
rect -64 1965 64 1999
rect -126 1139 -92 1915
rect 92 1139 126 1915
rect -64 1055 64 1089
rect -64 947 64 981
rect -126 121 -92 897
rect 92 121 126 897
rect -64 37 64 71
rect -64 -71 64 -37
rect -126 -897 -92 -121
rect 92 -897 126 -121
rect -64 -981 64 -947
rect -64 -1089 64 -1055
rect -126 -1915 -92 -1139
rect 92 -1915 126 -1139
rect -64 -1999 64 -1965
<< metal1 >>
rect -76 1999 76 2005
rect -76 1965 -64 1999
rect 64 1965 76 1999
rect -76 1959 76 1965
rect -132 1915 -86 1927
rect -132 1139 -126 1915
rect -92 1139 -86 1915
rect -132 1127 -86 1139
rect 86 1915 132 1927
rect 86 1139 92 1915
rect 126 1139 132 1915
rect 86 1127 132 1139
rect -76 1089 76 1095
rect -76 1055 -64 1089
rect 64 1055 76 1089
rect -76 1049 76 1055
rect -76 981 76 987
rect -76 947 -64 981
rect 64 947 76 981
rect -76 941 76 947
rect -132 897 -86 909
rect -132 121 -126 897
rect -92 121 -86 897
rect -132 109 -86 121
rect 86 897 132 909
rect 86 121 92 897
rect 126 121 132 897
rect 86 109 132 121
rect -76 71 76 77
rect -76 37 -64 71
rect 64 37 76 71
rect -76 31 76 37
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -121 -86 -109
rect -132 -897 -126 -121
rect -92 -897 -86 -121
rect -132 -909 -86 -897
rect 86 -121 132 -109
rect 86 -897 92 -121
rect 126 -897 132 -121
rect 86 -909 132 -897
rect -76 -947 76 -941
rect -76 -981 -64 -947
rect 64 -981 76 -947
rect -76 -987 76 -981
rect -76 -1055 76 -1049
rect -76 -1089 -64 -1055
rect 64 -1089 76 -1055
rect -76 -1095 76 -1089
rect -132 -1139 -86 -1127
rect -132 -1915 -126 -1139
rect -92 -1915 -86 -1139
rect -132 -1927 -86 -1915
rect 86 -1139 132 -1127
rect 86 -1915 92 -1139
rect 126 -1915 132 -1139
rect 86 -1927 132 -1915
rect -76 -1965 76 -1959
rect -76 -1999 -64 -1965
rect 64 -1999 76 -1965
rect -76 -2005 76 -1999
<< labels >>
rlabel psubdiffcont 0 -2084 0 -2084 0 B
port 1 nsew
rlabel ndiffc -109 -1527 -109 -1527 0 D0
port 2 nsew
rlabel ndiffc 109 -1527 109 -1527 0 S0
port 3 nsew
rlabel polycont 0 -1072 0 -1072 0 G0
port 4 nsew
rlabel ndiffc -109 -509 -109 -509 0 D1
port 5 nsew
rlabel ndiffc 109 -509 109 -509 0 S1
port 6 nsew
rlabel polycont 0 -54 0 -54 0 G1
port 7 nsew
rlabel ndiffc -109 509 -109 509 0 D2
port 8 nsew
rlabel ndiffc 109 509 109 509 0 S2
port 9 nsew
rlabel polycont 0 964 0 964 0 G2
port 10 nsew
rlabel ndiffc -109 1527 -109 1527 0 D3
port 11 nsew
rlabel ndiffc 109 1527 109 1527 0 S3
port 12 nsew
rlabel polycont 0 1982 0 1982 0 G3
port 13 nsew
<< properties >>
string FIXED_BBOX -223 -2084 223 2084
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.8 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 4
<< end >>
