# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 ;
  ORIGIN  0.000000  0.485000 ;
  SIZE  1.470000 BY  6.155000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.400000 ;
    PORT
      LAYER met2 ;
        RECT 0.605000 4.520000 0.865000 5.160000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.500000 ;
    PORT
      LAYER met1 ;
        RECT 0.410000 5.360000 1.060000 5.650000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.650000 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.485000 1.280000 -0.225000 ;
        RECT 0.190000 -0.225000 0.420000  5.170000 ;
        RECT 1.050000 -0.225000 1.280000  5.170000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.180000 0.390000 5.170000 ;
      RECT 0.400000 5.340000 1.070000 5.670000 ;
      RECT 0.650000 0.180000 0.820000 5.170000 ;
      RECT 1.080000 0.180000 1.250000 5.170000 ;
    LAYER mcon ;
      RECT 0.220000 0.435000 0.390000 0.605000 ;
      RECT 0.220000 0.795000 0.390000 0.965000 ;
      RECT 0.220000 1.155000 0.390000 1.325000 ;
      RECT 0.220000 1.515000 0.390000 1.685000 ;
      RECT 0.220000 1.875000 0.390000 2.045000 ;
      RECT 0.220000 2.235000 0.390000 2.405000 ;
      RECT 0.220000 2.595000 0.390000 2.765000 ;
      RECT 0.220000 2.955000 0.390000 3.125000 ;
      RECT 0.220000 3.315000 0.390000 3.485000 ;
      RECT 0.220000 3.675000 0.390000 3.845000 ;
      RECT 0.220000 4.035000 0.390000 4.205000 ;
      RECT 0.220000 4.395000 0.390000 4.565000 ;
      RECT 0.220000 4.755000 0.390000 4.925000 ;
      RECT 0.470000 5.420000 0.640000 5.590000 ;
      RECT 0.650000 0.435000 0.820000 0.605000 ;
      RECT 0.650000 0.795000 0.820000 0.965000 ;
      RECT 0.650000 1.155000 0.820000 1.325000 ;
      RECT 0.650000 1.515000 0.820000 1.685000 ;
      RECT 0.650000 1.875000 0.820000 2.045000 ;
      RECT 0.650000 2.235000 0.820000 2.405000 ;
      RECT 0.650000 2.595000 0.820000 2.765000 ;
      RECT 0.650000 2.955000 0.820000 3.125000 ;
      RECT 0.650000 3.315000 0.820000 3.485000 ;
      RECT 0.650000 3.675000 0.820000 3.845000 ;
      RECT 0.650000 4.035000 0.820000 4.205000 ;
      RECT 0.650000 4.395000 0.820000 4.565000 ;
      RECT 0.650000 4.755000 0.820000 4.925000 ;
      RECT 0.830000 5.420000 1.000000 5.590000 ;
      RECT 1.080000 0.435000 1.250000 0.605000 ;
      RECT 1.080000 0.795000 1.250000 0.965000 ;
      RECT 1.080000 1.155000 1.250000 1.325000 ;
      RECT 1.080000 1.515000 1.250000 1.685000 ;
      RECT 1.080000 1.875000 1.250000 2.045000 ;
      RECT 1.080000 2.235000 1.250000 2.405000 ;
      RECT 1.080000 2.595000 1.250000 2.765000 ;
      RECT 1.080000 2.955000 1.250000 3.125000 ;
      RECT 1.080000 3.315000 1.250000 3.485000 ;
      RECT 1.080000 3.675000 1.250000 3.845000 ;
      RECT 1.080000 4.035000 1.250000 4.205000 ;
      RECT 1.080000 4.395000 1.250000 4.565000 ;
      RECT 1.080000 4.755000 1.250000 4.925000 ;
    LAYER met1 ;
      RECT 0.605000 0.180000 0.865000 5.170000 ;
    LAYER via ;
      RECT 0.605000 4.550000 0.865000 4.810000 ;
      RECT 0.605000 4.870000 0.865000 5.130000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
END LIBRARY
