MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 45.71 BY 60.23 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 15.34 2.78 15.62 13.18 ;
      LAYER M3 ;
        RECT 29.1 2.78 29.38 8.98 ;
      LAYER M3 ;
        RECT 15.34 6.115 15.62 6.485 ;
      LAYER M2 ;
        RECT 15.48 6.16 29.24 6.44 ;
      LAYER M3 ;
        RECT 29.1 6.115 29.38 6.485 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 35.12 27.98 35.4 34.18 ;
      LAYER M3 ;
        RECT 33.83 34.7 34.11 52.66 ;
      LAYER M3 ;
        RECT 35.12 34.02 35.4 34.44 ;
      LAYER M2 ;
        RECT 33.97 34.3 35.26 34.58 ;
      LAYER M3 ;
        RECT 33.83 34.44 34.11 34.86 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 16.24 21.24 16.52 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 23.48 16.24 35 16.52 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 9.32 27.98 9.6 34.18 ;
  LAYER M3 ;
        RECT 11.04 34.7 11.32 56.86 ;
  LAYER M3 ;
        RECT 33.4 38.9 33.68 56.86 ;
  LAYER M3 ;
        RECT 9.32 34.02 9.6 34.44 ;
  LAYER M2 ;
        RECT 9.46 34.3 11.18 34.58 ;
  LAYER M3 ;
        RECT 11.04 34.44 11.32 34.86 ;
  LAYER M3 ;
        RECT 11.04 41.395 11.32 41.765 ;
  LAYER M2 ;
        RECT 11.18 41.44 33.54 41.72 ;
  LAYER M3 ;
        RECT 33.4 41.395 33.68 41.765 ;
  LAYER M2 ;
        RECT 9.3 34.3 9.62 34.58 ;
  LAYER M3 ;
        RECT 9.32 34.28 9.6 34.6 ;
  LAYER M2 ;
        RECT 11.02 34.3 11.34 34.58 ;
  LAYER M3 ;
        RECT 11.04 34.28 11.32 34.6 ;
  LAYER M2 ;
        RECT 9.3 34.3 9.62 34.58 ;
  LAYER M3 ;
        RECT 9.32 34.28 9.6 34.6 ;
  LAYER M2 ;
        RECT 11.02 34.3 11.34 34.58 ;
  LAYER M3 ;
        RECT 11.04 34.28 11.32 34.6 ;
  LAYER M2 ;
        RECT 9.3 34.3 9.62 34.58 ;
  LAYER M3 ;
        RECT 9.32 34.28 9.6 34.6 ;
  LAYER M2 ;
        RECT 11.02 34.3 11.34 34.58 ;
  LAYER M3 ;
        RECT 11.04 34.28 11.32 34.6 ;
  LAYER M2 ;
        RECT 11.02 41.44 11.34 41.72 ;
  LAYER M3 ;
        RECT 11.04 41.42 11.32 41.74 ;
  LAYER M2 ;
        RECT 33.38 41.44 33.7 41.72 ;
  LAYER M3 ;
        RECT 33.4 41.42 33.68 41.74 ;
  LAYER M2 ;
        RECT 9.3 34.3 9.62 34.58 ;
  LAYER M3 ;
        RECT 9.32 34.28 9.6 34.6 ;
  LAYER M2 ;
        RECT 11.02 34.3 11.34 34.58 ;
  LAYER M3 ;
        RECT 11.04 34.28 11.32 34.6 ;
  LAYER M2 ;
        RECT 11.02 41.44 11.34 41.72 ;
  LAYER M3 ;
        RECT 11.04 41.42 11.32 41.74 ;
  LAYER M2 ;
        RECT 33.38 41.44 33.7 41.72 ;
  LAYER M3 ;
        RECT 33.4 41.42 33.68 41.74 ;
  LAYER M3 ;
        RECT 8.89 23.78 9.17 29.98 ;
  LAYER M2 ;
        RECT 9.72 20.44 21.24 20.72 ;
  LAYER M3 ;
        RECT 19.21 21.26 19.49 25.78 ;
  LAYER M3 ;
        RECT 8.89 20.58 9.17 23.94 ;
  LAYER M2 ;
        RECT 9.03 20.44 9.89 20.72 ;
  LAYER M2 ;
        RECT 19.19 20.44 19.51 20.72 ;
  LAYER M3 ;
        RECT 19.21 20.58 19.49 21.42 ;
  LAYER M2 ;
        RECT 8.87 20.44 9.19 20.72 ;
  LAYER M3 ;
        RECT 8.89 20.42 9.17 20.74 ;
  LAYER M2 ;
        RECT 8.87 20.44 9.19 20.72 ;
  LAYER M3 ;
        RECT 8.89 20.42 9.17 20.74 ;
  LAYER M2 ;
        RECT 8.87 20.44 9.19 20.72 ;
  LAYER M3 ;
        RECT 8.89 20.42 9.17 20.74 ;
  LAYER M2 ;
        RECT 19.19 20.44 19.51 20.72 ;
  LAYER M3 ;
        RECT 19.21 20.42 19.49 20.74 ;
  LAYER M2 ;
        RECT 8.87 20.44 9.19 20.72 ;
  LAYER M3 ;
        RECT 8.89 20.42 9.17 20.74 ;
  LAYER M2 ;
        RECT 19.19 20.44 19.51 20.72 ;
  LAYER M3 ;
        RECT 19.21 20.42 19.49 20.74 ;
  LAYER M3 ;
        RECT 25.23 21.26 25.51 25.78 ;
  LAYER M2 ;
        RECT 23.48 20.44 35 20.72 ;
  LAYER M3 ;
        RECT 35.55 23.78 35.83 29.98 ;
  LAYER M3 ;
        RECT 25.23 20.58 25.51 21.42 ;
  LAYER M2 ;
        RECT 25.21 20.44 25.53 20.72 ;
  LAYER M2 ;
        RECT 34.83 20.44 35.69 20.72 ;
  LAYER M3 ;
        RECT 35.55 20.58 35.83 23.94 ;
  LAYER M2 ;
        RECT 25.21 20.44 25.53 20.72 ;
  LAYER M3 ;
        RECT 25.23 20.42 25.51 20.74 ;
  LAYER M2 ;
        RECT 25.21 20.44 25.53 20.72 ;
  LAYER M3 ;
        RECT 25.23 20.42 25.51 20.74 ;
  LAYER M2 ;
        RECT 25.21 20.44 25.53 20.72 ;
  LAYER M3 ;
        RECT 25.23 20.42 25.51 20.74 ;
  LAYER M2 ;
        RECT 35.53 20.44 35.85 20.72 ;
  LAYER M3 ;
        RECT 35.55 20.42 35.83 20.74 ;
  LAYER M2 ;
        RECT 25.21 20.44 25.53 20.72 ;
  LAYER M3 ;
        RECT 25.23 20.42 25.51 20.74 ;
  LAYER M2 ;
        RECT 35.53 20.44 35.85 20.72 ;
  LAYER M3 ;
        RECT 35.55 20.42 35.83 20.74 ;
  LAYER M2 ;
        RECT 9.29 20.02 21.67 20.3 ;
  LAYER M2 ;
        RECT 23.05 20.02 35.43 20.3 ;
  LAYER M3 ;
        RECT 28.67 6.98 28.95 13.18 ;
  LAYER M2 ;
        RECT 21.5 20.02 23.22 20.3 ;
  LAYER M2 ;
        RECT 28.65 20.02 28.97 20.3 ;
  LAYER M3 ;
        RECT 28.67 13.02 28.95 20.16 ;
  LAYER M2 ;
        RECT 28.65 20.02 28.97 20.3 ;
  LAYER M3 ;
        RECT 28.67 20 28.95 20.32 ;
  LAYER M2 ;
        RECT 28.65 20.02 28.97 20.3 ;
  LAYER M3 ;
        RECT 28.67 20 28.95 20.32 ;
  LAYER M1 ;
        RECT 20.945 9.575 21.195 13.105 ;
  LAYER M1 ;
        RECT 20.945 8.315 21.195 9.325 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 21.375 9.575 21.625 13.105 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 20.515 9.575 20.765 13.105 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 20.085 9.575 20.335 13.105 ;
  LAYER M1 ;
        RECT 20.085 8.315 20.335 9.325 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 19.655 9.575 19.905 13.105 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 19.225 9.575 19.475 13.105 ;
  LAYER M1 ;
        RECT 19.225 8.315 19.475 9.325 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 9.575 19.045 13.105 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 18.365 9.575 18.615 13.105 ;
  LAYER M1 ;
        RECT 18.365 8.315 18.615 9.325 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 17.935 9.575 18.185 13.105 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.505 9.575 17.755 13.105 ;
  LAYER M1 ;
        RECT 17.505 8.315 17.755 9.325 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 9.575 16.895 13.105 ;
  LAYER M1 ;
        RECT 16.645 8.315 16.895 9.325 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 9.575 15.175 13.105 ;
  LAYER M1 ;
        RECT 14.925 8.315 15.175 9.325 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 9.575 12.595 13.105 ;
  LAYER M1 ;
        RECT 12.345 8.315 12.595 9.325 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 9.575 12.165 13.105 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.485 9.575 11.735 13.105 ;
  LAYER M1 ;
        RECT 11.485 8.315 11.735 9.325 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.72 12.88 21.24 13.16 ;
  LAYER M2 ;
        RECT 9.72 8.68 21.24 8.96 ;
  LAYER M2 ;
        RECT 9.29 12.46 21.67 12.74 ;
  LAYER M2 ;
        RECT 9.72 7 21.24 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 21.24 3.08 ;
  LAYER M2 ;
        RECT 9.72 0.7 21.24 0.98 ;
  LAYER M2 ;
        RECT 9.29 6.58 21.67 6.86 ;
  LAYER M3 ;
        RECT 15.34 2.78 15.62 13.18 ;
  LAYER M3 ;
        RECT 14.91 0.68 15.19 12.76 ;
  LAYER M1 ;
        RECT 1.165 34.775 1.415 38.305 ;
  LAYER M1 ;
        RECT 1.165 38.555 1.415 39.565 ;
  LAYER M1 ;
        RECT 1.165 40.655 1.415 44.185 ;
  LAYER M1 ;
        RECT 1.165 44.435 1.415 45.445 ;
  LAYER M1 ;
        RECT 1.165 46.535 1.415 50.065 ;
  LAYER M1 ;
        RECT 1.165 50.315 1.415 51.325 ;
  LAYER M1 ;
        RECT 1.165 52.415 1.415 55.945 ;
  LAYER M1 ;
        RECT 1.165 56.195 1.415 57.205 ;
  LAYER M1 ;
        RECT 1.165 58.295 1.415 59.305 ;
  LAYER M1 ;
        RECT 0.735 34.775 0.985 38.305 ;
  LAYER M1 ;
        RECT 0.735 40.655 0.985 44.185 ;
  LAYER M1 ;
        RECT 0.735 46.535 0.985 50.065 ;
  LAYER M1 ;
        RECT 0.735 52.415 0.985 55.945 ;
  LAYER M1 ;
        RECT 1.595 34.775 1.845 38.305 ;
  LAYER M1 ;
        RECT 1.595 40.655 1.845 44.185 ;
  LAYER M1 ;
        RECT 1.595 46.535 1.845 50.065 ;
  LAYER M1 ;
        RECT 1.595 52.415 1.845 55.945 ;
  LAYER M1 ;
        RECT 2.025 34.775 2.275 38.305 ;
  LAYER M1 ;
        RECT 2.025 38.555 2.275 39.565 ;
  LAYER M1 ;
        RECT 2.025 40.655 2.275 44.185 ;
  LAYER M1 ;
        RECT 2.025 44.435 2.275 45.445 ;
  LAYER M1 ;
        RECT 2.025 46.535 2.275 50.065 ;
  LAYER M1 ;
        RECT 2.025 50.315 2.275 51.325 ;
  LAYER M1 ;
        RECT 2.025 52.415 2.275 55.945 ;
  LAYER M1 ;
        RECT 2.025 56.195 2.275 57.205 ;
  LAYER M1 ;
        RECT 2.025 58.295 2.275 59.305 ;
  LAYER M1 ;
        RECT 2.455 34.775 2.705 38.305 ;
  LAYER M1 ;
        RECT 2.455 40.655 2.705 44.185 ;
  LAYER M1 ;
        RECT 2.455 46.535 2.705 50.065 ;
  LAYER M1 ;
        RECT 2.455 52.415 2.705 55.945 ;
  LAYER M1 ;
        RECT 2.885 34.775 3.135 38.305 ;
  LAYER M1 ;
        RECT 2.885 38.555 3.135 39.565 ;
  LAYER M1 ;
        RECT 2.885 40.655 3.135 44.185 ;
  LAYER M1 ;
        RECT 2.885 44.435 3.135 45.445 ;
  LAYER M1 ;
        RECT 2.885 46.535 3.135 50.065 ;
  LAYER M1 ;
        RECT 2.885 50.315 3.135 51.325 ;
  LAYER M1 ;
        RECT 2.885 52.415 3.135 55.945 ;
  LAYER M1 ;
        RECT 2.885 56.195 3.135 57.205 ;
  LAYER M1 ;
        RECT 2.885 58.295 3.135 59.305 ;
  LAYER M1 ;
        RECT 3.315 34.775 3.565 38.305 ;
  LAYER M1 ;
        RECT 3.315 40.655 3.565 44.185 ;
  LAYER M1 ;
        RECT 3.315 46.535 3.565 50.065 ;
  LAYER M1 ;
        RECT 3.315 52.415 3.565 55.945 ;
  LAYER M1 ;
        RECT 3.745 34.775 3.995 38.305 ;
  LAYER M1 ;
        RECT 3.745 38.555 3.995 39.565 ;
  LAYER M1 ;
        RECT 3.745 40.655 3.995 44.185 ;
  LAYER M1 ;
        RECT 3.745 44.435 3.995 45.445 ;
  LAYER M1 ;
        RECT 3.745 46.535 3.995 50.065 ;
  LAYER M1 ;
        RECT 3.745 50.315 3.995 51.325 ;
  LAYER M1 ;
        RECT 3.745 52.415 3.995 55.945 ;
  LAYER M1 ;
        RECT 3.745 56.195 3.995 57.205 ;
  LAYER M1 ;
        RECT 3.745 58.295 3.995 59.305 ;
  LAYER M1 ;
        RECT 4.175 34.775 4.425 38.305 ;
  LAYER M1 ;
        RECT 4.175 40.655 4.425 44.185 ;
  LAYER M1 ;
        RECT 4.175 46.535 4.425 50.065 ;
  LAYER M1 ;
        RECT 4.175 52.415 4.425 55.945 ;
  LAYER M1 ;
        RECT 4.605 34.775 4.855 38.305 ;
  LAYER M1 ;
        RECT 4.605 38.555 4.855 39.565 ;
  LAYER M1 ;
        RECT 4.605 40.655 4.855 44.185 ;
  LAYER M1 ;
        RECT 4.605 44.435 4.855 45.445 ;
  LAYER M1 ;
        RECT 4.605 46.535 4.855 50.065 ;
  LAYER M1 ;
        RECT 4.605 50.315 4.855 51.325 ;
  LAYER M1 ;
        RECT 4.605 52.415 4.855 55.945 ;
  LAYER M1 ;
        RECT 4.605 56.195 4.855 57.205 ;
  LAYER M1 ;
        RECT 4.605 58.295 4.855 59.305 ;
  LAYER M1 ;
        RECT 5.035 34.775 5.285 38.305 ;
  LAYER M1 ;
        RECT 5.035 40.655 5.285 44.185 ;
  LAYER M1 ;
        RECT 5.035 46.535 5.285 50.065 ;
  LAYER M1 ;
        RECT 5.035 52.415 5.285 55.945 ;
  LAYER M1 ;
        RECT 5.465 34.775 5.715 38.305 ;
  LAYER M1 ;
        RECT 5.465 38.555 5.715 39.565 ;
  LAYER M1 ;
        RECT 5.465 40.655 5.715 44.185 ;
  LAYER M1 ;
        RECT 5.465 44.435 5.715 45.445 ;
  LAYER M1 ;
        RECT 5.465 46.535 5.715 50.065 ;
  LAYER M1 ;
        RECT 5.465 50.315 5.715 51.325 ;
  LAYER M1 ;
        RECT 5.465 52.415 5.715 55.945 ;
  LAYER M1 ;
        RECT 5.465 56.195 5.715 57.205 ;
  LAYER M1 ;
        RECT 5.465 58.295 5.715 59.305 ;
  LAYER M1 ;
        RECT 5.895 34.775 6.145 38.305 ;
  LAYER M1 ;
        RECT 5.895 40.655 6.145 44.185 ;
  LAYER M1 ;
        RECT 5.895 46.535 6.145 50.065 ;
  LAYER M1 ;
        RECT 5.895 52.415 6.145 55.945 ;
  LAYER M1 ;
        RECT 6.325 34.775 6.575 38.305 ;
  LAYER M1 ;
        RECT 6.325 38.555 6.575 39.565 ;
  LAYER M1 ;
        RECT 6.325 40.655 6.575 44.185 ;
  LAYER M1 ;
        RECT 6.325 44.435 6.575 45.445 ;
  LAYER M1 ;
        RECT 6.325 46.535 6.575 50.065 ;
  LAYER M1 ;
        RECT 6.325 50.315 6.575 51.325 ;
  LAYER M1 ;
        RECT 6.325 52.415 6.575 55.945 ;
  LAYER M1 ;
        RECT 6.325 56.195 6.575 57.205 ;
  LAYER M1 ;
        RECT 6.325 58.295 6.575 59.305 ;
  LAYER M1 ;
        RECT 6.755 34.775 7.005 38.305 ;
  LAYER M1 ;
        RECT 6.755 40.655 7.005 44.185 ;
  LAYER M1 ;
        RECT 6.755 46.535 7.005 50.065 ;
  LAYER M1 ;
        RECT 6.755 52.415 7.005 55.945 ;
  LAYER M1 ;
        RECT 7.185 34.775 7.435 38.305 ;
  LAYER M1 ;
        RECT 7.185 38.555 7.435 39.565 ;
  LAYER M1 ;
        RECT 7.185 40.655 7.435 44.185 ;
  LAYER M1 ;
        RECT 7.185 44.435 7.435 45.445 ;
  LAYER M1 ;
        RECT 7.185 46.535 7.435 50.065 ;
  LAYER M1 ;
        RECT 7.185 50.315 7.435 51.325 ;
  LAYER M1 ;
        RECT 7.185 52.415 7.435 55.945 ;
  LAYER M1 ;
        RECT 7.185 56.195 7.435 57.205 ;
  LAYER M1 ;
        RECT 7.185 58.295 7.435 59.305 ;
  LAYER M1 ;
        RECT 7.615 34.775 7.865 38.305 ;
  LAYER M1 ;
        RECT 7.615 40.655 7.865 44.185 ;
  LAYER M1 ;
        RECT 7.615 46.535 7.865 50.065 ;
  LAYER M1 ;
        RECT 7.615 52.415 7.865 55.945 ;
  LAYER M1 ;
        RECT 8.045 34.775 8.295 38.305 ;
  LAYER M1 ;
        RECT 8.045 38.555 8.295 39.565 ;
  LAYER M1 ;
        RECT 8.045 40.655 8.295 44.185 ;
  LAYER M1 ;
        RECT 8.045 44.435 8.295 45.445 ;
  LAYER M1 ;
        RECT 8.045 46.535 8.295 50.065 ;
  LAYER M1 ;
        RECT 8.045 50.315 8.295 51.325 ;
  LAYER M1 ;
        RECT 8.045 52.415 8.295 55.945 ;
  LAYER M1 ;
        RECT 8.045 56.195 8.295 57.205 ;
  LAYER M1 ;
        RECT 8.045 58.295 8.295 59.305 ;
  LAYER M1 ;
        RECT 8.475 34.775 8.725 38.305 ;
  LAYER M1 ;
        RECT 8.475 40.655 8.725 44.185 ;
  LAYER M1 ;
        RECT 8.475 46.535 8.725 50.065 ;
  LAYER M1 ;
        RECT 8.475 52.415 8.725 55.945 ;
  LAYER M1 ;
        RECT 8.905 34.775 9.155 38.305 ;
  LAYER M1 ;
        RECT 8.905 38.555 9.155 39.565 ;
  LAYER M1 ;
        RECT 8.905 40.655 9.155 44.185 ;
  LAYER M1 ;
        RECT 8.905 44.435 9.155 45.445 ;
  LAYER M1 ;
        RECT 8.905 46.535 9.155 50.065 ;
  LAYER M1 ;
        RECT 8.905 50.315 9.155 51.325 ;
  LAYER M1 ;
        RECT 8.905 52.415 9.155 55.945 ;
  LAYER M1 ;
        RECT 8.905 56.195 9.155 57.205 ;
  LAYER M1 ;
        RECT 8.905 58.295 9.155 59.305 ;
  LAYER M1 ;
        RECT 9.335 34.775 9.585 38.305 ;
  LAYER M1 ;
        RECT 9.335 40.655 9.585 44.185 ;
  LAYER M1 ;
        RECT 9.335 46.535 9.585 50.065 ;
  LAYER M1 ;
        RECT 9.335 52.415 9.585 55.945 ;
  LAYER M1 ;
        RECT 9.765 34.775 10.015 38.305 ;
  LAYER M1 ;
        RECT 9.765 38.555 10.015 39.565 ;
  LAYER M1 ;
        RECT 9.765 40.655 10.015 44.185 ;
  LAYER M1 ;
        RECT 9.765 44.435 10.015 45.445 ;
  LAYER M1 ;
        RECT 9.765 46.535 10.015 50.065 ;
  LAYER M1 ;
        RECT 9.765 50.315 10.015 51.325 ;
  LAYER M1 ;
        RECT 9.765 52.415 10.015 55.945 ;
  LAYER M1 ;
        RECT 9.765 56.195 10.015 57.205 ;
  LAYER M1 ;
        RECT 9.765 58.295 10.015 59.305 ;
  LAYER M1 ;
        RECT 10.195 34.775 10.445 38.305 ;
  LAYER M1 ;
        RECT 10.195 40.655 10.445 44.185 ;
  LAYER M1 ;
        RECT 10.195 46.535 10.445 50.065 ;
  LAYER M1 ;
        RECT 10.195 52.415 10.445 55.945 ;
  LAYER M1 ;
        RECT 10.625 34.775 10.875 38.305 ;
  LAYER M1 ;
        RECT 10.625 38.555 10.875 39.565 ;
  LAYER M1 ;
        RECT 10.625 40.655 10.875 44.185 ;
  LAYER M1 ;
        RECT 10.625 44.435 10.875 45.445 ;
  LAYER M1 ;
        RECT 10.625 46.535 10.875 50.065 ;
  LAYER M1 ;
        RECT 10.625 50.315 10.875 51.325 ;
  LAYER M1 ;
        RECT 10.625 52.415 10.875 55.945 ;
  LAYER M1 ;
        RECT 10.625 56.195 10.875 57.205 ;
  LAYER M1 ;
        RECT 10.625 58.295 10.875 59.305 ;
  LAYER M1 ;
        RECT 11.055 34.775 11.305 38.305 ;
  LAYER M1 ;
        RECT 11.055 40.655 11.305 44.185 ;
  LAYER M1 ;
        RECT 11.055 46.535 11.305 50.065 ;
  LAYER M1 ;
        RECT 11.055 52.415 11.305 55.945 ;
  LAYER M1 ;
        RECT 11.485 34.775 11.735 38.305 ;
  LAYER M1 ;
        RECT 11.485 38.555 11.735 39.565 ;
  LAYER M1 ;
        RECT 11.485 40.655 11.735 44.185 ;
  LAYER M1 ;
        RECT 11.485 44.435 11.735 45.445 ;
  LAYER M1 ;
        RECT 11.485 46.535 11.735 50.065 ;
  LAYER M1 ;
        RECT 11.485 50.315 11.735 51.325 ;
  LAYER M1 ;
        RECT 11.485 52.415 11.735 55.945 ;
  LAYER M1 ;
        RECT 11.485 56.195 11.735 57.205 ;
  LAYER M1 ;
        RECT 11.485 58.295 11.735 59.305 ;
  LAYER M1 ;
        RECT 11.915 34.775 12.165 38.305 ;
  LAYER M1 ;
        RECT 11.915 40.655 12.165 44.185 ;
  LAYER M1 ;
        RECT 11.915 46.535 12.165 50.065 ;
  LAYER M1 ;
        RECT 11.915 52.415 12.165 55.945 ;
  LAYER M1 ;
        RECT 12.345 34.775 12.595 38.305 ;
  LAYER M1 ;
        RECT 12.345 38.555 12.595 39.565 ;
  LAYER M1 ;
        RECT 12.345 40.655 12.595 44.185 ;
  LAYER M1 ;
        RECT 12.345 44.435 12.595 45.445 ;
  LAYER M1 ;
        RECT 12.345 46.535 12.595 50.065 ;
  LAYER M1 ;
        RECT 12.345 50.315 12.595 51.325 ;
  LAYER M1 ;
        RECT 12.345 52.415 12.595 55.945 ;
  LAYER M1 ;
        RECT 12.345 56.195 12.595 57.205 ;
  LAYER M1 ;
        RECT 12.345 58.295 12.595 59.305 ;
  LAYER M1 ;
        RECT 12.775 34.775 13.025 38.305 ;
  LAYER M1 ;
        RECT 12.775 40.655 13.025 44.185 ;
  LAYER M1 ;
        RECT 12.775 46.535 13.025 50.065 ;
  LAYER M1 ;
        RECT 12.775 52.415 13.025 55.945 ;
  LAYER M1 ;
        RECT 13.205 34.775 13.455 38.305 ;
  LAYER M1 ;
        RECT 13.205 38.555 13.455 39.565 ;
  LAYER M1 ;
        RECT 13.205 40.655 13.455 44.185 ;
  LAYER M1 ;
        RECT 13.205 44.435 13.455 45.445 ;
  LAYER M1 ;
        RECT 13.205 46.535 13.455 50.065 ;
  LAYER M1 ;
        RECT 13.205 50.315 13.455 51.325 ;
  LAYER M1 ;
        RECT 13.205 52.415 13.455 55.945 ;
  LAYER M1 ;
        RECT 13.205 56.195 13.455 57.205 ;
  LAYER M1 ;
        RECT 13.205 58.295 13.455 59.305 ;
  LAYER M1 ;
        RECT 13.635 34.775 13.885 38.305 ;
  LAYER M1 ;
        RECT 13.635 40.655 13.885 44.185 ;
  LAYER M1 ;
        RECT 13.635 46.535 13.885 50.065 ;
  LAYER M1 ;
        RECT 13.635 52.415 13.885 55.945 ;
  LAYER M1 ;
        RECT 14.065 34.775 14.315 38.305 ;
  LAYER M1 ;
        RECT 14.065 38.555 14.315 39.565 ;
  LAYER M1 ;
        RECT 14.065 40.655 14.315 44.185 ;
  LAYER M1 ;
        RECT 14.065 44.435 14.315 45.445 ;
  LAYER M1 ;
        RECT 14.065 46.535 14.315 50.065 ;
  LAYER M1 ;
        RECT 14.065 50.315 14.315 51.325 ;
  LAYER M1 ;
        RECT 14.065 52.415 14.315 55.945 ;
  LAYER M1 ;
        RECT 14.065 56.195 14.315 57.205 ;
  LAYER M1 ;
        RECT 14.065 58.295 14.315 59.305 ;
  LAYER M1 ;
        RECT 14.495 34.775 14.745 38.305 ;
  LAYER M1 ;
        RECT 14.495 40.655 14.745 44.185 ;
  LAYER M1 ;
        RECT 14.495 46.535 14.745 50.065 ;
  LAYER M1 ;
        RECT 14.495 52.415 14.745 55.945 ;
  LAYER M1 ;
        RECT 14.925 34.775 15.175 38.305 ;
  LAYER M1 ;
        RECT 14.925 38.555 15.175 39.565 ;
  LAYER M1 ;
        RECT 14.925 40.655 15.175 44.185 ;
  LAYER M1 ;
        RECT 14.925 44.435 15.175 45.445 ;
  LAYER M1 ;
        RECT 14.925 46.535 15.175 50.065 ;
  LAYER M1 ;
        RECT 14.925 50.315 15.175 51.325 ;
  LAYER M1 ;
        RECT 14.925 52.415 15.175 55.945 ;
  LAYER M1 ;
        RECT 14.925 56.195 15.175 57.205 ;
  LAYER M1 ;
        RECT 14.925 58.295 15.175 59.305 ;
  LAYER M1 ;
        RECT 15.355 34.775 15.605 38.305 ;
  LAYER M1 ;
        RECT 15.355 40.655 15.605 44.185 ;
  LAYER M1 ;
        RECT 15.355 46.535 15.605 50.065 ;
  LAYER M1 ;
        RECT 15.355 52.415 15.605 55.945 ;
  LAYER M1 ;
        RECT 15.785 34.775 16.035 38.305 ;
  LAYER M1 ;
        RECT 15.785 38.555 16.035 39.565 ;
  LAYER M1 ;
        RECT 15.785 40.655 16.035 44.185 ;
  LAYER M1 ;
        RECT 15.785 44.435 16.035 45.445 ;
  LAYER M1 ;
        RECT 15.785 46.535 16.035 50.065 ;
  LAYER M1 ;
        RECT 15.785 50.315 16.035 51.325 ;
  LAYER M1 ;
        RECT 15.785 52.415 16.035 55.945 ;
  LAYER M1 ;
        RECT 15.785 56.195 16.035 57.205 ;
  LAYER M1 ;
        RECT 15.785 58.295 16.035 59.305 ;
  LAYER M1 ;
        RECT 16.215 34.775 16.465 38.305 ;
  LAYER M1 ;
        RECT 16.215 40.655 16.465 44.185 ;
  LAYER M1 ;
        RECT 16.215 46.535 16.465 50.065 ;
  LAYER M1 ;
        RECT 16.215 52.415 16.465 55.945 ;
  LAYER M1 ;
        RECT 16.645 34.775 16.895 38.305 ;
  LAYER M1 ;
        RECT 16.645 38.555 16.895 39.565 ;
  LAYER M1 ;
        RECT 16.645 40.655 16.895 44.185 ;
  LAYER M1 ;
        RECT 16.645 44.435 16.895 45.445 ;
  LAYER M1 ;
        RECT 16.645 46.535 16.895 50.065 ;
  LAYER M1 ;
        RECT 16.645 50.315 16.895 51.325 ;
  LAYER M1 ;
        RECT 16.645 52.415 16.895 55.945 ;
  LAYER M1 ;
        RECT 16.645 56.195 16.895 57.205 ;
  LAYER M1 ;
        RECT 16.645 58.295 16.895 59.305 ;
  LAYER M1 ;
        RECT 17.075 34.775 17.325 38.305 ;
  LAYER M1 ;
        RECT 17.075 40.655 17.325 44.185 ;
  LAYER M1 ;
        RECT 17.075 46.535 17.325 50.065 ;
  LAYER M1 ;
        RECT 17.075 52.415 17.325 55.945 ;
  LAYER M1 ;
        RECT 17.505 34.775 17.755 38.305 ;
  LAYER M1 ;
        RECT 17.505 38.555 17.755 39.565 ;
  LAYER M1 ;
        RECT 17.505 40.655 17.755 44.185 ;
  LAYER M1 ;
        RECT 17.505 44.435 17.755 45.445 ;
  LAYER M1 ;
        RECT 17.505 46.535 17.755 50.065 ;
  LAYER M1 ;
        RECT 17.505 50.315 17.755 51.325 ;
  LAYER M1 ;
        RECT 17.505 52.415 17.755 55.945 ;
  LAYER M1 ;
        RECT 17.505 56.195 17.755 57.205 ;
  LAYER M1 ;
        RECT 17.505 58.295 17.755 59.305 ;
  LAYER M1 ;
        RECT 17.935 34.775 18.185 38.305 ;
  LAYER M1 ;
        RECT 17.935 40.655 18.185 44.185 ;
  LAYER M1 ;
        RECT 17.935 46.535 18.185 50.065 ;
  LAYER M1 ;
        RECT 17.935 52.415 18.185 55.945 ;
  LAYER M1 ;
        RECT 18.365 34.775 18.615 38.305 ;
  LAYER M1 ;
        RECT 18.365 38.555 18.615 39.565 ;
  LAYER M1 ;
        RECT 18.365 40.655 18.615 44.185 ;
  LAYER M1 ;
        RECT 18.365 44.435 18.615 45.445 ;
  LAYER M1 ;
        RECT 18.365 46.535 18.615 50.065 ;
  LAYER M1 ;
        RECT 18.365 50.315 18.615 51.325 ;
  LAYER M1 ;
        RECT 18.365 52.415 18.615 55.945 ;
  LAYER M1 ;
        RECT 18.365 56.195 18.615 57.205 ;
  LAYER M1 ;
        RECT 18.365 58.295 18.615 59.305 ;
  LAYER M1 ;
        RECT 18.795 34.775 19.045 38.305 ;
  LAYER M1 ;
        RECT 18.795 40.655 19.045 44.185 ;
  LAYER M1 ;
        RECT 18.795 46.535 19.045 50.065 ;
  LAYER M1 ;
        RECT 18.795 52.415 19.045 55.945 ;
  LAYER M1 ;
        RECT 19.225 34.775 19.475 38.305 ;
  LAYER M1 ;
        RECT 19.225 38.555 19.475 39.565 ;
  LAYER M1 ;
        RECT 19.225 40.655 19.475 44.185 ;
  LAYER M1 ;
        RECT 19.225 44.435 19.475 45.445 ;
  LAYER M1 ;
        RECT 19.225 46.535 19.475 50.065 ;
  LAYER M1 ;
        RECT 19.225 50.315 19.475 51.325 ;
  LAYER M1 ;
        RECT 19.225 52.415 19.475 55.945 ;
  LAYER M1 ;
        RECT 19.225 56.195 19.475 57.205 ;
  LAYER M1 ;
        RECT 19.225 58.295 19.475 59.305 ;
  LAYER M1 ;
        RECT 19.655 34.775 19.905 38.305 ;
  LAYER M1 ;
        RECT 19.655 40.655 19.905 44.185 ;
  LAYER M1 ;
        RECT 19.655 46.535 19.905 50.065 ;
  LAYER M1 ;
        RECT 19.655 52.415 19.905 55.945 ;
  LAYER M1 ;
        RECT 20.085 34.775 20.335 38.305 ;
  LAYER M1 ;
        RECT 20.085 38.555 20.335 39.565 ;
  LAYER M1 ;
        RECT 20.085 40.655 20.335 44.185 ;
  LAYER M1 ;
        RECT 20.085 44.435 20.335 45.445 ;
  LAYER M1 ;
        RECT 20.085 46.535 20.335 50.065 ;
  LAYER M1 ;
        RECT 20.085 50.315 20.335 51.325 ;
  LAYER M1 ;
        RECT 20.085 52.415 20.335 55.945 ;
  LAYER M1 ;
        RECT 20.085 56.195 20.335 57.205 ;
  LAYER M1 ;
        RECT 20.085 58.295 20.335 59.305 ;
  LAYER M1 ;
        RECT 20.515 34.775 20.765 38.305 ;
  LAYER M1 ;
        RECT 20.515 40.655 20.765 44.185 ;
  LAYER M1 ;
        RECT 20.515 46.535 20.765 50.065 ;
  LAYER M1 ;
        RECT 20.515 52.415 20.765 55.945 ;
  LAYER M1 ;
        RECT 20.945 34.775 21.195 38.305 ;
  LAYER M1 ;
        RECT 20.945 38.555 21.195 39.565 ;
  LAYER M1 ;
        RECT 20.945 40.655 21.195 44.185 ;
  LAYER M1 ;
        RECT 20.945 44.435 21.195 45.445 ;
  LAYER M1 ;
        RECT 20.945 46.535 21.195 50.065 ;
  LAYER M1 ;
        RECT 20.945 50.315 21.195 51.325 ;
  LAYER M1 ;
        RECT 20.945 52.415 21.195 55.945 ;
  LAYER M1 ;
        RECT 20.945 56.195 21.195 57.205 ;
  LAYER M1 ;
        RECT 20.945 58.295 21.195 59.305 ;
  LAYER M1 ;
        RECT 21.375 34.775 21.625 38.305 ;
  LAYER M1 ;
        RECT 21.375 40.655 21.625 44.185 ;
  LAYER M1 ;
        RECT 21.375 46.535 21.625 50.065 ;
  LAYER M1 ;
        RECT 21.375 52.415 21.625 55.945 ;
  LAYER M2 ;
        RECT 1.12 34.72 21.24 35 ;
  LAYER M2 ;
        RECT 1.12 38.92 21.24 39.2 ;
  LAYER M2 ;
        RECT 0.69 35.14 21.67 35.42 ;
  LAYER M2 ;
        RECT 1.12 40.6 21.24 40.88 ;
  LAYER M2 ;
        RECT 1.12 44.8 21.24 45.08 ;
  LAYER M2 ;
        RECT 0.69 41.02 21.67 41.3 ;
  LAYER M2 ;
        RECT 1.12 46.48 21.24 46.76 ;
  LAYER M2 ;
        RECT 1.12 50.68 21.24 50.96 ;
  LAYER M2 ;
        RECT 0.69 46.9 21.67 47.18 ;
  LAYER M2 ;
        RECT 1.12 52.36 21.24 52.64 ;
  LAYER M2 ;
        RECT 1.12 56.56 21.24 56.84 ;
  LAYER M2 ;
        RECT 1.12 58.66 21.24 58.94 ;
  LAYER M2 ;
        RECT 0.69 52.78 21.67 53.06 ;
  LAYER M3 ;
        RECT 11.04 34.7 11.32 56.86 ;
  LAYER M3 ;
        RECT 11.47 35.12 11.75 58.96 ;
  LAYER M1 ;
        RECT 20.945 21.335 21.195 24.865 ;
  LAYER M1 ;
        RECT 20.945 25.115 21.195 26.125 ;
  LAYER M1 ;
        RECT 20.945 27.215 21.195 28.225 ;
  LAYER M1 ;
        RECT 21.375 21.335 21.625 24.865 ;
  LAYER M1 ;
        RECT 20.515 21.335 20.765 24.865 ;
  LAYER M1 ;
        RECT 20.085 21.335 20.335 24.865 ;
  LAYER M1 ;
        RECT 20.085 25.115 20.335 26.125 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 28.225 ;
  LAYER M1 ;
        RECT 19.655 21.335 19.905 24.865 ;
  LAYER M1 ;
        RECT 19.225 21.335 19.475 24.865 ;
  LAYER M1 ;
        RECT 19.225 25.115 19.475 26.125 ;
  LAYER M1 ;
        RECT 19.225 27.215 19.475 28.225 ;
  LAYER M1 ;
        RECT 18.795 21.335 19.045 24.865 ;
  LAYER M1 ;
        RECT 18.365 21.335 18.615 24.865 ;
  LAYER M1 ;
        RECT 18.365 25.115 18.615 26.125 ;
  LAYER M1 ;
        RECT 18.365 27.215 18.615 28.225 ;
  LAYER M1 ;
        RECT 17.935 21.335 18.185 24.865 ;
  LAYER M1 ;
        RECT 17.505 21.335 17.755 24.865 ;
  LAYER M1 ;
        RECT 17.505 25.115 17.755 26.125 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 28.225 ;
  LAYER M1 ;
        RECT 17.075 21.335 17.325 24.865 ;
  LAYER M2 ;
        RECT 17.46 21.28 21.24 21.56 ;
  LAYER M2 ;
        RECT 17.46 25.48 21.24 25.76 ;
  LAYER M2 ;
        RECT 17.46 27.58 21.24 27.86 ;
  LAYER M2 ;
        RECT 17.03 21.7 21.67 21.98 ;
  LAYER M3 ;
        RECT 19.21 21.26 19.49 25.78 ;
  LAYER M3 ;
        RECT 18.78 21.68 19.06 27.88 ;
  LAYER M1 ;
        RECT 23.525 21.335 23.775 24.865 ;
  LAYER M1 ;
        RECT 23.525 25.115 23.775 26.125 ;
  LAYER M1 ;
        RECT 23.525 27.215 23.775 28.225 ;
  LAYER M1 ;
        RECT 23.095 21.335 23.345 24.865 ;
  LAYER M1 ;
        RECT 23.955 21.335 24.205 24.865 ;
  LAYER M1 ;
        RECT 24.385 21.335 24.635 24.865 ;
  LAYER M1 ;
        RECT 24.385 25.115 24.635 26.125 ;
  LAYER M1 ;
        RECT 24.385 27.215 24.635 28.225 ;
  LAYER M1 ;
        RECT 24.815 21.335 25.065 24.865 ;
  LAYER M1 ;
        RECT 25.245 21.335 25.495 24.865 ;
  LAYER M1 ;
        RECT 25.245 25.115 25.495 26.125 ;
  LAYER M1 ;
        RECT 25.245 27.215 25.495 28.225 ;
  LAYER M1 ;
        RECT 25.675 21.335 25.925 24.865 ;
  LAYER M1 ;
        RECT 26.105 21.335 26.355 24.865 ;
  LAYER M1 ;
        RECT 26.105 25.115 26.355 26.125 ;
  LAYER M1 ;
        RECT 26.105 27.215 26.355 28.225 ;
  LAYER M1 ;
        RECT 26.535 21.335 26.785 24.865 ;
  LAYER M1 ;
        RECT 26.965 21.335 27.215 24.865 ;
  LAYER M1 ;
        RECT 26.965 25.115 27.215 26.125 ;
  LAYER M1 ;
        RECT 26.965 27.215 27.215 28.225 ;
  LAYER M1 ;
        RECT 27.395 21.335 27.645 24.865 ;
  LAYER M2 ;
        RECT 23.48 21.28 27.26 21.56 ;
  LAYER M2 ;
        RECT 23.48 25.48 27.26 25.76 ;
  LAYER M2 ;
        RECT 23.48 27.58 27.26 27.86 ;
  LAYER M2 ;
        RECT 23.05 21.7 27.69 21.98 ;
  LAYER M3 ;
        RECT 25.23 21.26 25.51 25.78 ;
  LAYER M3 ;
        RECT 25.66 21.68 25.94 27.88 ;
  LAYER M1 ;
        RECT 43.305 34.775 43.555 38.305 ;
  LAYER M1 ;
        RECT 43.305 38.555 43.555 39.565 ;
  LAYER M1 ;
        RECT 43.305 40.655 43.555 44.185 ;
  LAYER M1 ;
        RECT 43.305 44.435 43.555 45.445 ;
  LAYER M1 ;
        RECT 43.305 46.535 43.555 50.065 ;
  LAYER M1 ;
        RECT 43.305 50.315 43.555 51.325 ;
  LAYER M1 ;
        RECT 43.305 52.415 43.555 55.945 ;
  LAYER M1 ;
        RECT 43.305 56.195 43.555 57.205 ;
  LAYER M1 ;
        RECT 43.305 58.295 43.555 59.305 ;
  LAYER M1 ;
        RECT 43.735 34.775 43.985 38.305 ;
  LAYER M1 ;
        RECT 43.735 40.655 43.985 44.185 ;
  LAYER M1 ;
        RECT 43.735 46.535 43.985 50.065 ;
  LAYER M1 ;
        RECT 43.735 52.415 43.985 55.945 ;
  LAYER M1 ;
        RECT 42.875 34.775 43.125 38.305 ;
  LAYER M1 ;
        RECT 42.875 40.655 43.125 44.185 ;
  LAYER M1 ;
        RECT 42.875 46.535 43.125 50.065 ;
  LAYER M1 ;
        RECT 42.875 52.415 43.125 55.945 ;
  LAYER M1 ;
        RECT 42.445 34.775 42.695 38.305 ;
  LAYER M1 ;
        RECT 42.445 38.555 42.695 39.565 ;
  LAYER M1 ;
        RECT 42.445 40.655 42.695 44.185 ;
  LAYER M1 ;
        RECT 42.445 44.435 42.695 45.445 ;
  LAYER M1 ;
        RECT 42.445 46.535 42.695 50.065 ;
  LAYER M1 ;
        RECT 42.445 50.315 42.695 51.325 ;
  LAYER M1 ;
        RECT 42.445 52.415 42.695 55.945 ;
  LAYER M1 ;
        RECT 42.445 56.195 42.695 57.205 ;
  LAYER M1 ;
        RECT 42.445 58.295 42.695 59.305 ;
  LAYER M1 ;
        RECT 42.015 34.775 42.265 38.305 ;
  LAYER M1 ;
        RECT 42.015 40.655 42.265 44.185 ;
  LAYER M1 ;
        RECT 42.015 46.535 42.265 50.065 ;
  LAYER M1 ;
        RECT 42.015 52.415 42.265 55.945 ;
  LAYER M1 ;
        RECT 41.585 34.775 41.835 38.305 ;
  LAYER M1 ;
        RECT 41.585 38.555 41.835 39.565 ;
  LAYER M1 ;
        RECT 41.585 40.655 41.835 44.185 ;
  LAYER M1 ;
        RECT 41.585 44.435 41.835 45.445 ;
  LAYER M1 ;
        RECT 41.585 46.535 41.835 50.065 ;
  LAYER M1 ;
        RECT 41.585 50.315 41.835 51.325 ;
  LAYER M1 ;
        RECT 41.585 52.415 41.835 55.945 ;
  LAYER M1 ;
        RECT 41.585 56.195 41.835 57.205 ;
  LAYER M1 ;
        RECT 41.585 58.295 41.835 59.305 ;
  LAYER M1 ;
        RECT 41.155 34.775 41.405 38.305 ;
  LAYER M1 ;
        RECT 41.155 40.655 41.405 44.185 ;
  LAYER M1 ;
        RECT 41.155 46.535 41.405 50.065 ;
  LAYER M1 ;
        RECT 41.155 52.415 41.405 55.945 ;
  LAYER M1 ;
        RECT 40.725 34.775 40.975 38.305 ;
  LAYER M1 ;
        RECT 40.725 38.555 40.975 39.565 ;
  LAYER M1 ;
        RECT 40.725 40.655 40.975 44.185 ;
  LAYER M1 ;
        RECT 40.725 44.435 40.975 45.445 ;
  LAYER M1 ;
        RECT 40.725 46.535 40.975 50.065 ;
  LAYER M1 ;
        RECT 40.725 50.315 40.975 51.325 ;
  LAYER M1 ;
        RECT 40.725 52.415 40.975 55.945 ;
  LAYER M1 ;
        RECT 40.725 56.195 40.975 57.205 ;
  LAYER M1 ;
        RECT 40.725 58.295 40.975 59.305 ;
  LAYER M1 ;
        RECT 40.295 34.775 40.545 38.305 ;
  LAYER M1 ;
        RECT 40.295 40.655 40.545 44.185 ;
  LAYER M1 ;
        RECT 40.295 46.535 40.545 50.065 ;
  LAYER M1 ;
        RECT 40.295 52.415 40.545 55.945 ;
  LAYER M1 ;
        RECT 39.865 34.775 40.115 38.305 ;
  LAYER M1 ;
        RECT 39.865 38.555 40.115 39.565 ;
  LAYER M1 ;
        RECT 39.865 40.655 40.115 44.185 ;
  LAYER M1 ;
        RECT 39.865 44.435 40.115 45.445 ;
  LAYER M1 ;
        RECT 39.865 46.535 40.115 50.065 ;
  LAYER M1 ;
        RECT 39.865 50.315 40.115 51.325 ;
  LAYER M1 ;
        RECT 39.865 52.415 40.115 55.945 ;
  LAYER M1 ;
        RECT 39.865 56.195 40.115 57.205 ;
  LAYER M1 ;
        RECT 39.865 58.295 40.115 59.305 ;
  LAYER M1 ;
        RECT 39.435 34.775 39.685 38.305 ;
  LAYER M1 ;
        RECT 39.435 40.655 39.685 44.185 ;
  LAYER M1 ;
        RECT 39.435 46.535 39.685 50.065 ;
  LAYER M1 ;
        RECT 39.435 52.415 39.685 55.945 ;
  LAYER M1 ;
        RECT 39.005 34.775 39.255 38.305 ;
  LAYER M1 ;
        RECT 39.005 38.555 39.255 39.565 ;
  LAYER M1 ;
        RECT 39.005 40.655 39.255 44.185 ;
  LAYER M1 ;
        RECT 39.005 44.435 39.255 45.445 ;
  LAYER M1 ;
        RECT 39.005 46.535 39.255 50.065 ;
  LAYER M1 ;
        RECT 39.005 50.315 39.255 51.325 ;
  LAYER M1 ;
        RECT 39.005 52.415 39.255 55.945 ;
  LAYER M1 ;
        RECT 39.005 56.195 39.255 57.205 ;
  LAYER M1 ;
        RECT 39.005 58.295 39.255 59.305 ;
  LAYER M1 ;
        RECT 38.575 34.775 38.825 38.305 ;
  LAYER M1 ;
        RECT 38.575 40.655 38.825 44.185 ;
  LAYER M1 ;
        RECT 38.575 46.535 38.825 50.065 ;
  LAYER M1 ;
        RECT 38.575 52.415 38.825 55.945 ;
  LAYER M1 ;
        RECT 38.145 34.775 38.395 38.305 ;
  LAYER M1 ;
        RECT 38.145 38.555 38.395 39.565 ;
  LAYER M1 ;
        RECT 38.145 40.655 38.395 44.185 ;
  LAYER M1 ;
        RECT 38.145 44.435 38.395 45.445 ;
  LAYER M1 ;
        RECT 38.145 46.535 38.395 50.065 ;
  LAYER M1 ;
        RECT 38.145 50.315 38.395 51.325 ;
  LAYER M1 ;
        RECT 38.145 52.415 38.395 55.945 ;
  LAYER M1 ;
        RECT 38.145 56.195 38.395 57.205 ;
  LAYER M1 ;
        RECT 38.145 58.295 38.395 59.305 ;
  LAYER M1 ;
        RECT 37.715 34.775 37.965 38.305 ;
  LAYER M1 ;
        RECT 37.715 40.655 37.965 44.185 ;
  LAYER M1 ;
        RECT 37.715 46.535 37.965 50.065 ;
  LAYER M1 ;
        RECT 37.715 52.415 37.965 55.945 ;
  LAYER M1 ;
        RECT 37.285 34.775 37.535 38.305 ;
  LAYER M1 ;
        RECT 37.285 38.555 37.535 39.565 ;
  LAYER M1 ;
        RECT 37.285 40.655 37.535 44.185 ;
  LAYER M1 ;
        RECT 37.285 44.435 37.535 45.445 ;
  LAYER M1 ;
        RECT 37.285 46.535 37.535 50.065 ;
  LAYER M1 ;
        RECT 37.285 50.315 37.535 51.325 ;
  LAYER M1 ;
        RECT 37.285 52.415 37.535 55.945 ;
  LAYER M1 ;
        RECT 37.285 56.195 37.535 57.205 ;
  LAYER M1 ;
        RECT 37.285 58.295 37.535 59.305 ;
  LAYER M1 ;
        RECT 36.855 34.775 37.105 38.305 ;
  LAYER M1 ;
        RECT 36.855 40.655 37.105 44.185 ;
  LAYER M1 ;
        RECT 36.855 46.535 37.105 50.065 ;
  LAYER M1 ;
        RECT 36.855 52.415 37.105 55.945 ;
  LAYER M1 ;
        RECT 36.425 34.775 36.675 38.305 ;
  LAYER M1 ;
        RECT 36.425 38.555 36.675 39.565 ;
  LAYER M1 ;
        RECT 36.425 40.655 36.675 44.185 ;
  LAYER M1 ;
        RECT 36.425 44.435 36.675 45.445 ;
  LAYER M1 ;
        RECT 36.425 46.535 36.675 50.065 ;
  LAYER M1 ;
        RECT 36.425 50.315 36.675 51.325 ;
  LAYER M1 ;
        RECT 36.425 52.415 36.675 55.945 ;
  LAYER M1 ;
        RECT 36.425 56.195 36.675 57.205 ;
  LAYER M1 ;
        RECT 36.425 58.295 36.675 59.305 ;
  LAYER M1 ;
        RECT 35.995 34.775 36.245 38.305 ;
  LAYER M1 ;
        RECT 35.995 40.655 36.245 44.185 ;
  LAYER M1 ;
        RECT 35.995 46.535 36.245 50.065 ;
  LAYER M1 ;
        RECT 35.995 52.415 36.245 55.945 ;
  LAYER M1 ;
        RECT 35.565 34.775 35.815 38.305 ;
  LAYER M1 ;
        RECT 35.565 38.555 35.815 39.565 ;
  LAYER M1 ;
        RECT 35.565 40.655 35.815 44.185 ;
  LAYER M1 ;
        RECT 35.565 44.435 35.815 45.445 ;
  LAYER M1 ;
        RECT 35.565 46.535 35.815 50.065 ;
  LAYER M1 ;
        RECT 35.565 50.315 35.815 51.325 ;
  LAYER M1 ;
        RECT 35.565 52.415 35.815 55.945 ;
  LAYER M1 ;
        RECT 35.565 56.195 35.815 57.205 ;
  LAYER M1 ;
        RECT 35.565 58.295 35.815 59.305 ;
  LAYER M1 ;
        RECT 35.135 34.775 35.385 38.305 ;
  LAYER M1 ;
        RECT 35.135 40.655 35.385 44.185 ;
  LAYER M1 ;
        RECT 35.135 46.535 35.385 50.065 ;
  LAYER M1 ;
        RECT 35.135 52.415 35.385 55.945 ;
  LAYER M1 ;
        RECT 34.705 34.775 34.955 38.305 ;
  LAYER M1 ;
        RECT 34.705 38.555 34.955 39.565 ;
  LAYER M1 ;
        RECT 34.705 40.655 34.955 44.185 ;
  LAYER M1 ;
        RECT 34.705 44.435 34.955 45.445 ;
  LAYER M1 ;
        RECT 34.705 46.535 34.955 50.065 ;
  LAYER M1 ;
        RECT 34.705 50.315 34.955 51.325 ;
  LAYER M1 ;
        RECT 34.705 52.415 34.955 55.945 ;
  LAYER M1 ;
        RECT 34.705 56.195 34.955 57.205 ;
  LAYER M1 ;
        RECT 34.705 58.295 34.955 59.305 ;
  LAYER M1 ;
        RECT 34.275 34.775 34.525 38.305 ;
  LAYER M1 ;
        RECT 34.275 40.655 34.525 44.185 ;
  LAYER M1 ;
        RECT 34.275 46.535 34.525 50.065 ;
  LAYER M1 ;
        RECT 34.275 52.415 34.525 55.945 ;
  LAYER M1 ;
        RECT 33.845 34.775 34.095 38.305 ;
  LAYER M1 ;
        RECT 33.845 38.555 34.095 39.565 ;
  LAYER M1 ;
        RECT 33.845 40.655 34.095 44.185 ;
  LAYER M1 ;
        RECT 33.845 44.435 34.095 45.445 ;
  LAYER M1 ;
        RECT 33.845 46.535 34.095 50.065 ;
  LAYER M1 ;
        RECT 33.845 50.315 34.095 51.325 ;
  LAYER M1 ;
        RECT 33.845 52.415 34.095 55.945 ;
  LAYER M1 ;
        RECT 33.845 56.195 34.095 57.205 ;
  LAYER M1 ;
        RECT 33.845 58.295 34.095 59.305 ;
  LAYER M1 ;
        RECT 33.415 34.775 33.665 38.305 ;
  LAYER M1 ;
        RECT 33.415 40.655 33.665 44.185 ;
  LAYER M1 ;
        RECT 33.415 46.535 33.665 50.065 ;
  LAYER M1 ;
        RECT 33.415 52.415 33.665 55.945 ;
  LAYER M1 ;
        RECT 32.985 34.775 33.235 38.305 ;
  LAYER M1 ;
        RECT 32.985 38.555 33.235 39.565 ;
  LAYER M1 ;
        RECT 32.985 40.655 33.235 44.185 ;
  LAYER M1 ;
        RECT 32.985 44.435 33.235 45.445 ;
  LAYER M1 ;
        RECT 32.985 46.535 33.235 50.065 ;
  LAYER M1 ;
        RECT 32.985 50.315 33.235 51.325 ;
  LAYER M1 ;
        RECT 32.985 52.415 33.235 55.945 ;
  LAYER M1 ;
        RECT 32.985 56.195 33.235 57.205 ;
  LAYER M1 ;
        RECT 32.985 58.295 33.235 59.305 ;
  LAYER M1 ;
        RECT 32.555 34.775 32.805 38.305 ;
  LAYER M1 ;
        RECT 32.555 40.655 32.805 44.185 ;
  LAYER M1 ;
        RECT 32.555 46.535 32.805 50.065 ;
  LAYER M1 ;
        RECT 32.555 52.415 32.805 55.945 ;
  LAYER M1 ;
        RECT 32.125 34.775 32.375 38.305 ;
  LAYER M1 ;
        RECT 32.125 38.555 32.375 39.565 ;
  LAYER M1 ;
        RECT 32.125 40.655 32.375 44.185 ;
  LAYER M1 ;
        RECT 32.125 44.435 32.375 45.445 ;
  LAYER M1 ;
        RECT 32.125 46.535 32.375 50.065 ;
  LAYER M1 ;
        RECT 32.125 50.315 32.375 51.325 ;
  LAYER M1 ;
        RECT 32.125 52.415 32.375 55.945 ;
  LAYER M1 ;
        RECT 32.125 56.195 32.375 57.205 ;
  LAYER M1 ;
        RECT 32.125 58.295 32.375 59.305 ;
  LAYER M1 ;
        RECT 31.695 34.775 31.945 38.305 ;
  LAYER M1 ;
        RECT 31.695 40.655 31.945 44.185 ;
  LAYER M1 ;
        RECT 31.695 46.535 31.945 50.065 ;
  LAYER M1 ;
        RECT 31.695 52.415 31.945 55.945 ;
  LAYER M1 ;
        RECT 31.265 34.775 31.515 38.305 ;
  LAYER M1 ;
        RECT 31.265 38.555 31.515 39.565 ;
  LAYER M1 ;
        RECT 31.265 40.655 31.515 44.185 ;
  LAYER M1 ;
        RECT 31.265 44.435 31.515 45.445 ;
  LAYER M1 ;
        RECT 31.265 46.535 31.515 50.065 ;
  LAYER M1 ;
        RECT 31.265 50.315 31.515 51.325 ;
  LAYER M1 ;
        RECT 31.265 52.415 31.515 55.945 ;
  LAYER M1 ;
        RECT 31.265 56.195 31.515 57.205 ;
  LAYER M1 ;
        RECT 31.265 58.295 31.515 59.305 ;
  LAYER M1 ;
        RECT 30.835 34.775 31.085 38.305 ;
  LAYER M1 ;
        RECT 30.835 40.655 31.085 44.185 ;
  LAYER M1 ;
        RECT 30.835 46.535 31.085 50.065 ;
  LAYER M1 ;
        RECT 30.835 52.415 31.085 55.945 ;
  LAYER M1 ;
        RECT 30.405 34.775 30.655 38.305 ;
  LAYER M1 ;
        RECT 30.405 38.555 30.655 39.565 ;
  LAYER M1 ;
        RECT 30.405 40.655 30.655 44.185 ;
  LAYER M1 ;
        RECT 30.405 44.435 30.655 45.445 ;
  LAYER M1 ;
        RECT 30.405 46.535 30.655 50.065 ;
  LAYER M1 ;
        RECT 30.405 50.315 30.655 51.325 ;
  LAYER M1 ;
        RECT 30.405 52.415 30.655 55.945 ;
  LAYER M1 ;
        RECT 30.405 56.195 30.655 57.205 ;
  LAYER M1 ;
        RECT 30.405 58.295 30.655 59.305 ;
  LAYER M1 ;
        RECT 29.975 34.775 30.225 38.305 ;
  LAYER M1 ;
        RECT 29.975 40.655 30.225 44.185 ;
  LAYER M1 ;
        RECT 29.975 46.535 30.225 50.065 ;
  LAYER M1 ;
        RECT 29.975 52.415 30.225 55.945 ;
  LAYER M1 ;
        RECT 29.545 34.775 29.795 38.305 ;
  LAYER M1 ;
        RECT 29.545 38.555 29.795 39.565 ;
  LAYER M1 ;
        RECT 29.545 40.655 29.795 44.185 ;
  LAYER M1 ;
        RECT 29.545 44.435 29.795 45.445 ;
  LAYER M1 ;
        RECT 29.545 46.535 29.795 50.065 ;
  LAYER M1 ;
        RECT 29.545 50.315 29.795 51.325 ;
  LAYER M1 ;
        RECT 29.545 52.415 29.795 55.945 ;
  LAYER M1 ;
        RECT 29.545 56.195 29.795 57.205 ;
  LAYER M1 ;
        RECT 29.545 58.295 29.795 59.305 ;
  LAYER M1 ;
        RECT 29.115 34.775 29.365 38.305 ;
  LAYER M1 ;
        RECT 29.115 40.655 29.365 44.185 ;
  LAYER M1 ;
        RECT 29.115 46.535 29.365 50.065 ;
  LAYER M1 ;
        RECT 29.115 52.415 29.365 55.945 ;
  LAYER M1 ;
        RECT 28.685 34.775 28.935 38.305 ;
  LAYER M1 ;
        RECT 28.685 38.555 28.935 39.565 ;
  LAYER M1 ;
        RECT 28.685 40.655 28.935 44.185 ;
  LAYER M1 ;
        RECT 28.685 44.435 28.935 45.445 ;
  LAYER M1 ;
        RECT 28.685 46.535 28.935 50.065 ;
  LAYER M1 ;
        RECT 28.685 50.315 28.935 51.325 ;
  LAYER M1 ;
        RECT 28.685 52.415 28.935 55.945 ;
  LAYER M1 ;
        RECT 28.685 56.195 28.935 57.205 ;
  LAYER M1 ;
        RECT 28.685 58.295 28.935 59.305 ;
  LAYER M1 ;
        RECT 28.255 34.775 28.505 38.305 ;
  LAYER M1 ;
        RECT 28.255 40.655 28.505 44.185 ;
  LAYER M1 ;
        RECT 28.255 46.535 28.505 50.065 ;
  LAYER M1 ;
        RECT 28.255 52.415 28.505 55.945 ;
  LAYER M1 ;
        RECT 27.825 34.775 28.075 38.305 ;
  LAYER M1 ;
        RECT 27.825 38.555 28.075 39.565 ;
  LAYER M1 ;
        RECT 27.825 40.655 28.075 44.185 ;
  LAYER M1 ;
        RECT 27.825 44.435 28.075 45.445 ;
  LAYER M1 ;
        RECT 27.825 46.535 28.075 50.065 ;
  LAYER M1 ;
        RECT 27.825 50.315 28.075 51.325 ;
  LAYER M1 ;
        RECT 27.825 52.415 28.075 55.945 ;
  LAYER M1 ;
        RECT 27.825 56.195 28.075 57.205 ;
  LAYER M1 ;
        RECT 27.825 58.295 28.075 59.305 ;
  LAYER M1 ;
        RECT 27.395 34.775 27.645 38.305 ;
  LAYER M1 ;
        RECT 27.395 40.655 27.645 44.185 ;
  LAYER M1 ;
        RECT 27.395 46.535 27.645 50.065 ;
  LAYER M1 ;
        RECT 27.395 52.415 27.645 55.945 ;
  LAYER M1 ;
        RECT 26.965 34.775 27.215 38.305 ;
  LAYER M1 ;
        RECT 26.965 38.555 27.215 39.565 ;
  LAYER M1 ;
        RECT 26.965 40.655 27.215 44.185 ;
  LAYER M1 ;
        RECT 26.965 44.435 27.215 45.445 ;
  LAYER M1 ;
        RECT 26.965 46.535 27.215 50.065 ;
  LAYER M1 ;
        RECT 26.965 50.315 27.215 51.325 ;
  LAYER M1 ;
        RECT 26.965 52.415 27.215 55.945 ;
  LAYER M1 ;
        RECT 26.965 56.195 27.215 57.205 ;
  LAYER M1 ;
        RECT 26.965 58.295 27.215 59.305 ;
  LAYER M1 ;
        RECT 26.535 34.775 26.785 38.305 ;
  LAYER M1 ;
        RECT 26.535 40.655 26.785 44.185 ;
  LAYER M1 ;
        RECT 26.535 46.535 26.785 50.065 ;
  LAYER M1 ;
        RECT 26.535 52.415 26.785 55.945 ;
  LAYER M1 ;
        RECT 26.105 34.775 26.355 38.305 ;
  LAYER M1 ;
        RECT 26.105 38.555 26.355 39.565 ;
  LAYER M1 ;
        RECT 26.105 40.655 26.355 44.185 ;
  LAYER M1 ;
        RECT 26.105 44.435 26.355 45.445 ;
  LAYER M1 ;
        RECT 26.105 46.535 26.355 50.065 ;
  LAYER M1 ;
        RECT 26.105 50.315 26.355 51.325 ;
  LAYER M1 ;
        RECT 26.105 52.415 26.355 55.945 ;
  LAYER M1 ;
        RECT 26.105 56.195 26.355 57.205 ;
  LAYER M1 ;
        RECT 26.105 58.295 26.355 59.305 ;
  LAYER M1 ;
        RECT 25.675 34.775 25.925 38.305 ;
  LAYER M1 ;
        RECT 25.675 40.655 25.925 44.185 ;
  LAYER M1 ;
        RECT 25.675 46.535 25.925 50.065 ;
  LAYER M1 ;
        RECT 25.675 52.415 25.925 55.945 ;
  LAYER M1 ;
        RECT 25.245 34.775 25.495 38.305 ;
  LAYER M1 ;
        RECT 25.245 38.555 25.495 39.565 ;
  LAYER M1 ;
        RECT 25.245 40.655 25.495 44.185 ;
  LAYER M1 ;
        RECT 25.245 44.435 25.495 45.445 ;
  LAYER M1 ;
        RECT 25.245 46.535 25.495 50.065 ;
  LAYER M1 ;
        RECT 25.245 50.315 25.495 51.325 ;
  LAYER M1 ;
        RECT 25.245 52.415 25.495 55.945 ;
  LAYER M1 ;
        RECT 25.245 56.195 25.495 57.205 ;
  LAYER M1 ;
        RECT 25.245 58.295 25.495 59.305 ;
  LAYER M1 ;
        RECT 24.815 34.775 25.065 38.305 ;
  LAYER M1 ;
        RECT 24.815 40.655 25.065 44.185 ;
  LAYER M1 ;
        RECT 24.815 46.535 25.065 50.065 ;
  LAYER M1 ;
        RECT 24.815 52.415 25.065 55.945 ;
  LAYER M1 ;
        RECT 24.385 34.775 24.635 38.305 ;
  LAYER M1 ;
        RECT 24.385 38.555 24.635 39.565 ;
  LAYER M1 ;
        RECT 24.385 40.655 24.635 44.185 ;
  LAYER M1 ;
        RECT 24.385 44.435 24.635 45.445 ;
  LAYER M1 ;
        RECT 24.385 46.535 24.635 50.065 ;
  LAYER M1 ;
        RECT 24.385 50.315 24.635 51.325 ;
  LAYER M1 ;
        RECT 24.385 52.415 24.635 55.945 ;
  LAYER M1 ;
        RECT 24.385 56.195 24.635 57.205 ;
  LAYER M1 ;
        RECT 24.385 58.295 24.635 59.305 ;
  LAYER M1 ;
        RECT 23.955 34.775 24.205 38.305 ;
  LAYER M1 ;
        RECT 23.955 40.655 24.205 44.185 ;
  LAYER M1 ;
        RECT 23.955 46.535 24.205 50.065 ;
  LAYER M1 ;
        RECT 23.955 52.415 24.205 55.945 ;
  LAYER M1 ;
        RECT 23.525 34.775 23.775 38.305 ;
  LAYER M1 ;
        RECT 23.525 38.555 23.775 39.565 ;
  LAYER M1 ;
        RECT 23.525 40.655 23.775 44.185 ;
  LAYER M1 ;
        RECT 23.525 44.435 23.775 45.445 ;
  LAYER M1 ;
        RECT 23.525 46.535 23.775 50.065 ;
  LAYER M1 ;
        RECT 23.525 50.315 23.775 51.325 ;
  LAYER M1 ;
        RECT 23.525 52.415 23.775 55.945 ;
  LAYER M1 ;
        RECT 23.525 56.195 23.775 57.205 ;
  LAYER M1 ;
        RECT 23.525 58.295 23.775 59.305 ;
  LAYER M1 ;
        RECT 23.095 34.775 23.345 38.305 ;
  LAYER M1 ;
        RECT 23.095 40.655 23.345 44.185 ;
  LAYER M1 ;
        RECT 23.095 46.535 23.345 50.065 ;
  LAYER M1 ;
        RECT 23.095 52.415 23.345 55.945 ;
  LAYER M2 ;
        RECT 23.48 34.72 43.6 35 ;
  LAYER M2 ;
        RECT 23.48 38.92 43.6 39.2 ;
  LAYER M2 ;
        RECT 23.05 35.14 44.03 35.42 ;
  LAYER M2 ;
        RECT 23.48 40.6 43.6 40.88 ;
  LAYER M2 ;
        RECT 23.48 44.8 43.6 45.08 ;
  LAYER M2 ;
        RECT 23.05 41.02 44.03 41.3 ;
  LAYER M2 ;
        RECT 23.48 46.48 43.6 46.76 ;
  LAYER M2 ;
        RECT 23.48 50.68 43.6 50.96 ;
  LAYER M2 ;
        RECT 23.05 46.9 44.03 47.18 ;
  LAYER M2 ;
        RECT 23.48 52.36 43.6 52.64 ;
  LAYER M2 ;
        RECT 23.48 56.56 43.6 56.84 ;
  LAYER M2 ;
        RECT 23.48 58.66 43.6 58.94 ;
  LAYER M2 ;
        RECT 23.05 52.78 44.03 53.06 ;
  LAYER M3 ;
        RECT 33.83 34.7 34.11 52.66 ;
  LAYER M3 ;
        RECT 33.4 38.9 33.68 56.86 ;
  LAYER M3 ;
        RECT 32.97 35.12 33.25 58.96 ;
  LAYER M1 ;
        RECT 23.525 9.575 23.775 13.105 ;
  LAYER M1 ;
        RECT 23.525 8.315 23.775 9.325 ;
  LAYER M1 ;
        RECT 23.525 3.695 23.775 7.225 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.525 0.335 23.775 1.345 ;
  LAYER M1 ;
        RECT 23.095 9.575 23.345 13.105 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 23.955 9.575 24.205 13.105 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.385 9.575 24.635 13.105 ;
  LAYER M1 ;
        RECT 24.385 8.315 24.635 9.325 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 24.815 9.575 25.065 13.105 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.245 9.575 25.495 13.105 ;
  LAYER M1 ;
        RECT 25.245 8.315 25.495 9.325 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 25.675 9.575 25.925 13.105 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.105 9.575 26.355 13.105 ;
  LAYER M1 ;
        RECT 26.105 8.315 26.355 9.325 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 26.535 9.575 26.785 13.105 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.965 9.575 27.215 13.105 ;
  LAYER M1 ;
        RECT 26.965 8.315 27.215 9.325 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 9.575 27.645 13.105 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 27.825 9.575 28.075 13.105 ;
  LAYER M1 ;
        RECT 27.825 8.315 28.075 9.325 ;
  LAYER M1 ;
        RECT 27.825 3.695 28.075 7.225 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 1.345 ;
  LAYER M1 ;
        RECT 28.255 9.575 28.505 13.105 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 28.685 9.575 28.935 13.105 ;
  LAYER M1 ;
        RECT 28.685 8.315 28.935 9.325 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 29.115 9.575 29.365 13.105 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.545 9.575 29.795 13.105 ;
  LAYER M1 ;
        RECT 29.545 8.315 29.795 9.325 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 9.575 30.225 13.105 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.405 9.575 30.655 13.105 ;
  LAYER M1 ;
        RECT 30.405 8.315 30.655 9.325 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 30.835 9.575 31.085 13.105 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 31.265 9.575 31.515 13.105 ;
  LAYER M1 ;
        RECT 31.265 8.315 31.515 9.325 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 31.695 9.575 31.945 13.105 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 32.125 9.575 32.375 13.105 ;
  LAYER M1 ;
        RECT 32.125 8.315 32.375 9.325 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 9.575 32.805 13.105 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.985 9.575 33.235 13.105 ;
  LAYER M1 ;
        RECT 32.985 8.315 33.235 9.325 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 9.575 33.665 13.105 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 33.845 9.575 34.095 13.105 ;
  LAYER M1 ;
        RECT 33.845 8.315 34.095 9.325 ;
  LAYER M1 ;
        RECT 33.845 3.695 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.845 2.435 34.095 3.445 ;
  LAYER M1 ;
        RECT 33.845 0.335 34.095 1.345 ;
  LAYER M1 ;
        RECT 34.275 9.575 34.525 13.105 ;
  LAYER M1 ;
        RECT 34.275 3.695 34.525 7.225 ;
  LAYER M1 ;
        RECT 34.705 9.575 34.955 13.105 ;
  LAYER M1 ;
        RECT 34.705 8.315 34.955 9.325 ;
  LAYER M1 ;
        RECT 34.705 3.695 34.955 7.225 ;
  LAYER M1 ;
        RECT 34.705 2.435 34.955 3.445 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 1.345 ;
  LAYER M1 ;
        RECT 35.135 9.575 35.385 13.105 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M2 ;
        RECT 23.48 12.88 35 13.16 ;
  LAYER M2 ;
        RECT 23.48 8.68 35 8.96 ;
  LAYER M2 ;
        RECT 23.05 12.46 35.43 12.74 ;
  LAYER M2 ;
        RECT 23.48 7 35 7.28 ;
  LAYER M2 ;
        RECT 23.48 2.8 35 3.08 ;
  LAYER M2 ;
        RECT 23.48 0.7 35 0.98 ;
  LAYER M2 ;
        RECT 23.05 6.58 35.43 6.86 ;
  LAYER M3 ;
        RECT 28.67 6.98 28.95 13.18 ;
  LAYER M3 ;
        RECT 29.1 2.78 29.38 8.98 ;
  LAYER M3 ;
        RECT 29.53 0.68 29.81 12.76 ;
  LAYER M1 ;
        RECT 14.925 30.575 15.175 34.105 ;
  LAYER M1 ;
        RECT 14.925 29.315 15.175 30.325 ;
  LAYER M1 ;
        RECT 14.925 24.695 15.175 28.225 ;
  LAYER M1 ;
        RECT 14.925 23.435 15.175 24.445 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 22.345 ;
  LAYER M1 ;
        RECT 15.355 30.575 15.605 34.105 ;
  LAYER M1 ;
        RECT 15.355 24.695 15.605 28.225 ;
  LAYER M1 ;
        RECT 14.495 30.575 14.745 34.105 ;
  LAYER M1 ;
        RECT 14.495 24.695 14.745 28.225 ;
  LAYER M1 ;
        RECT 14.065 30.575 14.315 34.105 ;
  LAYER M1 ;
        RECT 14.065 29.315 14.315 30.325 ;
  LAYER M1 ;
        RECT 14.065 24.695 14.315 28.225 ;
  LAYER M1 ;
        RECT 14.065 23.435 14.315 24.445 ;
  LAYER M1 ;
        RECT 14.065 21.335 14.315 22.345 ;
  LAYER M1 ;
        RECT 13.635 30.575 13.885 34.105 ;
  LAYER M1 ;
        RECT 13.635 24.695 13.885 28.225 ;
  LAYER M1 ;
        RECT 13.205 30.575 13.455 34.105 ;
  LAYER M1 ;
        RECT 13.205 29.315 13.455 30.325 ;
  LAYER M1 ;
        RECT 13.205 24.695 13.455 28.225 ;
  LAYER M1 ;
        RECT 13.205 23.435 13.455 24.445 ;
  LAYER M1 ;
        RECT 13.205 21.335 13.455 22.345 ;
  LAYER M1 ;
        RECT 12.775 30.575 13.025 34.105 ;
  LAYER M1 ;
        RECT 12.775 24.695 13.025 28.225 ;
  LAYER M1 ;
        RECT 12.345 30.575 12.595 34.105 ;
  LAYER M1 ;
        RECT 12.345 29.315 12.595 30.325 ;
  LAYER M1 ;
        RECT 12.345 24.695 12.595 28.225 ;
  LAYER M1 ;
        RECT 12.345 23.435 12.595 24.445 ;
  LAYER M1 ;
        RECT 12.345 21.335 12.595 22.345 ;
  LAYER M1 ;
        RECT 11.915 30.575 12.165 34.105 ;
  LAYER M1 ;
        RECT 11.915 24.695 12.165 28.225 ;
  LAYER M1 ;
        RECT 11.485 30.575 11.735 34.105 ;
  LAYER M1 ;
        RECT 11.485 29.315 11.735 30.325 ;
  LAYER M1 ;
        RECT 11.485 24.695 11.735 28.225 ;
  LAYER M1 ;
        RECT 11.485 23.435 11.735 24.445 ;
  LAYER M1 ;
        RECT 11.485 21.335 11.735 22.345 ;
  LAYER M1 ;
        RECT 11.055 30.575 11.305 34.105 ;
  LAYER M1 ;
        RECT 11.055 24.695 11.305 28.225 ;
  LAYER M1 ;
        RECT 10.625 30.575 10.875 34.105 ;
  LAYER M1 ;
        RECT 10.625 29.315 10.875 30.325 ;
  LAYER M1 ;
        RECT 10.625 24.695 10.875 28.225 ;
  LAYER M1 ;
        RECT 10.625 23.435 10.875 24.445 ;
  LAYER M1 ;
        RECT 10.625 21.335 10.875 22.345 ;
  LAYER M1 ;
        RECT 10.195 30.575 10.445 34.105 ;
  LAYER M1 ;
        RECT 10.195 24.695 10.445 28.225 ;
  LAYER M1 ;
        RECT 9.765 30.575 10.015 34.105 ;
  LAYER M1 ;
        RECT 9.765 29.315 10.015 30.325 ;
  LAYER M1 ;
        RECT 9.765 24.695 10.015 28.225 ;
  LAYER M1 ;
        RECT 9.765 23.435 10.015 24.445 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 22.345 ;
  LAYER M1 ;
        RECT 9.335 30.575 9.585 34.105 ;
  LAYER M1 ;
        RECT 9.335 24.695 9.585 28.225 ;
  LAYER M1 ;
        RECT 8.905 30.575 9.155 34.105 ;
  LAYER M1 ;
        RECT 8.905 29.315 9.155 30.325 ;
  LAYER M1 ;
        RECT 8.905 24.695 9.155 28.225 ;
  LAYER M1 ;
        RECT 8.905 23.435 9.155 24.445 ;
  LAYER M1 ;
        RECT 8.905 21.335 9.155 22.345 ;
  LAYER M1 ;
        RECT 8.475 30.575 8.725 34.105 ;
  LAYER M1 ;
        RECT 8.475 24.695 8.725 28.225 ;
  LAYER M1 ;
        RECT 8.045 30.575 8.295 34.105 ;
  LAYER M1 ;
        RECT 8.045 29.315 8.295 30.325 ;
  LAYER M1 ;
        RECT 8.045 24.695 8.295 28.225 ;
  LAYER M1 ;
        RECT 8.045 23.435 8.295 24.445 ;
  LAYER M1 ;
        RECT 8.045 21.335 8.295 22.345 ;
  LAYER M1 ;
        RECT 7.615 30.575 7.865 34.105 ;
  LAYER M1 ;
        RECT 7.615 24.695 7.865 28.225 ;
  LAYER M1 ;
        RECT 7.185 30.575 7.435 34.105 ;
  LAYER M1 ;
        RECT 7.185 29.315 7.435 30.325 ;
  LAYER M1 ;
        RECT 7.185 24.695 7.435 28.225 ;
  LAYER M1 ;
        RECT 7.185 23.435 7.435 24.445 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 22.345 ;
  LAYER M1 ;
        RECT 6.755 30.575 7.005 34.105 ;
  LAYER M1 ;
        RECT 6.755 24.695 7.005 28.225 ;
  LAYER M1 ;
        RECT 6.325 30.575 6.575 34.105 ;
  LAYER M1 ;
        RECT 6.325 29.315 6.575 30.325 ;
  LAYER M1 ;
        RECT 6.325 24.695 6.575 28.225 ;
  LAYER M1 ;
        RECT 6.325 23.435 6.575 24.445 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 22.345 ;
  LAYER M1 ;
        RECT 5.895 30.575 6.145 34.105 ;
  LAYER M1 ;
        RECT 5.895 24.695 6.145 28.225 ;
  LAYER M1 ;
        RECT 5.465 30.575 5.715 34.105 ;
  LAYER M1 ;
        RECT 5.465 29.315 5.715 30.325 ;
  LAYER M1 ;
        RECT 5.465 24.695 5.715 28.225 ;
  LAYER M1 ;
        RECT 5.465 23.435 5.715 24.445 ;
  LAYER M1 ;
        RECT 5.465 21.335 5.715 22.345 ;
  LAYER M1 ;
        RECT 5.035 30.575 5.285 34.105 ;
  LAYER M1 ;
        RECT 5.035 24.695 5.285 28.225 ;
  LAYER M1 ;
        RECT 4.605 30.575 4.855 34.105 ;
  LAYER M1 ;
        RECT 4.605 29.315 4.855 30.325 ;
  LAYER M1 ;
        RECT 4.605 24.695 4.855 28.225 ;
  LAYER M1 ;
        RECT 4.605 23.435 4.855 24.445 ;
  LAYER M1 ;
        RECT 4.605 21.335 4.855 22.345 ;
  LAYER M1 ;
        RECT 4.175 30.575 4.425 34.105 ;
  LAYER M1 ;
        RECT 4.175 24.695 4.425 28.225 ;
  LAYER M1 ;
        RECT 3.745 30.575 3.995 34.105 ;
  LAYER M1 ;
        RECT 3.745 29.315 3.995 30.325 ;
  LAYER M1 ;
        RECT 3.745 24.695 3.995 28.225 ;
  LAYER M1 ;
        RECT 3.745 23.435 3.995 24.445 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.315 30.575 3.565 34.105 ;
  LAYER M1 ;
        RECT 3.315 24.695 3.565 28.225 ;
  LAYER M1 ;
        RECT 2.885 30.575 3.135 34.105 ;
  LAYER M1 ;
        RECT 2.885 29.315 3.135 30.325 ;
  LAYER M1 ;
        RECT 2.885 24.695 3.135 28.225 ;
  LAYER M1 ;
        RECT 2.885 23.435 3.135 24.445 ;
  LAYER M1 ;
        RECT 2.885 21.335 3.135 22.345 ;
  LAYER M1 ;
        RECT 2.455 30.575 2.705 34.105 ;
  LAYER M1 ;
        RECT 2.455 24.695 2.705 28.225 ;
  LAYER M2 ;
        RECT 2.84 33.88 15.22 34.16 ;
  LAYER M2 ;
        RECT 2.84 29.68 15.22 29.96 ;
  LAYER M2 ;
        RECT 2.41 33.46 15.65 33.74 ;
  LAYER M2 ;
        RECT 2.84 28 15.22 28.28 ;
  LAYER M2 ;
        RECT 2.84 23.8 15.22 24.08 ;
  LAYER M2 ;
        RECT 2.84 21.7 15.22 21.98 ;
  LAYER M2 ;
        RECT 2.41 27.58 15.65 27.86 ;
  LAYER M3 ;
        RECT 9.32 27.98 9.6 34.18 ;
  LAYER M3 ;
        RECT 8.89 23.78 9.17 29.98 ;
  LAYER M3 ;
        RECT 8.46 21.68 8.74 33.76 ;
  LAYER M1 ;
        RECT 29.545 30.575 29.795 34.105 ;
  LAYER M1 ;
        RECT 29.545 29.315 29.795 30.325 ;
  LAYER M1 ;
        RECT 29.545 24.695 29.795 28.225 ;
  LAYER M1 ;
        RECT 29.545 23.435 29.795 24.445 ;
  LAYER M1 ;
        RECT 29.545 21.335 29.795 22.345 ;
  LAYER M1 ;
        RECT 29.115 30.575 29.365 34.105 ;
  LAYER M1 ;
        RECT 29.115 24.695 29.365 28.225 ;
  LAYER M1 ;
        RECT 29.975 30.575 30.225 34.105 ;
  LAYER M1 ;
        RECT 29.975 24.695 30.225 28.225 ;
  LAYER M1 ;
        RECT 30.405 30.575 30.655 34.105 ;
  LAYER M1 ;
        RECT 30.405 29.315 30.655 30.325 ;
  LAYER M1 ;
        RECT 30.405 24.695 30.655 28.225 ;
  LAYER M1 ;
        RECT 30.405 23.435 30.655 24.445 ;
  LAYER M1 ;
        RECT 30.405 21.335 30.655 22.345 ;
  LAYER M1 ;
        RECT 30.835 30.575 31.085 34.105 ;
  LAYER M1 ;
        RECT 30.835 24.695 31.085 28.225 ;
  LAYER M1 ;
        RECT 31.265 30.575 31.515 34.105 ;
  LAYER M1 ;
        RECT 31.265 29.315 31.515 30.325 ;
  LAYER M1 ;
        RECT 31.265 24.695 31.515 28.225 ;
  LAYER M1 ;
        RECT 31.265 23.435 31.515 24.445 ;
  LAYER M1 ;
        RECT 31.265 21.335 31.515 22.345 ;
  LAYER M1 ;
        RECT 31.695 30.575 31.945 34.105 ;
  LAYER M1 ;
        RECT 31.695 24.695 31.945 28.225 ;
  LAYER M1 ;
        RECT 32.125 30.575 32.375 34.105 ;
  LAYER M1 ;
        RECT 32.125 29.315 32.375 30.325 ;
  LAYER M1 ;
        RECT 32.125 24.695 32.375 28.225 ;
  LAYER M1 ;
        RECT 32.125 23.435 32.375 24.445 ;
  LAYER M1 ;
        RECT 32.125 21.335 32.375 22.345 ;
  LAYER M1 ;
        RECT 32.555 30.575 32.805 34.105 ;
  LAYER M1 ;
        RECT 32.555 24.695 32.805 28.225 ;
  LAYER M1 ;
        RECT 32.985 30.575 33.235 34.105 ;
  LAYER M1 ;
        RECT 32.985 29.315 33.235 30.325 ;
  LAYER M1 ;
        RECT 32.985 24.695 33.235 28.225 ;
  LAYER M1 ;
        RECT 32.985 23.435 33.235 24.445 ;
  LAYER M1 ;
        RECT 32.985 21.335 33.235 22.345 ;
  LAYER M1 ;
        RECT 33.415 30.575 33.665 34.105 ;
  LAYER M1 ;
        RECT 33.415 24.695 33.665 28.225 ;
  LAYER M1 ;
        RECT 33.845 30.575 34.095 34.105 ;
  LAYER M1 ;
        RECT 33.845 29.315 34.095 30.325 ;
  LAYER M1 ;
        RECT 33.845 24.695 34.095 28.225 ;
  LAYER M1 ;
        RECT 33.845 23.435 34.095 24.445 ;
  LAYER M1 ;
        RECT 33.845 21.335 34.095 22.345 ;
  LAYER M1 ;
        RECT 34.275 30.575 34.525 34.105 ;
  LAYER M1 ;
        RECT 34.275 24.695 34.525 28.225 ;
  LAYER M1 ;
        RECT 34.705 30.575 34.955 34.105 ;
  LAYER M1 ;
        RECT 34.705 29.315 34.955 30.325 ;
  LAYER M1 ;
        RECT 34.705 24.695 34.955 28.225 ;
  LAYER M1 ;
        RECT 34.705 23.435 34.955 24.445 ;
  LAYER M1 ;
        RECT 34.705 21.335 34.955 22.345 ;
  LAYER M1 ;
        RECT 35.135 30.575 35.385 34.105 ;
  LAYER M1 ;
        RECT 35.135 24.695 35.385 28.225 ;
  LAYER M1 ;
        RECT 35.565 30.575 35.815 34.105 ;
  LAYER M1 ;
        RECT 35.565 29.315 35.815 30.325 ;
  LAYER M1 ;
        RECT 35.565 24.695 35.815 28.225 ;
  LAYER M1 ;
        RECT 35.565 23.435 35.815 24.445 ;
  LAYER M1 ;
        RECT 35.565 21.335 35.815 22.345 ;
  LAYER M1 ;
        RECT 35.995 30.575 36.245 34.105 ;
  LAYER M1 ;
        RECT 35.995 24.695 36.245 28.225 ;
  LAYER M1 ;
        RECT 36.425 30.575 36.675 34.105 ;
  LAYER M1 ;
        RECT 36.425 29.315 36.675 30.325 ;
  LAYER M1 ;
        RECT 36.425 24.695 36.675 28.225 ;
  LAYER M1 ;
        RECT 36.425 23.435 36.675 24.445 ;
  LAYER M1 ;
        RECT 36.425 21.335 36.675 22.345 ;
  LAYER M1 ;
        RECT 36.855 30.575 37.105 34.105 ;
  LAYER M1 ;
        RECT 36.855 24.695 37.105 28.225 ;
  LAYER M1 ;
        RECT 37.285 30.575 37.535 34.105 ;
  LAYER M1 ;
        RECT 37.285 29.315 37.535 30.325 ;
  LAYER M1 ;
        RECT 37.285 24.695 37.535 28.225 ;
  LAYER M1 ;
        RECT 37.285 23.435 37.535 24.445 ;
  LAYER M1 ;
        RECT 37.285 21.335 37.535 22.345 ;
  LAYER M1 ;
        RECT 37.715 30.575 37.965 34.105 ;
  LAYER M1 ;
        RECT 37.715 24.695 37.965 28.225 ;
  LAYER M1 ;
        RECT 38.145 30.575 38.395 34.105 ;
  LAYER M1 ;
        RECT 38.145 29.315 38.395 30.325 ;
  LAYER M1 ;
        RECT 38.145 24.695 38.395 28.225 ;
  LAYER M1 ;
        RECT 38.145 23.435 38.395 24.445 ;
  LAYER M1 ;
        RECT 38.145 21.335 38.395 22.345 ;
  LAYER M1 ;
        RECT 38.575 30.575 38.825 34.105 ;
  LAYER M1 ;
        RECT 38.575 24.695 38.825 28.225 ;
  LAYER M1 ;
        RECT 39.005 30.575 39.255 34.105 ;
  LAYER M1 ;
        RECT 39.005 29.315 39.255 30.325 ;
  LAYER M1 ;
        RECT 39.005 24.695 39.255 28.225 ;
  LAYER M1 ;
        RECT 39.005 23.435 39.255 24.445 ;
  LAYER M1 ;
        RECT 39.005 21.335 39.255 22.345 ;
  LAYER M1 ;
        RECT 39.435 30.575 39.685 34.105 ;
  LAYER M1 ;
        RECT 39.435 24.695 39.685 28.225 ;
  LAYER M1 ;
        RECT 39.865 30.575 40.115 34.105 ;
  LAYER M1 ;
        RECT 39.865 29.315 40.115 30.325 ;
  LAYER M1 ;
        RECT 39.865 24.695 40.115 28.225 ;
  LAYER M1 ;
        RECT 39.865 23.435 40.115 24.445 ;
  LAYER M1 ;
        RECT 39.865 21.335 40.115 22.345 ;
  LAYER M1 ;
        RECT 40.295 30.575 40.545 34.105 ;
  LAYER M1 ;
        RECT 40.295 24.695 40.545 28.225 ;
  LAYER M1 ;
        RECT 40.725 30.575 40.975 34.105 ;
  LAYER M1 ;
        RECT 40.725 29.315 40.975 30.325 ;
  LAYER M1 ;
        RECT 40.725 24.695 40.975 28.225 ;
  LAYER M1 ;
        RECT 40.725 23.435 40.975 24.445 ;
  LAYER M1 ;
        RECT 40.725 21.335 40.975 22.345 ;
  LAYER M1 ;
        RECT 41.155 30.575 41.405 34.105 ;
  LAYER M1 ;
        RECT 41.155 24.695 41.405 28.225 ;
  LAYER M1 ;
        RECT 41.585 30.575 41.835 34.105 ;
  LAYER M1 ;
        RECT 41.585 29.315 41.835 30.325 ;
  LAYER M1 ;
        RECT 41.585 24.695 41.835 28.225 ;
  LAYER M1 ;
        RECT 41.585 23.435 41.835 24.445 ;
  LAYER M1 ;
        RECT 41.585 21.335 41.835 22.345 ;
  LAYER M1 ;
        RECT 42.015 30.575 42.265 34.105 ;
  LAYER M1 ;
        RECT 42.015 24.695 42.265 28.225 ;
  LAYER M2 ;
        RECT 29.5 33.88 41.88 34.16 ;
  LAYER M2 ;
        RECT 29.5 29.68 41.88 29.96 ;
  LAYER M2 ;
        RECT 29.07 33.46 42.31 33.74 ;
  LAYER M2 ;
        RECT 29.5 28 41.88 28.28 ;
  LAYER M2 ;
        RECT 29.5 23.8 41.88 24.08 ;
  LAYER M2 ;
        RECT 29.5 21.7 41.88 21.98 ;
  LAYER M2 ;
        RECT 29.07 27.58 42.31 27.86 ;
  LAYER M3 ;
        RECT 35.12 27.98 35.4 34.18 ;
  LAYER M3 ;
        RECT 35.55 23.78 35.83 29.98 ;
  LAYER M3 ;
        RECT 35.98 21.68 36.26 33.76 ;
  LAYER M1 ;
        RECT 9.765 17.135 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.765 15.875 10.015 16.885 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.335 17.135 9.585 20.665 ;
  LAYER M1 ;
        RECT 10.195 17.135 10.445 20.665 ;
  LAYER M1 ;
        RECT 10.625 17.135 10.875 20.665 ;
  LAYER M1 ;
        RECT 10.625 15.875 10.875 16.885 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 17.135 11.305 20.665 ;
  LAYER M1 ;
        RECT 11.485 17.135 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.485 15.875 11.735 16.885 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 17.135 12.165 20.665 ;
  LAYER M1 ;
        RECT 12.345 17.135 12.595 20.665 ;
  LAYER M1 ;
        RECT 12.345 15.875 12.595 16.885 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 14.785 ;
  LAYER M1 ;
        RECT 12.775 17.135 13.025 20.665 ;
  LAYER M1 ;
        RECT 13.205 17.135 13.455 20.665 ;
  LAYER M1 ;
        RECT 13.205 15.875 13.455 16.885 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.635 17.135 13.885 20.665 ;
  LAYER M1 ;
        RECT 14.065 17.135 14.315 20.665 ;
  LAYER M1 ;
        RECT 14.065 15.875 14.315 16.885 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.495 17.135 14.745 20.665 ;
  LAYER M1 ;
        RECT 14.925 17.135 15.175 20.665 ;
  LAYER M1 ;
        RECT 14.925 15.875 15.175 16.885 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 14.785 ;
  LAYER M1 ;
        RECT 15.355 17.135 15.605 20.665 ;
  LAYER M1 ;
        RECT 15.785 17.135 16.035 20.665 ;
  LAYER M1 ;
        RECT 15.785 15.875 16.035 16.885 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 14.785 ;
  LAYER M1 ;
        RECT 16.215 17.135 16.465 20.665 ;
  LAYER M1 ;
        RECT 16.645 17.135 16.895 20.665 ;
  LAYER M1 ;
        RECT 16.645 15.875 16.895 16.885 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 17.075 17.135 17.325 20.665 ;
  LAYER M1 ;
        RECT 17.505 17.135 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.505 15.875 17.755 16.885 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.935 17.135 18.185 20.665 ;
  LAYER M1 ;
        RECT 18.365 17.135 18.615 20.665 ;
  LAYER M1 ;
        RECT 18.365 15.875 18.615 16.885 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 14.785 ;
  LAYER M1 ;
        RECT 18.795 17.135 19.045 20.665 ;
  LAYER M1 ;
        RECT 19.225 17.135 19.475 20.665 ;
  LAYER M1 ;
        RECT 19.225 15.875 19.475 16.885 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 19.655 17.135 19.905 20.665 ;
  LAYER M1 ;
        RECT 20.085 17.135 20.335 20.665 ;
  LAYER M1 ;
        RECT 20.085 15.875 20.335 16.885 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 14.785 ;
  LAYER M1 ;
        RECT 20.515 17.135 20.765 20.665 ;
  LAYER M1 ;
        RECT 20.945 17.135 21.195 20.665 ;
  LAYER M1 ;
        RECT 20.945 15.875 21.195 16.885 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 14.785 ;
  LAYER M1 ;
        RECT 21.375 17.135 21.625 20.665 ;
  LAYER M2 ;
        RECT 9.72 14.14 21.24 14.42 ;
  LAYER M2 ;
        RECT 9.72 20.44 21.24 20.72 ;
  LAYER M2 ;
        RECT 9.72 16.24 21.24 16.52 ;
  LAYER M2 ;
        RECT 9.29 20.02 21.67 20.3 ;
  LAYER M1 ;
        RECT 34.705 17.135 34.955 20.665 ;
  LAYER M1 ;
        RECT 34.705 15.875 34.955 16.885 ;
  LAYER M1 ;
        RECT 34.705 13.775 34.955 14.785 ;
  LAYER M1 ;
        RECT 35.135 17.135 35.385 20.665 ;
  LAYER M1 ;
        RECT 34.275 17.135 34.525 20.665 ;
  LAYER M1 ;
        RECT 33.845 17.135 34.095 20.665 ;
  LAYER M1 ;
        RECT 33.845 15.875 34.095 16.885 ;
  LAYER M1 ;
        RECT 33.845 13.775 34.095 14.785 ;
  LAYER M1 ;
        RECT 33.415 17.135 33.665 20.665 ;
  LAYER M1 ;
        RECT 32.985 17.135 33.235 20.665 ;
  LAYER M1 ;
        RECT 32.985 15.875 33.235 16.885 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 14.785 ;
  LAYER M1 ;
        RECT 32.555 17.135 32.805 20.665 ;
  LAYER M1 ;
        RECT 32.125 17.135 32.375 20.665 ;
  LAYER M1 ;
        RECT 32.125 15.875 32.375 16.885 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 14.785 ;
  LAYER M1 ;
        RECT 31.695 17.135 31.945 20.665 ;
  LAYER M1 ;
        RECT 31.265 17.135 31.515 20.665 ;
  LAYER M1 ;
        RECT 31.265 15.875 31.515 16.885 ;
  LAYER M1 ;
        RECT 31.265 13.775 31.515 14.785 ;
  LAYER M1 ;
        RECT 30.835 17.135 31.085 20.665 ;
  LAYER M1 ;
        RECT 30.405 17.135 30.655 20.665 ;
  LAYER M1 ;
        RECT 30.405 15.875 30.655 16.885 ;
  LAYER M1 ;
        RECT 30.405 13.775 30.655 14.785 ;
  LAYER M1 ;
        RECT 29.975 17.135 30.225 20.665 ;
  LAYER M1 ;
        RECT 29.545 17.135 29.795 20.665 ;
  LAYER M1 ;
        RECT 29.545 15.875 29.795 16.885 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.115 17.135 29.365 20.665 ;
  LAYER M1 ;
        RECT 28.685 17.135 28.935 20.665 ;
  LAYER M1 ;
        RECT 28.685 15.875 28.935 16.885 ;
  LAYER M1 ;
        RECT 28.685 13.775 28.935 14.785 ;
  LAYER M1 ;
        RECT 28.255 17.135 28.505 20.665 ;
  LAYER M1 ;
        RECT 27.825 17.135 28.075 20.665 ;
  LAYER M1 ;
        RECT 27.825 15.875 28.075 16.885 ;
  LAYER M1 ;
        RECT 27.825 13.775 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.395 17.135 27.645 20.665 ;
  LAYER M1 ;
        RECT 26.965 17.135 27.215 20.665 ;
  LAYER M1 ;
        RECT 26.965 15.875 27.215 16.885 ;
  LAYER M1 ;
        RECT 26.965 13.775 27.215 14.785 ;
  LAYER M1 ;
        RECT 26.535 17.135 26.785 20.665 ;
  LAYER M1 ;
        RECT 26.105 17.135 26.355 20.665 ;
  LAYER M1 ;
        RECT 26.105 15.875 26.355 16.885 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 14.785 ;
  LAYER M1 ;
        RECT 25.675 17.135 25.925 20.665 ;
  LAYER M1 ;
        RECT 25.245 17.135 25.495 20.665 ;
  LAYER M1 ;
        RECT 25.245 15.875 25.495 16.885 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 14.785 ;
  LAYER M1 ;
        RECT 24.815 17.135 25.065 20.665 ;
  LAYER M1 ;
        RECT 24.385 17.135 24.635 20.665 ;
  LAYER M1 ;
        RECT 24.385 15.875 24.635 16.885 ;
  LAYER M1 ;
        RECT 24.385 13.775 24.635 14.785 ;
  LAYER M1 ;
        RECT 23.955 17.135 24.205 20.665 ;
  LAYER M1 ;
        RECT 23.525 17.135 23.775 20.665 ;
  LAYER M1 ;
        RECT 23.525 15.875 23.775 16.885 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 14.785 ;
  LAYER M1 ;
        RECT 23.095 17.135 23.345 20.665 ;
  LAYER M2 ;
        RECT 23.48 14.14 35 14.42 ;
  LAYER M2 ;
        RECT 23.48 20.44 35 20.72 ;
  LAYER M2 ;
        RECT 23.48 16.24 35 16.52 ;
  LAYER M2 ;
        RECT 23.05 20.02 35.43 20.3 ;
  END 
END CURRENT_MIRROR_OTA
