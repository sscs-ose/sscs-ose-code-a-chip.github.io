* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
X0 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=250000u
X1 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=150000u
X2 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=250000u
X3 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=150000u
.ends
