MACRO NMOS_S_17321006_X28_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_17321006_X28_Y1 0 0 ;
  SIZE 25800 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 280 24680 560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 4480 24680 4760 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 13190 680 13470 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 7225 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 7225 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 7225 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 7225 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 7225 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 7225 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 7225 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 7225 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 7225 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 7225 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 7225 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 7225 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 7225 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 7225 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 7225 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 7225 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 7225 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 7225 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 7225 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 20085 335 20335 3865 ;
    LAYER M1 ;
      RECT 20085 4115 20335 5125 ;
    LAYER M1 ;
      RECT 20085 6215 20335 7225 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20945 335 21195 3865 ;
    LAYER M1 ;
      RECT 20945 4115 21195 5125 ;
    LAYER M1 ;
      RECT 20945 6215 21195 7225 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 21805 335 22055 3865 ;
    LAYER M1 ;
      RECT 21805 4115 22055 5125 ;
    LAYER M1 ;
      RECT 21805 6215 22055 7225 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22665 335 22915 3865 ;
    LAYER M1 ;
      RECT 22665 4115 22915 5125 ;
    LAYER M1 ;
      RECT 22665 6215 22915 7225 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23525 335 23775 3865 ;
    LAYER M1 ;
      RECT 23525 4115 23775 5125 ;
    LAYER M1 ;
      RECT 23525 6215 23775 7225 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 24385 335 24635 3865 ;
    LAYER M1 ;
      RECT 24385 4115 24635 5125 ;
    LAYER M1 ;
      RECT 24385 6215 24635 7225 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M2 ;
      RECT 1120 6580 24680 6860 ;
    LAYER M2 ;
      RECT 690 700 25110 980 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6635 3955 6805 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6635 5675 6805 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6635 6535 6805 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6635 7395 6805 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6635 8255 6805 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6635 9115 6805 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6635 9975 6805 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6635 10835 6805 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6635 11695 6805 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6635 12555 6805 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6635 13415 6805 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6635 14275 6805 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6635 15135 6805 ;
    LAYER V1 ;
      RECT 15825 335 15995 505 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6635 15995 6805 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6635 16855 6805 ;
    LAYER V1 ;
      RECT 17545 335 17715 505 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6635 17715 6805 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6635 18575 6805 ;
    LAYER V1 ;
      RECT 19265 335 19435 505 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6635 19435 6805 ;
    LAYER V1 ;
      RECT 20125 335 20295 505 ;
    LAYER V1 ;
      RECT 20125 4535 20295 4705 ;
    LAYER V1 ;
      RECT 20125 6635 20295 6805 ;
    LAYER V1 ;
      RECT 20985 335 21155 505 ;
    LAYER V1 ;
      RECT 20985 4535 21155 4705 ;
    LAYER V1 ;
      RECT 20985 6635 21155 6805 ;
    LAYER V1 ;
      RECT 21845 335 22015 505 ;
    LAYER V1 ;
      RECT 21845 4535 22015 4705 ;
    LAYER V1 ;
      RECT 21845 6635 22015 6805 ;
    LAYER V1 ;
      RECT 22705 335 22875 505 ;
    LAYER V1 ;
      RECT 22705 4535 22875 4705 ;
    LAYER V1 ;
      RECT 22705 6635 22875 6805 ;
    LAYER V1 ;
      RECT 23565 335 23735 505 ;
    LAYER V1 ;
      RECT 23565 4535 23735 4705 ;
    LAYER V1 ;
      RECT 23565 6635 23735 6805 ;
    LAYER V1 ;
      RECT 24425 335 24595 505 ;
    LAYER V1 ;
      RECT 24425 4535 24595 4705 ;
    LAYER V1 ;
      RECT 24425 6635 24595 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 15395 755 15565 925 ;
    LAYER V1 ;
      RECT 16255 755 16425 925 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17975 755 18145 925 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 19695 755 19865 925 ;
    LAYER V1 ;
      RECT 20555 755 20725 925 ;
    LAYER V1 ;
      RECT 21415 755 21585 925 ;
    LAYER V1 ;
      RECT 22275 755 22445 925 ;
    LAYER V1 ;
      RECT 23135 755 23305 925 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 24855 755 25025 925 ;
    LAYER V2 ;
      RECT 13255 765 13405 915 ;
    LAYER V2 ;
      RECT 13255 6645 13405 6795 ;
  END
END NMOS_S_17321006_X28_Y1
