# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_20v0_noptap_iso
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_20v0_noptap_iso ;
  ORIGIN  12.38000  7.000000 ;
  SIZE  26.26000 BY  44.00500 ;
  OBS
    LAYER li1 ;
      RECT -5.340000  0.045000 -4.670000 29.955000 ;
      RECT -4.150000  0.045000 -3.480000 29.955000 ;
      RECT -1.045000 -3.285000  2.775000 -2.215000 ;
      RECT  0.075000  0.215000  1.425000 29.785000 ;
      RECT  4.980000  0.045000  5.650000 29.955000 ;
      RECT  6.170000  0.045000  6.840000 29.955000 ;
    LAYER mcon ;
      RECT -5.270000  0.155000 -4.740000 29.845000 ;
      RECT -4.080000  0.155000 -3.550000 29.845000 ;
      RECT -0.900000 -3.205000 -0.730000 -3.035000 ;
      RECT -0.900000 -2.835000 -0.730000 -2.665000 ;
      RECT -0.900000 -2.465000 -0.730000 -2.295000 ;
      RECT -0.530000 -3.205000 -0.360000 -3.035000 ;
      RECT -0.530000 -2.835000 -0.360000 -2.665000 ;
      RECT -0.530000 -2.465000 -0.360000 -2.295000 ;
      RECT -0.160000 -3.205000  0.010000 -3.035000 ;
      RECT -0.160000 -2.835000  0.010000 -2.665000 ;
      RECT -0.160000 -2.465000  0.010000 -2.295000 ;
      RECT  0.125000  0.335000  1.375000 29.665000 ;
      RECT  0.210000 -3.205000  0.380000 -3.035000 ;
      RECT  0.210000 -2.835000  0.380000 -2.665000 ;
      RECT  0.210000 -2.465000  0.380000 -2.295000 ;
      RECT  0.580000 -3.205000  0.750000 -3.035000 ;
      RECT  0.580000 -2.835000  0.750000 -2.665000 ;
      RECT  0.580000 -2.465000  0.750000 -2.295000 ;
      RECT  0.950000 -3.205000  1.120000 -3.035000 ;
      RECT  0.950000 -2.835000  1.120000 -2.665000 ;
      RECT  0.950000 -2.465000  1.120000 -2.295000 ;
      RECT  1.320000 -3.205000  1.490000 -3.035000 ;
      RECT  1.320000 -2.835000  1.490000 -2.665000 ;
      RECT  1.320000 -2.465000  1.490000 -2.295000 ;
      RECT  1.690000 -3.205000  1.860000 -3.035000 ;
      RECT  1.690000 -2.835000  1.860000 -2.665000 ;
      RECT  1.690000 -2.465000  1.860000 -2.295000 ;
      RECT  2.060000 -3.205000  2.230000 -3.035000 ;
      RECT  2.060000 -2.835000  2.230000 -2.665000 ;
      RECT  2.060000 -2.465000  2.230000 -2.295000 ;
      RECT  2.430000 -3.205000  2.600000 -3.035000 ;
      RECT  2.430000 -2.835000  2.600000 -2.665000 ;
      RECT  2.430000 -2.465000  2.600000 -2.295000 ;
      RECT  5.050000  0.155000  5.580000 29.845000 ;
      RECT  6.240000  0.155000  6.770000 29.845000 ;
    LAYER met1 ;
      RECT -5.330000  0.095000 -4.680000 29.905000 ;
      RECT -4.140000  0.095000 -3.490000 29.905000 ;
      RECT -1.045000 -3.285000  2.775000 -2.215000 ;
      RECT  0.065000  0.275000  1.435000 29.725000 ;
      RECT  4.990000  0.095000  5.640000 29.905000 ;
      RECT  6.180000  0.095000  6.830000 29.905000 ;
    LAYER met2 ;
      RECT -1.045000 -3.285000 2.775000 -2.215000 ;
      RECT  0.110000  0.285000 1.390000 29.725000 ;
    LAYER via ;
      RECT -0.945000 -3.250000 -0.685000 -2.990000 ;
      RECT -0.945000 -2.880000 -0.685000 -2.620000 ;
      RECT -0.945000 -2.510000 -0.685000 -2.250000 ;
      RECT -0.575000 -3.250000 -0.315000 -2.990000 ;
      RECT -0.575000 -2.880000 -0.315000 -2.620000 ;
      RECT -0.575000 -2.510000 -0.315000 -2.250000 ;
      RECT -0.205000 -3.250000  0.055000 -2.990000 ;
      RECT -0.205000 -2.880000  0.055000 -2.620000 ;
      RECT -0.205000 -2.510000  0.055000 -2.250000 ;
      RECT  0.140000  0.315000  1.360000 29.695000 ;
      RECT  0.165000 -3.250000  0.425000 -2.990000 ;
      RECT  0.165000 -2.880000  0.425000 -2.620000 ;
      RECT  0.165000 -2.510000  0.425000 -2.250000 ;
      RECT  0.535000 -3.250000  0.795000 -2.990000 ;
      RECT  0.535000 -2.880000  0.795000 -2.620000 ;
      RECT  0.535000 -2.510000  0.795000 -2.250000 ;
      RECT  0.905000 -3.250000  1.165000 -2.990000 ;
      RECT  0.905000 -2.880000  1.165000 -2.620000 ;
      RECT  0.905000 -2.510000  1.165000 -2.250000 ;
      RECT  1.275000 -3.250000  1.535000 -2.990000 ;
      RECT  1.275000 -2.880000  1.535000 -2.620000 ;
      RECT  1.275000 -2.510000  1.535000 -2.250000 ;
      RECT  1.645000 -3.250000  1.905000 -2.990000 ;
      RECT  1.645000 -2.880000  1.905000 -2.620000 ;
      RECT  1.645000 -2.510000  1.905000 -2.250000 ;
      RECT  2.015000 -3.250000  2.275000 -2.990000 ;
      RECT  2.015000 -2.880000  2.275000 -2.620000 ;
      RECT  2.015000 -2.510000  2.275000 -2.250000 ;
      RECT  2.385000 -3.250000  2.645000 -2.990000 ;
      RECT  2.385000 -2.880000  2.645000 -2.620000 ;
      RECT  2.385000 -2.510000  2.645000 -2.250000 ;
  END
END sky130_fd_pr__rf_nfet_20v0_noptap_iso
END LIBRARY
