module approxMult_signed8x8 (A, B, OUT);
  input  [7:0] A;
  input  [7:0] B;
  output [15:0] OUT;
  wire n0, n1, n10, n11, n12, n13, n14, n15, n2, n3, n4, n5, n6, n7, n8, n9, v0_0, v100_0, v101_0, v102_0, v103_0, v104_0, v105_0, v106_0, v107_0, v108_0, v109_0, v10_0, v110_0, v111_0, v112_0, v113_0, v114_0, v115_0, v116_0, v117_0, v118_0, v119_0, v11_0, v120_0, v121_0, v122_0, v123_0, v124_0, v125_0, v126_0, v127_0, v128_0, v129_0, v12_0, v130_0, v131_0, v132_0, v133_0, v134_0, v135_0, v136_0, v137_0, v138_0, v139_0, v13_0, v140_0, v141_0, v142_0, v143_0, v144_0, v145_0, v146_0, v147_0, v148_0, v149_0, v14_0, v150_0, v151_0, v152_0, v153_0, v154_0, v155_0, v156_0, v157_0, v158_0, v159_0, v15_0, v160_0, v161_0, v162_0, v163_0, v164_0, v165_0, v166_0, v167_0, v168_0, v169_0, v16_0, v170_0, v171_0, v172_0, v173_0, v174_0, v175_0, v176_0, v177_0, v178_0, v179_0, v17_0, v180_0, v181_0, v182_0, v183_0, v184_0, v185_0, v186_0, v187_0, v188_0, v189_0, v18_0, v190_0, v191_0, v192_0, v193_0, v194_0, v195_0, v196_0, v197_0, v198_0, v199_0, v19_0, v1_0, v200_0, v201_0, v202_0, v203_0, v204_0, v205_0, v206_0, v207_0, v208_0, v209_0, v20_0, v210_0, v211_0, v212_0, v213_0, v214_0, v215_0, v216_0, v217_0, v218_0, v219_0, v21_0, v220_0, v221_0, v222_0, v223_0, v224_0, v225_0, v226_0, v227_0, v228_0, v229_0, v22_0, v230_0, v231_0, v232_0, v233_0, v234_0, v235_0, v236_0, v237_0, v238_0, v239_0, v23_0, v240_0, v241_0, v242_0, v243_0, v244_0, v245_0, v246_0, v247_0, v248_0, v249_0, v24_0, v250_0, v251_0, v252_0, v253_0, v254_0, v255_0, v256_0, v257_0, v258_0, v259_0, v25_0, v260_0, v261_0, v262_0, v263_0, v264_0, v265_0, v266_0, v267_0, v268_0, v269_0, v26_0, v270_0, v271_0, v272_0, v273_0, v274_0, v275_0, v276_0, v277_0, v278_0, v279_0, v27_0, v280_0, v281_0, v282_0, v283_0, v284_0, v285_0, v286_0, v287_0, v288_0, v289_0, v28_0, v290_0, v291_0, v292_0, v293_0, v294_0, v295_0, v296_0, v297_0, v298_0, v299_0, v29_0, v2_0, v300_0, v301_0, v302_0, v303_0, v304_0, v305_0, v306_0, v307_0, v308_0, v309_0, v30_0, v310_0, v311_0, v312_0, v313_0, v314_0, v315_0, v316_0, v317_0, v318_0, v319_0, v31_0, v320_0, v321_0, v322_0, v323_0, v324_0, v325_0, v326_0, v327_0, v328_0, v329_0, v32_0, v330_0, v331_0, v332_0, v333_0, v334_0, v335_0, v336_0, v337_0, v338_0, v339_0, v33_0, v340_0, v341_0, v342_0, v343_0, v344_0, v345_0, v346_0, v347_0, v348_0, v349_0, v34_0, v350_0, v351_0, v352_0, v353_0, v354_0, v355_0, v356_0, v357_0, v358_0, v359_0, v35_0, v360_0, v361_0, v362_0, v363_0, v364_0, v365_0, v366_0, v367_0, v368_0, v369_0, v36_0, v370_0, v371_0, v372_0, v373_0, v374_0, v375_0, v376_0, v377_0, v378_0, v379_0, v37_0, v380_0, v381_0, v382_0, v383_0, v384_0, v385_0, v386_0, v387_0, v388_0, v389_0, v38_0, v390_0, v391_0, v392_0, v393_0, v394_0, v395_0, v396_0, v397_0, v398_0, v399_0, v39_0, v3_0, v400_0, v401_0, v402_0, v403_0, v404_0, v405_0, v406_0, v407_0, v408_0, v409_0, v40_0, v410_0, v411_0, v412_0, v413_0, v414_0, v415_0, v416_0, v417_0, v418_0, v419_0, v41_0, v420_0, v421_0, v422_0, v423_0, v424_0, v425_0, v426_0, v427_0, v428_0, v429_0, v42_0, v430_0, v431_0, v432_0, v433_0, v434_0, v435_0, v436_0, v437_0, v438_0, v439_0, v43_0, v440_0, v441_0, v442_0, v443_0, v444_0, v445_0, v446_0, v447_0, v448_0, v449_0, v44_0, v450_0, v451_0, v452_0, v453_0, v454_0, v455_0, v456_0, v457_0, v458_0, v459_0, v45_0, v460_0, v461_0, v462_0, v463_0, v464_0, v465_0, v466_0, v467_0, v468_0, v469_0, v46_0, v47_0, v48_0, v49_0, v4_0, v50_0, v51_0, v52_0, v53_0, v54_0, v55_0, v56_0, v57_0, v58_0, v59_0, v5_0, v60_0, v61_0, v62_0, v63_0, v64_0, v65_0, v66_0, v67_0, v68_0, v69_0, v6_0, v70_0, v71_0, v72_0, v73_0, v74_0, v75_0, v76_0, v77_0, v78_0, v79_0, v7_0, v80_0, v81_0, v82_0, v83_0, v84_0, v85_0, v86_0, v87_0, v88_0, v89_0, v8_0, v90_0, v91_0, v92_0, v93_0, v94_0, v95_0, v96_0, v97_0, v98_0, v99_0, v9_0;

  // Map n0..n7 to A[0..7], n8..n15 to B[0..7]
  assign n0 = A[0];
  assign n1 = A[1];
  assign n2 = A[2];
  assign n3 = A[3];
  assign n4 = A[4];
  assign n5 = A[5];
  assign n6 = A[6];
  assign n7 = A[7];
  assign n8 = B[0];
  assign n9 = B[1];
  assign n10 = B[2];
  assign n11 = B[3];
  assign n12 = B[4];
  assign n13 = B[5];
  assign n14 = B[6];
  assign n15 = B[7];

  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0001_ (
    .A1(n12),
    .A2(n1),
    .ZN(v0_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0002_ (
    .I(v0_0),
    .ZN(v1_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0003_ (
    .A1(n11),
    .A2(n0),
    .ZN(v2_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0004_ (
    .I(v2_0),
    .ZN(v3_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0005_ (
    .A1(v1_0),
    .A2(v3_0),
    .ZN(v4_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0006_ (
    .I(v4_0),
    .ZN(v5_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0007_ (
    .A1(n9),
    .A2(n3),
    .ZN(v6_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0008_ (
    .A1(n9),
    .A2(n2),
    .ZN(v7_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0009_ (
    .A1(n8),
    .A2(n3),
    .ZN(v8_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0010_ (
    .I(v8_0),
    .ZN(v9_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0011_ (
    .A1(n10),
    .A2(n1),
    .ZN(v10_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0012_ (
    .I(v10_0),
    .ZN(v11_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0013_ (
    .A1(v9_0),
    .A2(v11_0),
    .ZN(v12_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0014_ (
    .I(v12_0),
    .ZN(v13_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0015_ (
    .A1(n10),
    .A2(n2),
    .ZN(v14_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0016_ (
    .A1(n9),
    .A2(n4),
    .ZN(v15_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0017_ (
    .A1(v8_0),
    .A2(v15_0),
    .Z(v16_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0018_ (
    .A1(n8),
    .A2(n4),
    .ZN(v17_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0019_ (
    .A1(v6_0),
    .A2(v17_0),
    .ZN(v18_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0020_ (
    .A1(v16_0),
    .A2(v18_0),
    .ZN(v19_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0021_ (
    .A1(v14_0),
    .A2(v19_0),
    .Z(v20_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0022_ (
    .A1(v13_0),
    .A2(v20_0),
    .Z(v21_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0023_ (
    .A1(n12),
    .A2(n0),
    .ZN(v22_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0024_ (
    .A1(n11),
    .A2(n1),
    .ZN(v23_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0025_ (
    .A1(v22_0),
    .A2(v23_0),
    .Z(v24_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0026_ (
    .A1(v21_0),
    .A2(v24_0),
    .ZN(v25_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0027_ (
    .A1(v20_0),
    .A2(v13_0),
    .ZN(v26_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0028_ (
    .A1(v25_0),
    .A2(v26_0),
    .ZN(v27_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0029_ (
    .A1(n2),
    .A2(n11),
    .ZN(v28_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0030_ (
    .I(v28_0),
    .ZN(v29_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0031_ (
    .A1(v1_0),
    .A2(v29_0),
    .ZN(v30_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0032_ (
    .A1(v0_0),
    .A2(v28_0),
    .ZN(v31_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0033_ (
    .A1(v30_0),
    .A2(v31_0),
    .ZN(v32_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0034_ (
    .A1(n13),
    .A2(n0),
    .ZN(v33_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0035_ (
    .A1(v32_0),
    .A2(v33_0),
    .Z(v34_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0036_ (
    .A1(v32_0),
    .A2(v33_0),
    .ZN(v35_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0037_ (
    .A1(v34_0),
    .A2(v35_0),
    .ZN(v36_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0038_ (
    .I(v14_0),
    .ZN(v37_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0039_ (
    .A1(v18_0),
    .A2(v37_0),
    .ZN(v38_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0040_ (
    .A1(v38_0),
    .A2(v16_0),
    .Z(v39_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0041_ (
    .A1(n5),
    .A2(n8),
    .ZN(v40_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0042_ (
    .A1(v15_0),
    .A2(v40_0),
    .Z(v41_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0043_ (
    .A1(n10),
    .A2(n3),
    .ZN(v42_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0044_ (
    .I(v42_0),
    .ZN(v43_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0045_ (
    .A1(v41_0),
    .A2(v43_0),
    .ZN(v44_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0046_ (
    .A1(n5),
    .A2(n9),
    .ZN(v45_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0047_ (
    .A1(v17_0),
    .A2(v45_0),
    .Z(v46_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0048_ (
    .I(v41_0),
    .ZN(v47_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0049_ (
    .A1(v47_0),
    .A2(v42_0),
    .ZN(v48_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0050_ (
    .A1(v44_0),
    .A2(v48_0),
    .ZN(v49_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0051_ (
    .A1(v39_0),
    .A2(v49_0),
    .ZN(v50_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0052_ (
    .A1(v44_0),
    .A2(v48_0),
    .Z(v51_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0053_ (
    .A1(v38_0),
    .A2(v16_0),
    .ZN(v52_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0054_ (
    .A1(v51_0),
    .A2(v52_0),
    .ZN(v53_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0055_ (
    .A1(v50_0),
    .A2(v53_0),
    .ZN(v54_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0056_ (
    .A1(v36_0),
    .A2(v54_0),
    .Z(v55_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0057_ (
    .A1(v27_0),
    .A2(v55_0),
    .Z(v56_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0058_ (
    .A1(v5_0),
    .A2(v56_0),
    .Z(v57_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0059_ (
    .A1(v24_0),
    .A2(v21_0),
    .Z(v58_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0060_ (
    .I(n1),
    .ZN(v59_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0061_ (
    .A1(v7_0),
    .A2(v59_0),
    .Z(v60_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0062_ (
    .I(v60_0),
    .ZN(v61_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0063_ (
    .A1(v6_0),
    .A2(v61_0),
    .Z(v62_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0064_ (
    .A1(v62_0),
    .A2(v2_0),
    .Z(v63_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0065_ (
    .I(v61_0),
    .ZN(v64_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0066_ (
    .A1(v63_0),
    .A2(v64_0),
    .ZN(v65_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0067_ (
    .A1(v58_0),
    .A2(v65_0),
    .Z(v66_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0068_ (
    .A1(v2_0),
    .A2(v62_0),
    .Z(v67_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0069_ (
    .A1(v67_0),
    .A2(v24_0),
    .Z(v68_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0070_ (
    .A1(v66_0),
    .A2(v68_0),
    .ZN(v69_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0071_ (
    .A1(v65_0),
    .A2(v58_0),
    .ZN(v70_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0072_ (
    .A1(v69_0),
    .A2(v70_0),
    .ZN(v71_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0073_ (
    .A1(v57_0),
    .A2(v71_0),
    .Z(v72_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0074_ (
    .I(v24_0),
    .ZN(v73_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0075_ (
    .A1(v68_0),
    .A2(v66_0),
    .Z(v74_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0076_ (
    .I(v69_0),
    .ZN(v75_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0077_ (
    .A1(v75_0),
    .A2(v57_0),
    .Z(v76_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0078_ (
    .I(v70_0),
    .ZN(v77_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0079_ (
    .A1(v57_0),
    .A2(v77_0),
    .ZN(v78_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0080_ (
    .A1(v56_0),
    .A2(v5_0),
    .ZN(v79_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0081_ (
    .A1(v55_0),
    .A2(v27_0),
    .ZN(v80_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0082_ (
    .A1(v79_0),
    .A2(v80_0),
    .ZN(v81_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0083_ (
    .I(v81_0),
    .ZN(v82_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0084_ (
    .A1(v54_0),
    .A2(v36_0),
    .Z(v83_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0085_ (
    .A1(v83_0),
    .A2(v53_0),
    .ZN(v84_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0086_ (
    .A1(n3),
    .A2(n12),
    .ZN(v85_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0087_ (
    .I(v85_0),
    .ZN(v86_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0088_ (
    .A1(v86_0),
    .A2(v29_0),
    .ZN(v87_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0089_ (
    .A1(n2),
    .A2(n12),
    .ZN(v88_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0090_ (
    .A1(n3),
    .A2(n11),
    .ZN(v89_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0091_ (
    .A1(v88_0),
    .A2(v89_0),
    .ZN(v90_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0092_ (
    .A1(v87_0),
    .A2(v90_0),
    .ZN(v91_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0093_ (
    .A1(n1),
    .A2(n13),
    .ZN(v92_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0094_ (
    .A1(v91_0),
    .A2(v92_0),
    .Z(v93_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0095_ (
    .A1(v91_0),
    .A2(v92_0),
    .ZN(v94_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0096_ (
    .A1(v93_0),
    .A2(v94_0),
    .ZN(v95_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0097_ (
    .A1(v44_0),
    .A2(v46_0),
    .Z(v96_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0098_ (
    .A1(n8),
    .A2(n6),
    .ZN(v97_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0099_ (
    .A1(v45_0),
    .A2(v97_0),
    .ZN(v98_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0100_ (
    .A1(n4),
    .A2(n10),
    .ZN(v99_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0101_ (
    .I(v99_0),
    .ZN(v100_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0102_ (
    .A1(v98_0),
    .A2(v100_0),
    .ZN(v101_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0103_ (
    .A1(n5),
    .A2(n8),
    .Z(v102_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0104_ (
    .A1(n9),
    .A2(n6),
    .Z(v103_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0105_ (
    .A1(v102_0),
    .A2(v103_0),
    .ZN(v104_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0106_ (
    .A1(v104_0),
    .A2(v98_0),
    .ZN(v105_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0107_ (
    .A1(v105_0),
    .A2(v99_0),
    .ZN(v106_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0108_ (
    .A1(v101_0),
    .A2(v106_0),
    .ZN(v107_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0109_ (
    .A1(v96_0),
    .A2(v107_0),
    .ZN(v108_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0110_ (
    .A1(v99_0),
    .A2(v105_0),
    .Z(v109_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0111_ (
    .A1(v44_0),
    .A2(v46_0),
    .ZN(v110_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0112_ (
    .A1(v109_0),
    .A2(v110_0),
    .ZN(v111_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0113_ (
    .A1(v108_0),
    .A2(v111_0),
    .ZN(v112_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0114_ (
    .A1(v95_0),
    .A2(v112_0),
    .Z(v113_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0115_ (
    .A1(v84_0),
    .A2(v113_0),
    .Z(v114_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0116_ (
    .A1(n0),
    .A2(n14),
    .ZN(v115_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0117_ (
    .I(v115_0),
    .ZN(v116_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0118_ (
    .A1(v34_0),
    .A2(v30_0),
    .ZN(v117_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0119_ (
    .A1(v116_0),
    .A2(v117_0),
    .Z(v118_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0120_ (
    .A1(v114_0),
    .A2(v118_0),
    .ZN(v119_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0121_ (
    .A1(v113_0),
    .A2(v84_0),
    .ZN(v120_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0122_ (
    .I(v114_0),
    .ZN(v121_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0123_ (
    .I(v118_0),
    .ZN(v122_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0124_ (
    .A1(v121_0),
    .A2(v122_0),
    .ZN(v123_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0125_ (
    .A1(v119_0),
    .A2(v123_0),
    .ZN(v124_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0126_ (
    .A1(v82_0),
    .A2(v124_0),
    .ZN(v125_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0127_ (
    .I(v124_0),
    .ZN(v126_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0128_ (
    .A1(v126_0),
    .A2(v81_0),
    .ZN(v127_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0129_ (
    .A1(v125_0),
    .A2(v127_0),
    .ZN(v128_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0130_ (
    .A1(v78_0),
    .A2(v128_0),
    .Z(v129_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0131_ (
    .A1(v76_0),
    .A2(v129_0),
    .Z(v130_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0132_ (
    .A1(v129_0),
    .A2(v76_0),
    .ZN(v131_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0133_ (
    .A1(v128_0),
    .A2(v78_0),
    .Z(v132_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0134_ (
    .A1(v131_0),
    .A2(v132_0),
    .ZN(v133_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0135_ (
    .A1(v119_0),
    .A2(v120_0),
    .ZN(v134_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0136_ (
    .A1(v93_0),
    .A2(v87_0),
    .ZN(v135_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0137_ (
    .A1(n1),
    .A2(n14),
    .ZN(v136_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0138_ (
    .A1(n2),
    .A2(n13),
    .ZN(v137_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0139_ (
    .A1(v136_0),
    .A2(v137_0),
    .Z(v138_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0140_ (
    .I(v138_0),
    .ZN(v139_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0141_ (
    .I(n15),
    .ZN(v140_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0142_ (
    .A1(v140_0),
    .A2(n0),
    .Z(v141_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0143_ (
    .A1(v139_0),
    .A2(v141_0),
    .Z(v142_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0144_ (
    .A1(v139_0),
    .A2(v141_0),
    .ZN(v143_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0145_ (
    .A1(v142_0),
    .A2(v143_0),
    .ZN(v144_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0146_ (
    .A1(v135_0),
    .A2(v144_0),
    .Z(v145_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0147_ (
    .I(v95_0),
    .ZN(v146_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0148_ (
    .A1(v108_0),
    .A2(v146_0),
    .ZN(v147_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0149_ (
    .A1(v147_0),
    .A2(v111_0),
    .Z(v148_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0150_ (
    .A1(n8),
    .A2(n7),
    .ZN(v149_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0151_ (
    .A1(v140_0),
    .A2(v149_0),
    .Z(v150_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0152_ (
    .A1(v150_0),
    .A2(v103_0),
    .ZN(v151_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0153_ (
    .A1(n8),
    .A2(n7),
    .Z(v152_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0154_ (
    .A1(v152_0),
    .A2(n15),
    .ZN(v153_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0155_ (
    .I(v150_0),
    .ZN(v154_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0156_ (
    .I(v103_0),
    .ZN(v155_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0157_ (
    .A1(v154_0),
    .A2(v155_0),
    .ZN(v156_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0158_ (
    .A1(v151_0),
    .A2(v156_0),
    .ZN(v157_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0159_ (
    .A1(v101_0),
    .A2(v104_0),
    .ZN(v158_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0160_ (
    .A1(v157_0),
    .A2(v158_0),
    .Z(v159_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0161_ (
    .A1(n5),
    .A2(n11),
    .ZN(v160_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0162_ (
    .A1(v99_0),
    .A2(v160_0),
    .Z(v161_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0163_ (
    .A1(n4),
    .A2(n11),
    .ZN(v162_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0164_ (
    .A1(n5),
    .A2(n10),
    .ZN(v163_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0165_ (
    .A1(v162_0),
    .A2(v163_0),
    .ZN(v164_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0166_ (
    .A1(v161_0),
    .A2(v164_0),
    .ZN(v165_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0167_ (
    .A1(v165_0),
    .A2(v85_0),
    .Z(v166_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0168_ (
    .A1(v165_0),
    .A2(v85_0),
    .ZN(v167_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0169_ (
    .A1(v166_0),
    .A2(v167_0),
    .ZN(v168_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0170_ (
    .A1(v159_0),
    .A2(v168_0),
    .Z(v169_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0171_ (
    .A1(v159_0),
    .A2(v168_0),
    .ZN(v170_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0172_ (
    .A1(v169_0),
    .A2(v170_0),
    .ZN(v171_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0173_ (
    .A1(v148_0),
    .A2(v171_0),
    .ZN(v172_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0174_ (
    .A1(v168_0),
    .A2(v159_0),
    .Z(v173_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0175_ (
    .A1(v147_0),
    .A2(v111_0),
    .ZN(v174_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0176_ (
    .A1(v173_0),
    .A2(v174_0),
    .ZN(v175_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0177_ (
    .A1(v172_0),
    .A2(v175_0),
    .ZN(v176_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0178_ (
    .A1(v145_0),
    .A2(v176_0),
    .Z(v177_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0179_ (
    .A1(v134_0),
    .A2(v177_0),
    .Z(v178_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0180_ (
    .A1(v117_0),
    .A2(v122_0),
    .ZN(v179_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0181_ (
    .I(v179_0),
    .ZN(v180_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0182_ (
    .A1(v178_0),
    .A2(v180_0),
    .ZN(v181_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0183_ (
    .A1(v177_0),
    .A2(v134_0),
    .ZN(v182_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0184_ (
    .I(v178_0),
    .ZN(v183_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0185_ (
    .A1(v183_0),
    .A2(v179_0),
    .ZN(v184_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0186_ (
    .A1(v181_0),
    .A2(v184_0),
    .ZN(v185_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0187_ (
    .A1(v127_0),
    .A2(v185_0),
    .Z(v186_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0188_ (
    .A1(v133_0),
    .A2(v186_0),
    .Z(v187_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0189_ (
    .A1(v181_0),
    .A2(v182_0),
    .ZN(v188_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0190_ (
    .A1(v145_0),
    .A2(v135_0),
    .ZN(v189_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0191_ (
    .A1(v176_0),
    .A2(v145_0),
    .Z(v190_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0192_ (
    .A1(v190_0),
    .A2(v175_0),
    .ZN(v191_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0193_ (
    .A1(n5),
    .A2(n12),
    .ZN(v192_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0194_ (
    .A1(v162_0),
    .A2(v192_0),
    .Z(v193_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0195_ (
    .A1(n4),
    .A2(n12),
    .ZN(v194_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0196_ (
    .A1(v160_0),
    .A2(v194_0),
    .ZN(v195_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0197_ (
    .A1(v193_0),
    .A2(v195_0),
    .ZN(v196_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0198_ (
    .A1(n3),
    .A2(n13),
    .ZN(v197_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0199_ (
    .A1(v196_0),
    .A2(v197_0),
    .Z(v198_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0200_ (
    .A1(v196_0),
    .A2(v197_0),
    .ZN(v199_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0201_ (
    .A1(v198_0),
    .A2(v199_0),
    .ZN(v200_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0202_ (
    .A1(v151_0),
    .A2(v153_0),
    .ZN(v201_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0203_ (
    .A1(v152_0),
    .A2(n9),
    .ZN(v202_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0204_ (
    .A1(n9),
    .A2(n7),
    .ZN(v203_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0205_ (
    .A1(v149_0),
    .A2(v203_0),
    .ZN(v204_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0206_ (
    .A1(v202_0),
    .A2(v204_0),
    .ZN(v205_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0207_ (
    .A1(n10),
    .A2(n6),
    .ZN(v206_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0208_ (
    .A1(v205_0),
    .A2(v206_0),
    .Z(v207_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0209_ (
    .A1(v205_0),
    .A2(v206_0),
    .ZN(v208_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0210_ (
    .A1(v207_0),
    .A2(v208_0),
    .ZN(v209_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0211_ (
    .A1(v201_0),
    .A2(v209_0),
    .Z(v210_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0212_ (
    .A1(v200_0),
    .A2(v210_0),
    .Z(v211_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0213_ (
    .A1(v159_0),
    .A2(v158_0),
    .ZN(v212_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0214_ (
    .A1(v169_0),
    .A2(v212_0),
    .ZN(v213_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0215_ (
    .A1(v211_0),
    .A2(v213_0),
    .Z(v214_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0216_ (
    .A1(v211_0),
    .A2(v213_0),
    .ZN(v215_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0217_ (
    .A1(v214_0),
    .A2(v215_0),
    .ZN(v216_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0218_ (
    .A1(n2),
    .A2(n14),
    .ZN(v217_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0219_ (
    .A1(v92_0),
    .A2(v217_0),
    .Z(v218_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0220_ (
    .A1(v142_0),
    .A2(v218_0),
    .ZN(v219_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0221_ (
    .A1(v166_0),
    .A2(v161_0),
    .ZN(v220_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0222_ (
    .A1(v59_0),
    .A2(n15),
    .ZN(v221_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0223_ (
    .A1(v217_0),
    .A2(v221_0),
    .Z(v222_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0224_ (
    .A1(v220_0),
    .A2(v222_0),
    .Z(v223_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0225_ (
    .A1(v220_0),
    .A2(v222_0),
    .ZN(v224_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0226_ (
    .A1(v223_0),
    .A2(v224_0),
    .ZN(v225_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0227_ (
    .A1(v219_0),
    .A2(v225_0),
    .Z(v226_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0228_ (
    .A1(v216_0),
    .A2(v226_0),
    .Z(v227_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0229_ (
    .A1(v216_0),
    .A2(v226_0),
    .ZN(v228_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0230_ (
    .A1(v227_0),
    .A2(v228_0),
    .ZN(v229_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0231_ (
    .A1(v191_0),
    .A2(v229_0),
    .Z(v230_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0232_ (
    .A1(v189_0),
    .A2(v230_0),
    .Z(v231_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0233_ (
    .A1(v188_0),
    .A2(v231_0),
    .Z(v232_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0234_ (
    .A1(v186_0),
    .A2(v133_0),
    .ZN(v233_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0235_ (
    .A1(v185_0),
    .A2(v127_0),
    .Z(v234_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0236_ (
    .A1(v233_0),
    .A2(v234_0),
    .ZN(v235_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0237_ (
    .A1(v232_0),
    .A2(v235_0),
    .Z(v236_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0238_ (
    .A1(v226_0),
    .A2(v219_0),
    .ZN(v237_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0239_ (
    .A1(v237_0),
    .A2(v224_0),
    .ZN(v238_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0240_ (
    .I(v238_0),
    .ZN(v239_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0241_ (
    .A1(v227_0),
    .A2(v215_0),
    .ZN(v240_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0242_ (
    .A1(v210_0),
    .A2(v200_0),
    .Z(v241_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0243_ (
    .A1(v210_0),
    .A2(v201_0),
    .ZN(v242_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0244_ (
    .A1(v241_0),
    .A2(v242_0),
    .ZN(v243_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0245_ (
    .A1(n11),
    .A2(n6),
    .ZN(v244_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0246_ (
    .A1(v192_0),
    .A2(v244_0),
    .Z(v245_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0247_ (
    .I(v245_0),
    .ZN(v246_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0248_ (
    .A1(n4),
    .A2(n13),
    .ZN(v247_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0249_ (
    .A1(v246_0),
    .A2(v247_0),
    .Z(v248_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0250_ (
    .A1(v246_0),
    .A2(v247_0),
    .ZN(v249_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0251_ (
    .A1(v248_0),
    .A2(v249_0),
    .ZN(v250_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0252_ (
    .A1(n10),
    .A2(n7),
    .ZN(v251_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0253_ (
    .A1(v251_0),
    .A2(v205_0),
    .Z(v252_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0254_ (
    .A1(v207_0),
    .A2(v202_0),
    .ZN(v253_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0255_ (
    .A1(v252_0),
    .A2(v253_0),
    .Z(v254_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0256_ (
    .A1(v252_0),
    .A2(v253_0),
    .ZN(v255_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0257_ (
    .A1(v254_0),
    .A2(v255_0),
    .Z(v256_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0258_ (
    .A1(v250_0),
    .A2(v256_0),
    .Z(v257_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0259_ (
    .A1(v243_0),
    .A2(v257_0),
    .Z(v258_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0260_ (
    .A1(v221_0),
    .A2(v217_0),
    .Z(v259_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0261_ (
    .A1(n3),
    .A2(n14),
    .ZN(v260_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0262_ (
    .I(n2),
    .ZN(v261_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0263_ (
    .A1(v261_0),
    .A2(n15),
    .ZN(v262_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0264_ (
    .A1(v260_0),
    .A2(v262_0),
    .Z(v263_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0265_ (
    .A1(v198_0),
    .A2(v193_0),
    .ZN(v264_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0266_ (
    .A1(v263_0),
    .A2(v264_0),
    .Z(v265_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0267_ (
    .I(v265_0),
    .ZN(v266_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0268_ (
    .A1(v259_0),
    .A2(v266_0),
    .Z(v267_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0269_ (
    .I(v267_0),
    .ZN(v268_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0270_ (
    .A1(v258_0),
    .A2(v268_0),
    .Z(v269_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0271_ (
    .A1(v258_0),
    .A2(v268_0),
    .ZN(v270_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0272_ (
    .A1(v269_0),
    .A2(v270_0),
    .ZN(v271_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0273_ (
    .A1(v240_0),
    .A2(v271_0),
    .Z(v272_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0274_ (
    .A1(v239_0),
    .A2(v272_0),
    .Z(v273_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0275_ (
    .A1(v230_0),
    .A2(v189_0),
    .Z(v274_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0276_ (
    .A1(v230_0),
    .A2(v191_0),
    .ZN(v275_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0277_ (
    .A1(v274_0),
    .A2(v275_0),
    .ZN(v276_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0278_ (
    .A1(v273_0),
    .A2(v276_0),
    .Z(v277_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0279_ (
    .A1(v273_0),
    .A2(v276_0),
    .ZN(v278_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0280_ (
    .A1(v277_0),
    .A2(v278_0),
    .Z(v279_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0281_ (
    .A1(v235_0),
    .A2(v232_0),
    .Z(v280_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0282_ (
    .I(v280_0),
    .ZN(v281_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0283_ (
    .A1(v231_0),
    .A2(v188_0),
    .ZN(v282_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0284_ (
    .A1(v281_0),
    .A2(v282_0),
    .ZN(v283_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0285_ (
    .A1(v279_0),
    .A2(v283_0),
    .Z(v284_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0286_ (
    .A1(v272_0),
    .A2(v239_0),
    .Z(v285_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0287_ (
    .A1(v272_0),
    .A2(v240_0),
    .ZN(v286_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0288_ (
    .A1(v285_0),
    .A2(v286_0),
    .ZN(v287_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0289_ (
    .A1(v266_0),
    .A2(v259_0),
    .Z(v288_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0290_ (
    .A1(v264_0),
    .A2(v263_0),
    .ZN(v289_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0291_ (
    .A1(v288_0),
    .A2(v289_0),
    .ZN(v290_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0292_ (
    .A1(n4),
    .A2(n14),
    .ZN(v291_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0293_ (
    .I(n3),
    .ZN(v292_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0294_ (
    .A1(v292_0),
    .A2(n15),
    .ZN(v293_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0295_ (
    .A1(v291_0),
    .A2(v293_0),
    .Z(v294_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0296_ (
    .A1(n12),
    .A2(n6),
    .ZN(v295_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0297_ (
    .A1(v160_0),
    .A2(v295_0),
    .Z(v296_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0298_ (
    .A1(v248_0),
    .A2(v296_0),
    .ZN(v297_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0299_ (
    .A1(v294_0),
    .A2(v297_0),
    .Z(v298_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0300_ (
    .I(v298_0),
    .ZN(v299_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0301_ (
    .A1(v262_0),
    .A2(v260_0),
    .Z(v300_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0302_ (
    .A1(v299_0),
    .A2(v300_0),
    .Z(v301_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0303_ (
    .A1(v299_0),
    .A2(v300_0),
    .ZN(v302_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0304_ (
    .A1(v301_0),
    .A2(v302_0),
    .ZN(v303_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0305_ (
    .A1(v256_0),
    .A2(v257_0),
    .ZN(v304_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0306_ (
    .A1(v304_0),
    .A2(v255_0),
    .ZN(v305_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0307_ (
    .I(v204_0),
    .ZN(v306_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0308_ (
    .A1(v306_0),
    .A2(v251_0),
    .ZN(v307_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0309_ (
    .A1(v255_0),
    .A2(v307_0),
    .ZN(v308_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0310_ (
    .A1(n11),
    .A2(n7),
    .ZN(v309_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0311_ (
    .A1(v295_0),
    .A2(v309_0),
    .Z(v310_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0312_ (
    .I(v310_0),
    .ZN(v311_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0313_ (
    .A1(n5),
    .A2(n13),
    .ZN(v312_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0314_ (
    .A1(v311_0),
    .A2(v312_0),
    .Z(v313_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0315_ (
    .A1(v311_0),
    .A2(v312_0),
    .ZN(v314_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0316_ (
    .A1(v313_0),
    .A2(v314_0),
    .Z(v315_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0317_ (
    .I(v315_0),
    .ZN(v316_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0318_ (
    .A1(v308_0),
    .A2(v316_0),
    .Z(v317_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0319_ (
    .A1(v305_0),
    .A2(v317_0),
    .Z(v318_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0320_ (
    .A1(v305_0),
    .A2(v317_0),
    .ZN(v319_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0321_ (
    .A1(v318_0),
    .A2(v319_0),
    .ZN(v320_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0322_ (
    .A1(v303_0),
    .A2(v320_0),
    .Z(v321_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0323_ (
    .A1(v258_0),
    .A2(v243_0),
    .ZN(v322_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0324_ (
    .A1(v269_0),
    .A2(v322_0),
    .ZN(v323_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0325_ (
    .A1(v321_0),
    .A2(v323_0),
    .Z(v324_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0326_ (
    .A1(v290_0),
    .A2(v324_0),
    .Z(v325_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0327_ (
    .A1(v287_0),
    .A2(v325_0),
    .Z(v326_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0328_ (
    .A1(v280_0),
    .A2(v279_0),
    .ZN(v327_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0329_ (
    .A1(v278_0),
    .A2(v282_0),
    .ZN(v328_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0330_ (
    .A1(v328_0),
    .A2(v277_0),
    .ZN(v329_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0331_ (
    .A1(v327_0),
    .A2(v329_0),
    .ZN(v330_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0332_ (
    .A1(v326_0),
    .A2(v330_0),
    .Z(v331_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0333_ (
    .A1(v297_0),
    .A2(v294_0),
    .ZN(v332_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0334_ (
    .A1(v301_0),
    .A2(v332_0),
    .ZN(v333_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0335_ (
    .A1(v320_0),
    .A2(v303_0),
    .Z(v334_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0336_ (
    .A1(v334_0),
    .A2(v319_0),
    .ZN(v335_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0337_ (
    .A1(n5),
    .A2(n14),
    .ZN(v336_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0338_ (
    .I(n4),
    .ZN(v337_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0339_ (
    .A1(v337_0),
    .A2(n15),
    .ZN(v338_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0340_ (
    .A1(v336_0),
    .A2(v338_0),
    .Z(v339_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0341_ (
    .A1(v295_0),
    .A2(v309_0),
    .Z(v340_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0342_ (
    .A1(v313_0),
    .A2(v340_0),
    .ZN(v341_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0343_ (
    .A1(v339_0),
    .A2(v341_0),
    .Z(v342_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0344_ (
    .I(v342_0),
    .ZN(v343_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0345_ (
    .A1(v293_0),
    .A2(v291_0),
    .Z(v344_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0346_ (
    .A1(v343_0),
    .A2(v344_0),
    .Z(v345_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0347_ (
    .A1(v343_0),
    .A2(v344_0),
    .ZN(v346_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0348_ (
    .A1(v345_0),
    .A2(v346_0),
    .Z(v347_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0349_ (
    .I(v308_0),
    .ZN(v348_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0350_ (
    .A1(v348_0),
    .A2(v315_0),
    .ZN(v349_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0351_ (
    .A1(v349_0),
    .A2(v255_0),
    .ZN(v350_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0352_ (
    .I(v309_0),
    .ZN(v351_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0353_ (
    .A1(v351_0),
    .A2(n12),
    .ZN(v352_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0354_ (
    .A1(n12),
    .A2(n7),
    .ZN(v353_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0355_ (
    .A1(v309_0),
    .A2(v353_0),
    .ZN(v354_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0356_ (
    .A1(v352_0),
    .A2(v354_0),
    .ZN(v355_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0357_ (
    .A1(n13),
    .A2(n6),
    .ZN(v356_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0358_ (
    .A1(v355_0),
    .A2(v356_0),
    .Z(v357_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0359_ (
    .A1(v355_0),
    .A2(v356_0),
    .ZN(v358_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0360_ (
    .A1(v357_0),
    .A2(v358_0),
    .Z(v359_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0361_ (
    .I(v359_0),
    .ZN(v360_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0362_ (
    .A1(v360_0),
    .A2(v308_0),
    .Z(v361_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0363_ (
    .A1(v350_0),
    .A2(v361_0),
    .Z(v362_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0364_ (
    .A1(v350_0),
    .A2(v361_0),
    .ZN(v363_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0365_ (
    .A1(v362_0),
    .A2(v363_0),
    .Z(v364_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0366_ (
    .A1(v347_0),
    .A2(v364_0),
    .Z(v365_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0367_ (
    .A1(v335_0),
    .A2(v365_0),
    .Z(v366_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0368_ (
    .A1(v333_0),
    .A2(v366_0),
    .Z(v367_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0369_ (
    .A1(v324_0),
    .A2(v290_0),
    .ZN(v368_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0370_ (
    .A1(v323_0),
    .A2(v321_0),
    .ZN(v369_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0371_ (
    .A1(v368_0),
    .A2(v369_0),
    .ZN(v370_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0372_ (
    .A1(v367_0),
    .A2(v370_0),
    .Z(v371_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0373_ (
    .A1(v367_0),
    .A2(v370_0),
    .ZN(v372_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0374_ (
    .A1(v371_0),
    .A2(v372_0),
    .Z(v373_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0375_ (
    .A1(v330_0),
    .A2(v326_0),
    .ZN(v374_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0376_ (
    .A1(v325_0),
    .A2(v287_0),
    .ZN(v375_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0377_ (
    .A1(v374_0),
    .A2(v375_0),
    .ZN(v376_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0378_ (
    .A1(v373_0),
    .A2(v376_0),
    .Z(v377_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0379_ (
    .A1(v366_0),
    .A2(v333_0),
    .ZN(v378_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0380_ (
    .A1(v365_0),
    .A2(v335_0),
    .ZN(v379_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0381_ (
    .A1(v378_0),
    .A2(v379_0),
    .ZN(v380_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0382_ (
    .A1(v341_0),
    .A2(v339_0),
    .ZN(v381_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0383_ (
    .A1(v345_0),
    .A2(v381_0),
    .ZN(v382_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0384_ (
    .A1(v364_0),
    .A2(v347_0),
    .ZN(v383_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0385_ (
    .A1(v383_0),
    .A2(v363_0),
    .ZN(v384_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0386_ (
    .A1(n6),
    .A2(n14),
    .ZN(v385_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0387_ (
    .I(n5),
    .ZN(v386_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0388_ (
    .A1(v386_0),
    .A2(n15),
    .ZN(v387_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0389_ (
    .A1(v385_0),
    .A2(v387_0),
    .Z(v388_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0390_ (
    .A1(v357_0),
    .A2(v352_0),
    .ZN(v389_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0391_ (
    .A1(v388_0),
    .A2(v389_0),
    .Z(v390_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0392_ (
    .I(v390_0),
    .ZN(v391_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0393_ (
    .A1(v338_0),
    .A2(v336_0),
    .Z(v392_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0394_ (
    .A1(v391_0),
    .A2(v392_0),
    .Z(v393_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0395_ (
    .A1(v391_0),
    .A2(v392_0),
    .ZN(v394_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0396_ (
    .A1(v393_0),
    .A2(v394_0),
    .Z(v395_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0397_ (
    .A1(v307_0),
    .A2(v359_0),
    .ZN(v396_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0398_ (
    .A1(v396_0),
    .A2(v255_0),
    .ZN(v397_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0399_ (
    .A1(n13),
    .A2(n7),
    .ZN(v398_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0400_ (
    .A1(v398_0),
    .A2(v355_0),
    .Z(v399_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0401_ (
    .I(v399_0),
    .ZN(v400_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0402_ (
    .A1(v400_0),
    .A2(v308_0),
    .Z(v401_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0403_ (
    .A1(v397_0),
    .A2(v401_0),
    .Z(v402_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0404_ (
    .A1(v397_0),
    .A2(v401_0),
    .ZN(v403_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0405_ (
    .A1(v402_0),
    .A2(v403_0),
    .Z(v404_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0406_ (
    .A1(v395_0),
    .A2(v404_0),
    .Z(v405_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0407_ (
    .A1(v384_0),
    .A2(v405_0),
    .Z(v406_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0408_ (
    .A1(v382_0),
    .A2(v406_0),
    .Z(v407_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0409_ (
    .A1(v380_0),
    .A2(v407_0),
    .Z(v408_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0410_ (
    .A1(v375_0),
    .A2(v373_0),
    .Z(v409_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0411_ (
    .A1(v374_0),
    .A2(v409_0),
    .ZN(v410_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0412_ (
    .A1(v410_0),
    .A2(v371_0),
    .Z(v411_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0413_ (
    .A1(v408_0),
    .A2(v411_0),
    .Z(v412_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0414_ (
    .A1(v389_0),
    .A2(v388_0),
    .ZN(v413_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0415_ (
    .A1(v393_0),
    .A2(v413_0),
    .ZN(v414_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0416_ (
    .A1(v404_0),
    .A2(v395_0),
    .ZN(v415_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0417_ (
    .A1(v415_0),
    .A2(v403_0),
    .ZN(v416_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0418_ (
    .A1(v308_0),
    .A2(v400_0),
    .Z(v417_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0419_ (
    .A1(v417_0),
    .A2(v255_0),
    .ZN(v418_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0420_ (
    .A1(v400_0),
    .A2(v255_0),
    .Z(v419_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0421_ (
    .A1(v418_0),
    .A2(v419_0),
    .ZN(v420_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0422_ (
    .I(v420_0),
    .ZN(v421_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0423_ (
    .A1(v355_0),
    .A2(v398_0),
    .Z(v422_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0424_ (
    .A1(v422_0),
    .A2(v352_0),
    .ZN(v423_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0425_ (
    .I(v423_0),
    .ZN(v424_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0426_ (
    .A1(n14),
    .A2(n7),
    .ZN(v425_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0427_ (
    .I(v425_0),
    .ZN(v426_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0428_ (
    .A1(v140_0),
    .A2(n6),
    .Z(v427_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0429_ (
    .A1(v426_0),
    .A2(v427_0),
    .Z(v428_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0430_ (
    .A1(v424_0),
    .A2(v428_0),
    .Z(v429_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0431_ (
    .A1(v424_0),
    .A2(v428_0),
    .ZN(v430_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0432_ (
    .A1(v429_0),
    .A2(v430_0),
    .Z(v431_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0433_ (
    .I(v431_0),
    .ZN(v432_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0434_ (
    .A1(v387_0),
    .A2(v385_0),
    .Z(v433_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0435_ (
    .A1(v432_0),
    .A2(v433_0),
    .Z(v434_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0436_ (
    .A1(v432_0),
    .A2(v433_0),
    .ZN(v435_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0437_ (
    .A1(v434_0),
    .A2(v435_0),
    .Z(v436_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0438_ (
    .A1(v421_0),
    .A2(v436_0),
    .Z(v437_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0439_ (
    .A1(v416_0),
    .A2(v437_0),
    .Z(v438_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0440_ (
    .A1(v414_0),
    .A2(v438_0),
    .Z(v439_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0441_ (
    .A1(v406_0),
    .A2(v382_0),
    .ZN(v440_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0442_ (
    .A1(v405_0),
    .A2(v384_0),
    .ZN(v441_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0443_ (
    .A1(v440_0),
    .A2(v441_0),
    .ZN(v442_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0444_ (
    .A1(v439_0),
    .A2(v442_0),
    .Z(v443_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0445_ (
    .A1(v439_0),
    .A2(v442_0),
    .ZN(v444_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0446_ (
    .A1(v443_0),
    .A2(v444_0),
    .Z(v445_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0447_ (
    .A1(v411_0),
    .A2(v408_0),
    .ZN(v446_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0448_ (
    .A1(v407_0),
    .A2(v380_0),
    .ZN(v447_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0449_ (
    .A1(v446_0),
    .A2(v447_0),
    .ZN(v448_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0450_ (
    .A1(v445_0),
    .A2(v448_0),
    .Z(v449_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0451_ (
    .A1(v434_0),
    .A2(v429_0),
    .ZN(v450_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0452_ (
    .A1(v427_0),
    .A2(v426_0),
    .ZN(v451_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0453_ (
    .A1(v140_0),
    .A2(n7),
    .Z(v452_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0454_ (
    .A1(v451_0),
    .A2(v452_0),
    .ZN(v453_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0455_ (
    .A1(v453_0),
    .A2(v423_0),
    .Z(v454_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0456_ (
    .A1(v454_0),
    .A2(v421_0),
    .Z(v455_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0457_ (
    .A1(v436_0),
    .A2(v421_0),
    .ZN(v456_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0458_ (
    .A1(v456_0),
    .A2(v419_0),
    .ZN(v457_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0459_ (
    .A1(v455_0),
    .A2(v457_0),
    .Z(v458_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0460_ (
    .A1(v450_0),
    .A2(v458_0),
    .Z(v459_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0461_ (
    .A1(v438_0),
    .A2(v414_0),
    .ZN(v460_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0462_ (
    .A1(v437_0),
    .A2(v416_0),
    .ZN(v461_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0463_ (
    .A1(v460_0),
    .A2(v461_0),
    .ZN(v462_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0464_ (
    .A1(v459_0),
    .A2(v462_0),
    .Z(v463_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0465_ (
    .A1(v448_0),
    .A2(v443_0),
    .ZN(v464_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0466_ (
    .A1(v464_0),
    .A2(v444_0),
    .ZN(v465_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0467_ (
    .A1(v463_0),
    .A2(v465_0),
    .Z(v466_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0468_ (
    .I(v463_0),
    .ZN(v467_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0469_ (
    .A1(v467_0),
    .A2(v436_0),
    .ZN(v468_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0470_ (
    .A1(v466_0),
    .A2(v468_0),
    .Z(v469_0)
  );

  assign OUT[0] = v358_0;
  assign OUT[1] = v6_0;
  assign OUT[2] = n10;
  assign OUT[3] = v73_0;
  assign OUT[4] = v74_0;
  assign OUT[5] = v72_0;
  assign OUT[6] = v130_0;
  assign OUT[7] = v187_0;
  assign OUT[8] = v236_0;
  assign OUT[9] = v284_0;
  assign OUT[10] = v331_0;
  assign OUT[11] = v377_0;
  assign OUT[12] = v412_0;
  assign OUT[13] = v449_0;
  assign OUT[14] = v466_0;
  assign OUT[15] = v469_0;
endmodule
