* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_nfet_latch__tox_slope=5.989e-03
.param sky130_fd_pr__special_nfet_latch__vth0_slope=5.289e-03
.param sky130_fd_pr__special_nfet_latch__lint_slope=0
.param sky130_fd_pr__special_nfet_latch__wint_slope=0
.param sky130_fd_pr__special_nfet_latch__nfactor_slope=0.0
.param sky130_fd_pr__special_nfet_latch__voff_slope=0.00
