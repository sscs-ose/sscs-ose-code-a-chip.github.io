* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff = -0.0535
* Number of bins: 9
.param
+ sky130_fd_pr__nfet_03v3_nvt__toxe_mult = 1.0
+ sky130_fd_pr__nfet_03v3_nvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_03v3_nvt__overlap_mult = 0.77117
+ sky130_fd_pr__nfet_03v3_nvt__ajunction_mult = 0.97602
+ sky130_fd_pr__nfet_03v3_nvt__pjunction_mult = 1.0437
+ sky130_fd_pr__nfet_03v3_nvt__lint_diff = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__wint_diff = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__dlc_diff = -1.5781e-8
+ sky130_fd_pr__nfet_03v3_nvt__dwc_diff = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_0 = 0.038449
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_0 = 0.0019135
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0 = -1.3838
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0 = ' -0.015836 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_0 = -0.00065697
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0 = -3837.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_0 = -1.4132e-19
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_0 = 3.4977e-11
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_1 = 5.3407e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_1 = 0.033082
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_1 = 0.0096743
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1 = -1.3958
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1 = ' -0.015324 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_1 = -0.0011594
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1 = -6763.8
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_1 = 1.0429e-19
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_2 = 2.6095e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_2 = 5.8204e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_2 = 0.0057767
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2 = -0.46503
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2 = ' 0.0032323 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_2 = 0.0063254
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2 = -4056.8
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_2 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_3 = -3.3361e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_3 = 3.7397e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_3 = 0.040673
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_3 = 0.0032721
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3 = -1.3621
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3 = ' -0.01875 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_3 = -0.00011074
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3 = -4396.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_3 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_4 = 3.7224e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_4 = 2.2268e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_4 = 0.045453
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_4 = 0.010004
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4 = -1.3404
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4 = ' -0.018338 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_4 = -0.0018856
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4 = -8376.1
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_5 = 0.011241
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5 = -6843.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_5 = 3.0597e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_5 = 7.2969e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_5 = 0.012715
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5 = -1.6434
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5 = ' 0.051876 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6 = -0.746
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6 = ' 0.022008 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_6 = 0.007881
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6 = -3534.9
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_6 = 2.3973e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_6 = 8.5737e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_6 = 0.012066
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_7 = 0.04193
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_7 = 0.011117
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7 = -1.3436
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7 = ' -0.014154 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_7 = -0.0017689
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7 = -7893.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_7 = 2.6547e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_7 = 4.0061e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_7 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_8 = 0.0084797
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8 = -0.43724
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8 = ' -0.0034771 + sky130_fd_pr__nfet_03v3_nvt__vth0_correldiff'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_8 = 0.005952
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8 = -5528.9
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_8 = 2.4645e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_8 = 5.5525e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8 = 0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"
