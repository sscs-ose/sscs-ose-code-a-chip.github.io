# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.010000 BY  4.900000 ;
  PIN BULK
    ANTENNADIFFAREA  3.913000 ;
    ANTENNAGATEAREA  0.903000 ;
    PORT
      LAYER li1 ;
        RECT 0.205000 0.925000 0.800000 3.975000 ;
        RECT 0.600000 0.455000 0.930000 0.785000 ;
        RECT 0.600000 0.785000 0.800000 0.925000 ;
        RECT 0.600000 3.975000 0.800000 4.115000 ;
        RECT 0.600000 4.115000 0.930000 4.445000 ;
        RECT 3.080000 0.455000 3.410000 0.785000 ;
        RECT 3.080000 4.115000 3.410000 4.445000 ;
        RECT 3.210000 0.785000 3.410000 0.925000 ;
        RECT 3.210000 0.925000 3.805000 3.975000 ;
        RECT 3.210000 3.975000 3.410000 4.115000 ;
      LAYER mcon ;
        RECT 0.300000 1.105000 0.470000 1.275000 ;
        RECT 0.300000 1.465000 0.470000 1.635000 ;
        RECT 0.300000 1.825000 0.470000 1.995000 ;
        RECT 0.300000 2.185000 0.470000 2.355000 ;
        RECT 0.300000 2.545000 0.470000 2.715000 ;
        RECT 0.300000 2.905000 0.470000 3.075000 ;
        RECT 0.300000 3.265000 0.470000 3.435000 ;
        RECT 0.300000 3.625000 0.470000 3.795000 ;
        RECT 3.540000 1.105000 3.710000 1.275000 ;
        RECT 3.540000 1.465000 3.710000 1.635000 ;
        RECT 3.540000 1.825000 3.710000 1.995000 ;
        RECT 3.540000 2.185000 3.710000 2.355000 ;
        RECT 3.540000 2.545000 3.710000 2.715000 ;
        RECT 3.540000 2.905000 3.710000 3.075000 ;
        RECT 3.540000 3.265000 3.710000 3.435000 ;
        RECT 3.540000 3.625000 3.710000 3.795000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.205000 1.045000 0.500000 3.855000 ;
        RECT 3.510000 1.045000 3.805000 3.855000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.575000 3.940000 3.855000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.806000 ;
    PORT
      LAYER li1 ;
        RECT 1.215000 0.000000 2.795000 0.695000 ;
        RECT 1.215000 4.205000 2.795000 4.900000 ;
      LAYER mcon ;
        RECT 1.275000 0.095000 1.445000 0.265000 ;
        RECT 1.275000 0.455000 1.445000 0.625000 ;
        RECT 1.275000 4.275000 1.445000 4.445000 ;
        RECT 1.275000 4.635000 1.445000 4.805000 ;
        RECT 1.685000 0.095000 1.855000 0.265000 ;
        RECT 1.685000 0.455000 1.855000 0.625000 ;
        RECT 1.685000 4.275000 1.855000 4.445000 ;
        RECT 1.685000 4.635000 1.855000 4.805000 ;
        RECT 2.155000 0.095000 2.325000 0.265000 ;
        RECT 2.155000 0.455000 2.325000 0.625000 ;
        RECT 2.155000 4.275000 2.325000 4.445000 ;
        RECT 2.155000 4.635000 2.325000 4.805000 ;
        RECT 2.565000 0.095000 2.735000 0.265000 ;
        RECT 2.565000 0.455000 2.735000 0.625000 ;
        RECT 2.565000 4.275000 2.735000 4.445000 ;
        RECT 2.565000 4.635000 2.735000 4.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.215000 0.000000 2.795000 0.685000 ;
        RECT 1.215000 4.215000 2.795000 4.900000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.528400 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.045000 3.940000 2.325000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 1.060000 0.925000 1.230000 3.975000 ;
      RECT 1.490000 0.925000 1.660000 3.975000 ;
      RECT 1.920000 0.925000 2.090000 3.975000 ;
      RECT 2.350000 0.925000 2.520000 3.975000 ;
      RECT 2.780000 0.925000 2.950000 3.975000 ;
    LAYER mcon ;
      RECT 1.060000 1.105000 1.230000 1.275000 ;
      RECT 1.060000 1.465000 1.230000 1.635000 ;
      RECT 1.060000 1.825000 1.230000 1.995000 ;
      RECT 1.060000 2.185000 1.230000 2.355000 ;
      RECT 1.060000 2.545000 1.230000 2.715000 ;
      RECT 1.060000 2.905000 1.230000 3.075000 ;
      RECT 1.060000 3.265000 1.230000 3.435000 ;
      RECT 1.060000 3.625000 1.230000 3.795000 ;
      RECT 1.490000 1.105000 1.660000 1.275000 ;
      RECT 1.490000 1.465000 1.660000 1.635000 ;
      RECT 1.490000 1.825000 1.660000 1.995000 ;
      RECT 1.490000 2.185000 1.660000 2.355000 ;
      RECT 1.490000 2.545000 1.660000 2.715000 ;
      RECT 1.490000 2.905000 1.660000 3.075000 ;
      RECT 1.490000 3.265000 1.660000 3.435000 ;
      RECT 1.490000 3.625000 1.660000 3.795000 ;
      RECT 1.920000 1.105000 2.090000 1.275000 ;
      RECT 1.920000 1.465000 2.090000 1.635000 ;
      RECT 1.920000 1.825000 2.090000 1.995000 ;
      RECT 1.920000 2.185000 2.090000 2.355000 ;
      RECT 1.920000 2.545000 2.090000 2.715000 ;
      RECT 1.920000 2.905000 2.090000 3.075000 ;
      RECT 1.920000 3.265000 2.090000 3.435000 ;
      RECT 1.920000 3.625000 2.090000 3.795000 ;
      RECT 2.350000 1.105000 2.520000 1.275000 ;
      RECT 2.350000 1.465000 2.520000 1.635000 ;
      RECT 2.350000 1.825000 2.520000 1.995000 ;
      RECT 2.350000 2.185000 2.520000 2.355000 ;
      RECT 2.350000 2.545000 2.520000 2.715000 ;
      RECT 2.350000 2.905000 2.520000 3.075000 ;
      RECT 2.350000 3.265000 2.520000 3.435000 ;
      RECT 2.350000 3.625000 2.520000 3.795000 ;
      RECT 2.780000 1.105000 2.950000 1.275000 ;
      RECT 2.780000 1.465000 2.950000 1.635000 ;
      RECT 2.780000 1.825000 2.950000 1.995000 ;
      RECT 2.780000 2.185000 2.950000 2.355000 ;
      RECT 2.780000 2.545000 2.950000 2.715000 ;
      RECT 2.780000 2.905000 2.950000 3.075000 ;
      RECT 2.780000 3.265000 2.950000 3.435000 ;
      RECT 2.780000 3.625000 2.950000 3.795000 ;
    LAYER met1 ;
      RECT 1.015000 1.045000 1.275000 3.855000 ;
      RECT 1.445000 1.045000 1.705000 3.855000 ;
      RECT 1.875000 1.045000 2.135000 3.855000 ;
      RECT 2.305000 1.045000 2.565000 3.855000 ;
      RECT 2.735000 1.045000 2.995000 3.855000 ;
    LAYER via ;
      RECT 1.015000 1.075000 1.275000 1.335000 ;
      RECT 1.015000 1.395000 1.275000 1.655000 ;
      RECT 1.015000 1.715000 1.275000 1.975000 ;
      RECT 1.015000 2.035000 1.275000 2.295000 ;
      RECT 1.445000 2.605000 1.705000 2.865000 ;
      RECT 1.445000 2.925000 1.705000 3.185000 ;
      RECT 1.445000 3.245000 1.705000 3.505000 ;
      RECT 1.445000 3.565000 1.705000 3.825000 ;
      RECT 1.875000 1.075000 2.135000 1.335000 ;
      RECT 1.875000 1.395000 2.135000 1.655000 ;
      RECT 1.875000 1.715000 2.135000 1.975000 ;
      RECT 1.875000 2.035000 2.135000 2.295000 ;
      RECT 2.305000 2.605000 2.565000 2.865000 ;
      RECT 2.305000 2.925000 2.565000 3.185000 ;
      RECT 2.305000 3.245000 2.565000 3.505000 ;
      RECT 2.305000 3.565000 2.565000 3.825000 ;
      RECT 2.735000 1.075000 2.995000 1.335000 ;
      RECT 2.735000 1.395000 2.995000 1.655000 ;
      RECT 2.735000 1.715000 2.995000 1.975000 ;
      RECT 2.735000 2.035000 2.995000 2.295000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15
END LIBRARY
