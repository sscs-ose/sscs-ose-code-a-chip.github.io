# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_aura_lvs_drc
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_aura_lvs_drc ;
  ORIGIN  0.000000  213.9700 ;
  SIZE  1555.530 BY  412.1700 ;
  PIN B_P
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 -205.320000 11.985000 -202.345000 ;
    END
  END B_P
  PIN D_P
    ANTENNADIFFAREA  3.886400 ;
    PORT
      LAYER met3 ;
        RECT 74.460000 -124.310000 80.885000 -123.665000 ;
        RECT 76.195000 -124.455000 76.525000 -124.310000 ;
        RECT 77.055000 -124.455000 77.385000 -124.310000 ;
    END
  END D_P
  PIN G
    ANTENNAGATEAREA  8.190000 ;
    PORT
      LAYER met1 ;
        RECT 68.260000 100.485000 72.550000 100.785000 ;
        RECT 72.180000 100.785000 72.550000 100.905000 ;
        RECT 72.180000 100.905000 85.210000 101.195000 ;
        RECT 84.840000 101.195000 85.210000 103.065000 ;
        RECT 84.840000 103.065000 97.335000 103.355000 ;
    END
  END G
  PIN G_P
    ANTENNAGATEAREA  4.164000 ;
    PORT
      LAYER met1 ;
        RECT 66.630000 -124.305000 70.790000 -124.015000 ;
        RECT 70.445000 -124.015000 70.790000 -123.445000 ;
        RECT 70.445000 -123.445000 79.720000 -123.155000 ;
        RECT 76.105000 -123.465000 77.475000 -123.445000 ;
        RECT 79.375000 -123.155000 79.720000 -122.145000 ;
        RECT 79.375000 -122.145000 85.050000 -121.855000 ;
        RECT 84.705000 -121.855000 85.050000 -120.110000 ;
        RECT 84.705000 -120.110000 87.235000 -119.820000 ;
    END
  END G_P
  PIN NWELL
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 8.650000 11.985000 11.625000 ;
    END
  END NWELL
  PIN S
    ANTENNADIFFAREA  10.98720 ;
    PORT
      LAYER met1 ;
        RECT 68.260000 99.265000 97.765000  99.565000 ;
        RECT 69.045000 99.565000 69.275000 100.310000 ;
        RECT 69.905000 99.565000 70.135000 100.310000 ;
        RECT 74.165000 99.565000 74.395000 100.655000 ;
        RECT 75.025000 99.565000 75.255000 100.655000 ;
        RECT 76.885000 99.565000 77.115000 100.655000 ;
        RECT 77.745000 99.565000 77.975000 100.655000 ;
        RECT 78.605000 99.565000 78.835000 100.655000 ;
        RECT 80.100000 99.565000 80.330000 100.655000 ;
        RECT 80.960000 99.565000 81.190000 100.655000 ;
        RECT 81.820000 99.565000 82.050000 100.655000 ;
        RECT 82.680000 99.565000 82.910000 100.655000 ;
        RECT 83.540000 99.565000 83.770000 100.655000 ;
        RECT 86.605000 99.565000 86.835000 102.815000 ;
        RECT 87.465000 99.565000 87.695000 102.815000 ;
        RECT 90.095000 99.565000 90.325000 102.815000 ;
        RECT 90.955000 99.565000 91.185000 102.815000 ;
        RECT 91.815000 99.565000 92.045000 102.815000 ;
        RECT 94.095000 99.565000 94.325000 102.815000 ;
        RECT 94.955000 99.565000 95.185000 102.815000 ;
        RECT 95.815000 99.565000 96.045000 102.815000 ;
        RECT 96.675000 99.565000 96.905000 102.815000 ;
        RECT 97.535000 99.565000 97.765000 102.815000 ;
    END
  END S
  PIN S_P
    ANTENNADIFFAREA  6.936400 ;
    PORT
      LAYER met1 ;
        RECT 66.630000 -125.955000 87.455000 -125.655000 ;
        RECT 68.055000 -125.655000 68.285000 -124.565000 ;
        RECT 68.915000 -125.655000 69.145000 -124.565000 ;
        RECT 71.905000 -125.655000 72.135000 -123.660000 ;
        RECT 72.765000 -125.655000 72.995000 -123.660000 ;
        RECT 75.815000 -125.655000 76.045000 -123.725000 ;
        RECT 76.675000 -125.655000 76.905000 -123.725000 ;
        RECT 77.535000 -125.655000 77.765000 -123.725000 ;
        RECT 81.950000 -125.655000 82.180000 -122.405000 ;
        RECT 82.810000 -125.655000 83.040000 -122.405000 ;
        RECT 86.365000 -125.655000 86.595000 -120.300000 ;
        RECT 87.225000 -125.655000 87.455000 -120.300000 ;
    END
  END S_P
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 60.140000 90.690000 62.950000 93.665000 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 75.895000  99.965000 86.220000 100.685000 ;
        RECT 77.265000  99.915000 77.595000  99.965000 ;
        RECT 78.125000  99.915000 78.455000  99.965000 ;
        RECT 80.480000  99.915000 80.810000  99.965000 ;
        RECT 81.340000  99.915000 81.670000  99.965000 ;
        RECT 82.200000  99.915000 82.530000  99.965000 ;
        RECT 83.060000  99.915000 83.390000  99.965000 ;
        RECT 85.830000 100.685000 86.220000 102.875000 ;
        RECT 88.780000 102.075000 97.385000 102.875000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 68.085000 -125.255000 68.255000 -124.565000 ;
      RECT 68.265000 -124.335000 68.935000 -123.995000 ;
      RECT 68.515000 -125.255000 68.685000 -124.565000 ;
      RECT 68.945000 -125.255000 69.115000 -124.565000 ;
      RECT 69.075000   99.965000 69.245000  100.295000 ;
      RECT 69.255000  100.465000 69.925000  100.795000 ;
      RECT 69.505000   99.965000 69.675000  100.295000 ;
      RECT 69.935000   99.965000 70.105000  100.295000 ;
      RECT 71.935000 -125.330000 72.105000 -123.660000 ;
      RECT 72.115000 -123.465000 72.785000 -123.135000 ;
      RECT 72.365000 -125.330000 72.535000 -123.660000 ;
      RECT 72.795000 -125.330000 72.965000 -123.660000 ;
      RECT 74.195000   99.965000 74.365000  100.655000 ;
      RECT 74.375000  100.885000 75.045000  101.215000 ;
      RECT 74.625000   99.965000 74.795000  100.655000 ;
      RECT 75.055000   99.965000 75.225000  100.655000 ;
      RECT 75.845000 -125.255000 76.015000 -123.725000 ;
      RECT 76.115000 -123.495000 77.465000 -123.155000 ;
      RECT 76.275000 -125.255000 76.445000 -123.725000 ;
      RECT 76.705000 -125.255000 76.875000 -123.725000 ;
      RECT 76.915000   99.965000 77.085000  100.655000 ;
      RECT 77.135000 -125.255000 77.305000 -123.725000 ;
      RECT 77.185000  100.885000 78.535000  101.215000 ;
      RECT 77.345000   99.965000 77.515000  100.655000 ;
      RECT 77.565000 -125.255000 77.735000 -123.725000 ;
      RECT 77.775000   99.965000 77.945000  100.655000 ;
      RECT 78.205000   99.965000 78.375000  100.655000 ;
      RECT 78.635000   99.965000 78.805000  100.655000 ;
      RECT 80.130000   99.965000 80.300000  100.655000 ;
      RECT 80.560000   99.965000 80.730000  100.655000 ;
      RECT 80.580000  100.885000 83.290000  101.215000 ;
      RECT 80.990000   99.965000 81.160000  100.655000 ;
      RECT 81.420000   99.965000 81.590000  100.655000 ;
      RECT 81.850000   99.965000 82.020000  100.655000 ;
      RECT 81.980000 -125.275000 82.150000 -122.405000 ;
      RECT 82.160000 -122.175000 82.830000 -121.835000 ;
      RECT 82.280000   99.965000 82.450000  100.655000 ;
      RECT 82.410000 -125.255000 82.580000 -122.405000 ;
      RECT 82.710000   99.965000 82.880000  100.655000 ;
      RECT 82.840000 -125.255000 83.010000 -122.405000 ;
      RECT 83.140000   99.965000 83.310000  100.655000 ;
      RECT 83.570000   99.965000 83.740000  100.655000 ;
      RECT 86.395000 -125.290000 86.565000 -120.300000 ;
      RECT 86.575000 -120.130000 87.245000 -119.800000 ;
      RECT 86.635000   99.945000 86.805000  102.815000 ;
      RECT 86.815000  103.045000 87.485000  103.375000 ;
      RECT 86.825000 -125.290000 86.995000 -120.300000 ;
      RECT 87.065000   99.965000 87.235000  102.815000 ;
      RECT 87.255000 -125.290000 87.425000 -120.300000 ;
      RECT 87.495000   99.965000 87.665000  102.815000 ;
      RECT 90.125000   99.965000 90.295000  102.815000 ;
      RECT 90.395000  103.045000 91.745000  103.375000 ;
      RECT 90.555000   99.965000 90.725000  102.815000 ;
      RECT 90.985000   99.965000 91.155000  102.815000 ;
      RECT 91.415000   99.965000 91.585000  102.815000 ;
      RECT 91.845000   99.965000 92.015000  102.815000 ;
      RECT 94.125000   99.965000 94.295000  102.815000 ;
      RECT 94.555000   99.965000 94.725000  102.815000 ;
      RECT 94.575000  103.045000 97.285000  103.375000 ;
      RECT 94.985000   99.965000 95.155000  102.815000 ;
      RECT 95.415000   99.965000 95.585000  102.815000 ;
      RECT 95.845000   99.965000 96.015000  102.815000 ;
      RECT 96.275000   99.965000 96.445000  102.815000 ;
      RECT 96.705000   99.965000 96.875000  102.815000 ;
      RECT 97.135000   99.965000 97.305000  102.815000 ;
      RECT 97.565000   99.965000 97.735000  102.815000 ;
    LAYER mcon ;
      RECT 68.085000 -125.175000 68.255000 -125.005000 ;
      RECT 68.085000 -124.815000 68.255000 -124.645000 ;
      RECT 68.335000 -124.245000 68.505000 -124.075000 ;
      RECT 68.515000 -125.175000 68.685000 -125.005000 ;
      RECT 68.515000 -124.815000 68.685000 -124.645000 ;
      RECT 68.695000 -124.245000 68.865000 -124.075000 ;
      RECT 68.945000 -125.175000 69.115000 -125.005000 ;
      RECT 68.945000 -124.815000 69.115000 -124.645000 ;
      RECT 69.075000  100.045000 69.245000  100.215000 ;
      RECT 69.325000  100.545000 69.495000  100.715000 ;
      RECT 69.505000  100.045000 69.675000  100.215000 ;
      RECT 69.685000  100.545000 69.855000  100.715000 ;
      RECT 69.935000  100.045000 70.105000  100.215000 ;
      RECT 71.935000 -125.115000 72.105000 -124.945000 ;
      RECT 71.935000 -124.755000 72.105000 -124.585000 ;
      RECT 71.935000 -124.395000 72.105000 -124.225000 ;
      RECT 71.935000 -124.035000 72.105000 -123.865000 ;
      RECT 72.185000 -123.385000 72.355000 -123.215000 ;
      RECT 72.365000 -125.115000 72.535000 -124.945000 ;
      RECT 72.365000 -124.755000 72.535000 -124.585000 ;
      RECT 72.365000 -124.395000 72.535000 -124.225000 ;
      RECT 72.365000 -124.035000 72.535000 -123.865000 ;
      RECT 72.545000 -123.385000 72.715000 -123.215000 ;
      RECT 72.795000 -125.115000 72.965000 -124.945000 ;
      RECT 72.795000 -124.755000 72.965000 -124.585000 ;
      RECT 72.795000 -124.395000 72.965000 -124.225000 ;
      RECT 72.795000 -124.035000 72.965000 -123.865000 ;
      RECT 74.195000  100.045000 74.365000  100.215000 ;
      RECT 74.195000  100.405000 74.365000  100.575000 ;
      RECT 74.445000  100.965000 74.615000  101.135000 ;
      RECT 74.625000  100.045000 74.795000  100.215000 ;
      RECT 74.625000  100.405000 74.795000  100.575000 ;
      RECT 74.805000  100.965000 74.975000  101.135000 ;
      RECT 75.055000  100.045000 75.225000  100.215000 ;
      RECT 75.055000  100.405000 75.225000  100.575000 ;
      RECT 75.845000 -125.115000 76.015000 -124.945000 ;
      RECT 75.845000 -124.755000 76.015000 -124.585000 ;
      RECT 75.845000 -124.395000 76.015000 -124.225000 ;
      RECT 75.845000 -124.035000 76.015000 -123.865000 ;
      RECT 76.165000 -123.405000 76.335000 -123.235000 ;
      RECT 76.275000 -125.115000 76.445000 -124.945000 ;
      RECT 76.275000 -124.755000 76.445000 -124.585000 ;
      RECT 76.275000 -124.395000 76.445000 -124.225000 ;
      RECT 76.275000 -124.035000 76.445000 -123.865000 ;
      RECT 76.525000 -123.405000 76.695000 -123.235000 ;
      RECT 76.705000 -125.115000 76.875000 -124.945000 ;
      RECT 76.705000 -124.755000 76.875000 -124.585000 ;
      RECT 76.705000 -124.395000 76.875000 -124.225000 ;
      RECT 76.705000 -124.035000 76.875000 -123.865000 ;
      RECT 76.885000 -123.405000 77.055000 -123.235000 ;
      RECT 76.915000  100.045000 77.085000  100.215000 ;
      RECT 76.915000  100.405000 77.085000  100.575000 ;
      RECT 77.135000 -125.115000 77.305000 -124.945000 ;
      RECT 77.135000 -124.755000 77.305000 -124.585000 ;
      RECT 77.135000 -124.395000 77.305000 -124.225000 ;
      RECT 77.135000 -124.035000 77.305000 -123.865000 ;
      RECT 77.235000  100.965000 77.405000  101.135000 ;
      RECT 77.245000 -123.405000 77.415000 -123.235000 ;
      RECT 77.345000  100.045000 77.515000  100.215000 ;
      RECT 77.345000  100.405000 77.515000  100.575000 ;
      RECT 77.565000 -125.115000 77.735000 -124.945000 ;
      RECT 77.565000 -124.755000 77.735000 -124.585000 ;
      RECT 77.565000 -124.395000 77.735000 -124.225000 ;
      RECT 77.565000 -124.035000 77.735000 -123.865000 ;
      RECT 77.595000  100.965000 77.765000  101.135000 ;
      RECT 77.775000  100.045000 77.945000  100.215000 ;
      RECT 77.775000  100.405000 77.945000  100.575000 ;
      RECT 77.955000  100.965000 78.125000  101.135000 ;
      RECT 78.205000  100.045000 78.375000  100.215000 ;
      RECT 78.205000  100.405000 78.375000  100.575000 ;
      RECT 78.315000  100.965000 78.485000  101.135000 ;
      RECT 78.635000  100.045000 78.805000  100.215000 ;
      RECT 78.635000  100.405000 78.805000  100.575000 ;
      RECT 80.130000  100.045000 80.300000  100.215000 ;
      RECT 80.130000  100.405000 80.300000  100.575000 ;
      RECT 80.560000  100.045000 80.730000  100.215000 ;
      RECT 80.560000  100.405000 80.730000  100.575000 ;
      RECT 80.590000  100.965000 80.760000  101.135000 ;
      RECT 80.950000  100.965000 81.120000  101.135000 ;
      RECT 80.990000  100.045000 81.160000  100.215000 ;
      RECT 80.990000  100.405000 81.160000  100.575000 ;
      RECT 81.310000  100.965000 81.480000  101.135000 ;
      RECT 81.420000  100.045000 81.590000  100.215000 ;
      RECT 81.420000  100.405000 81.590000  100.575000 ;
      RECT 81.670000  100.965000 81.840000  101.135000 ;
      RECT 81.850000  100.045000 82.020000  100.215000 ;
      RECT 81.850000  100.405000 82.020000  100.575000 ;
      RECT 81.980000 -125.175000 82.150000 -125.005000 ;
      RECT 81.980000 -124.815000 82.150000 -124.645000 ;
      RECT 81.980000 -124.455000 82.150000 -124.285000 ;
      RECT 81.980000 -124.095000 82.150000 -123.925000 ;
      RECT 81.980000 -123.735000 82.150000 -123.565000 ;
      RECT 81.980000 -123.375000 82.150000 -123.205000 ;
      RECT 81.980000 -123.015000 82.150000 -122.845000 ;
      RECT 81.980000 -122.655000 82.150000 -122.485000 ;
      RECT 82.030000  100.965000 82.200000  101.135000 ;
      RECT 82.230000 -122.085000 82.400000 -121.915000 ;
      RECT 82.280000  100.045000 82.450000  100.215000 ;
      RECT 82.280000  100.405000 82.450000  100.575000 ;
      RECT 82.390000  100.965000 82.560000  101.135000 ;
      RECT 82.410000 -125.175000 82.580000 -125.005000 ;
      RECT 82.410000 -124.815000 82.580000 -124.645000 ;
      RECT 82.410000 -124.455000 82.580000 -124.285000 ;
      RECT 82.410000 -124.095000 82.580000 -123.925000 ;
      RECT 82.410000 -123.735000 82.580000 -123.565000 ;
      RECT 82.410000 -123.375000 82.580000 -123.205000 ;
      RECT 82.410000 -123.015000 82.580000 -122.845000 ;
      RECT 82.410000 -122.655000 82.580000 -122.485000 ;
      RECT 82.590000 -122.085000 82.760000 -121.915000 ;
      RECT 82.710000  100.045000 82.880000  100.215000 ;
      RECT 82.710000  100.405000 82.880000  100.575000 ;
      RECT 82.750000  100.965000 82.920000  101.135000 ;
      RECT 82.840000 -125.175000 83.010000 -125.005000 ;
      RECT 82.840000 -124.815000 83.010000 -124.645000 ;
      RECT 82.840000 -124.455000 83.010000 -124.285000 ;
      RECT 82.840000 -124.095000 83.010000 -123.925000 ;
      RECT 82.840000 -123.735000 83.010000 -123.565000 ;
      RECT 82.840000 -123.375000 83.010000 -123.205000 ;
      RECT 82.840000 -123.015000 83.010000 -122.845000 ;
      RECT 82.840000 -122.655000 83.010000 -122.485000 ;
      RECT 83.110000  100.965000 83.280000  101.135000 ;
      RECT 83.140000  100.045000 83.310000  100.215000 ;
      RECT 83.140000  100.405000 83.310000  100.575000 ;
      RECT 83.570000  100.045000 83.740000  100.215000 ;
      RECT 83.570000  100.405000 83.740000  100.575000 ;
      RECT 86.395000 -125.035000 86.565000 -124.865000 ;
      RECT 86.395000 -124.675000 86.565000 -124.505000 ;
      RECT 86.395000 -124.315000 86.565000 -124.145000 ;
      RECT 86.395000 -123.955000 86.565000 -123.785000 ;
      RECT 86.395000 -123.595000 86.565000 -123.425000 ;
      RECT 86.395000 -123.235000 86.565000 -123.065000 ;
      RECT 86.395000 -122.875000 86.565000 -122.705000 ;
      RECT 86.395000 -122.515000 86.565000 -122.345000 ;
      RECT 86.395000 -122.155000 86.565000 -121.985000 ;
      RECT 86.395000 -121.795000 86.565000 -121.625000 ;
      RECT 86.395000 -121.435000 86.565000 -121.265000 ;
      RECT 86.395000 -121.075000 86.565000 -120.905000 ;
      RECT 86.395000 -120.715000 86.565000 -120.545000 ;
      RECT 86.635000  100.045000 86.805000  100.215000 ;
      RECT 86.635000  100.405000 86.805000  100.575000 ;
      RECT 86.635000  100.765000 86.805000  100.935000 ;
      RECT 86.635000  101.125000 86.805000  101.295000 ;
      RECT 86.635000  101.485000 86.805000  101.655000 ;
      RECT 86.635000  101.845000 86.805000  102.015000 ;
      RECT 86.635000  102.205000 86.805000  102.375000 ;
      RECT 86.635000  102.565000 86.805000  102.735000 ;
      RECT 86.645000 -120.050000 86.815000 -119.880000 ;
      RECT 86.825000 -125.035000 86.995000 -124.865000 ;
      RECT 86.825000 -124.675000 86.995000 -124.505000 ;
      RECT 86.825000 -124.315000 86.995000 -124.145000 ;
      RECT 86.825000 -123.955000 86.995000 -123.785000 ;
      RECT 86.825000 -123.595000 86.995000 -123.425000 ;
      RECT 86.825000 -123.235000 86.995000 -123.065000 ;
      RECT 86.825000 -122.875000 86.995000 -122.705000 ;
      RECT 86.825000 -122.515000 86.995000 -122.345000 ;
      RECT 86.825000 -122.155000 86.995000 -121.985000 ;
      RECT 86.825000 -121.795000 86.995000 -121.625000 ;
      RECT 86.825000 -121.435000 86.995000 -121.265000 ;
      RECT 86.825000 -121.075000 86.995000 -120.905000 ;
      RECT 86.825000 -120.715000 86.995000 -120.545000 ;
      RECT 86.885000  103.125000 87.055000  103.295000 ;
      RECT 87.005000 -120.050000 87.175000 -119.880000 ;
      RECT 87.065000  100.045000 87.235000  100.215000 ;
      RECT 87.065000  100.405000 87.235000  100.575000 ;
      RECT 87.065000  100.765000 87.235000  100.935000 ;
      RECT 87.065000  101.125000 87.235000  101.295000 ;
      RECT 87.065000  101.485000 87.235000  101.655000 ;
      RECT 87.065000  101.845000 87.235000  102.015000 ;
      RECT 87.065000  102.205000 87.235000  102.375000 ;
      RECT 87.065000  102.565000 87.235000  102.735000 ;
      RECT 87.245000  103.125000 87.415000  103.295000 ;
      RECT 87.255000 -125.035000 87.425000 -124.865000 ;
      RECT 87.255000 -124.675000 87.425000 -124.505000 ;
      RECT 87.255000 -124.315000 87.425000 -124.145000 ;
      RECT 87.255000 -123.955000 87.425000 -123.785000 ;
      RECT 87.255000 -123.595000 87.425000 -123.425000 ;
      RECT 87.255000 -123.235000 87.425000 -123.065000 ;
      RECT 87.255000 -122.875000 87.425000 -122.705000 ;
      RECT 87.255000 -122.515000 87.425000 -122.345000 ;
      RECT 87.255000 -122.155000 87.425000 -121.985000 ;
      RECT 87.255000 -121.795000 87.425000 -121.625000 ;
      RECT 87.255000 -121.435000 87.425000 -121.265000 ;
      RECT 87.255000 -121.075000 87.425000 -120.905000 ;
      RECT 87.255000 -120.715000 87.425000 -120.545000 ;
      RECT 87.495000  100.045000 87.665000  100.215000 ;
      RECT 87.495000  100.405000 87.665000  100.575000 ;
      RECT 87.495000  100.765000 87.665000  100.935000 ;
      RECT 87.495000  101.125000 87.665000  101.295000 ;
      RECT 87.495000  101.485000 87.665000  101.655000 ;
      RECT 87.495000  101.845000 87.665000  102.015000 ;
      RECT 87.495000  102.205000 87.665000  102.375000 ;
      RECT 87.495000  102.565000 87.665000  102.735000 ;
      RECT 90.125000  100.045000 90.295000  100.215000 ;
      RECT 90.125000  100.405000 90.295000  100.575000 ;
      RECT 90.125000  100.765000 90.295000  100.935000 ;
      RECT 90.125000  101.125000 90.295000  101.295000 ;
      RECT 90.125000  101.485000 90.295000  101.655000 ;
      RECT 90.125000  101.845000 90.295000  102.015000 ;
      RECT 90.125000  102.205000 90.295000  102.375000 ;
      RECT 90.125000  102.565000 90.295000  102.735000 ;
      RECT 90.445000  103.125000 90.615000  103.295000 ;
      RECT 90.555000  100.045000 90.725000  100.215000 ;
      RECT 90.555000  100.405000 90.725000  100.575000 ;
      RECT 90.555000  100.765000 90.725000  100.935000 ;
      RECT 90.555000  101.125000 90.725000  101.295000 ;
      RECT 90.555000  101.485000 90.725000  101.655000 ;
      RECT 90.555000  101.845000 90.725000  102.015000 ;
      RECT 90.555000  102.205000 90.725000  102.375000 ;
      RECT 90.555000  102.565000 90.725000  102.735000 ;
      RECT 90.805000  103.125000 90.975000  103.295000 ;
      RECT 90.985000  100.045000 91.155000  100.215000 ;
      RECT 90.985000  100.405000 91.155000  100.575000 ;
      RECT 90.985000  100.765000 91.155000  100.935000 ;
      RECT 90.985000  101.125000 91.155000  101.295000 ;
      RECT 90.985000  101.485000 91.155000  101.655000 ;
      RECT 90.985000  101.845000 91.155000  102.015000 ;
      RECT 90.985000  102.205000 91.155000  102.375000 ;
      RECT 90.985000  102.565000 91.155000  102.735000 ;
      RECT 91.165000  103.125000 91.335000  103.295000 ;
      RECT 91.415000  100.045000 91.585000  100.215000 ;
      RECT 91.415000  100.405000 91.585000  100.575000 ;
      RECT 91.415000  100.765000 91.585000  100.935000 ;
      RECT 91.415000  101.125000 91.585000  101.295000 ;
      RECT 91.415000  101.485000 91.585000  101.655000 ;
      RECT 91.415000  101.845000 91.585000  102.015000 ;
      RECT 91.415000  102.205000 91.585000  102.375000 ;
      RECT 91.415000  102.565000 91.585000  102.735000 ;
      RECT 91.525000  103.125000 91.695000  103.295000 ;
      RECT 91.845000  100.045000 92.015000  100.215000 ;
      RECT 91.845000  100.405000 92.015000  100.575000 ;
      RECT 91.845000  100.765000 92.015000  100.935000 ;
      RECT 91.845000  101.125000 92.015000  101.295000 ;
      RECT 91.845000  101.485000 92.015000  101.655000 ;
      RECT 91.845000  101.845000 92.015000  102.015000 ;
      RECT 91.845000  102.205000 92.015000  102.375000 ;
      RECT 91.845000  102.565000 92.015000  102.735000 ;
      RECT 94.125000  100.045000 94.295000  100.215000 ;
      RECT 94.125000  100.405000 94.295000  100.575000 ;
      RECT 94.125000  100.765000 94.295000  100.935000 ;
      RECT 94.125000  101.125000 94.295000  101.295000 ;
      RECT 94.125000  101.485000 94.295000  101.655000 ;
      RECT 94.125000  101.845000 94.295000  102.015000 ;
      RECT 94.125000  102.205000 94.295000  102.375000 ;
      RECT 94.125000  102.565000 94.295000  102.735000 ;
      RECT 94.555000  100.045000 94.725000  100.215000 ;
      RECT 94.555000  100.405000 94.725000  100.575000 ;
      RECT 94.555000  100.765000 94.725000  100.935000 ;
      RECT 94.555000  101.125000 94.725000  101.295000 ;
      RECT 94.555000  101.485000 94.725000  101.655000 ;
      RECT 94.555000  101.845000 94.725000  102.015000 ;
      RECT 94.555000  102.205000 94.725000  102.375000 ;
      RECT 94.555000  102.565000 94.725000  102.735000 ;
      RECT 94.585000  103.125000 94.755000  103.295000 ;
      RECT 94.945000  103.125000 95.115000  103.295000 ;
      RECT 94.985000  100.045000 95.155000  100.215000 ;
      RECT 94.985000  100.405000 95.155000  100.575000 ;
      RECT 94.985000  100.765000 95.155000  100.935000 ;
      RECT 94.985000  101.125000 95.155000  101.295000 ;
      RECT 94.985000  101.485000 95.155000  101.655000 ;
      RECT 94.985000  101.845000 95.155000  102.015000 ;
      RECT 94.985000  102.205000 95.155000  102.375000 ;
      RECT 94.985000  102.565000 95.155000  102.735000 ;
      RECT 95.305000  103.125000 95.475000  103.295000 ;
      RECT 95.415000  100.045000 95.585000  100.215000 ;
      RECT 95.415000  100.405000 95.585000  100.575000 ;
      RECT 95.415000  100.765000 95.585000  100.935000 ;
      RECT 95.415000  101.125000 95.585000  101.295000 ;
      RECT 95.415000  101.485000 95.585000  101.655000 ;
      RECT 95.415000  101.845000 95.585000  102.015000 ;
      RECT 95.415000  102.205000 95.585000  102.375000 ;
      RECT 95.415000  102.565000 95.585000  102.735000 ;
      RECT 95.665000  103.125000 95.835000  103.295000 ;
      RECT 95.845000  100.045000 96.015000  100.215000 ;
      RECT 95.845000  100.405000 96.015000  100.575000 ;
      RECT 95.845000  100.765000 96.015000  100.935000 ;
      RECT 95.845000  101.125000 96.015000  101.295000 ;
      RECT 95.845000  101.485000 96.015000  101.655000 ;
      RECT 95.845000  101.845000 96.015000  102.015000 ;
      RECT 95.845000  102.205000 96.015000  102.375000 ;
      RECT 95.845000  102.565000 96.015000  102.735000 ;
      RECT 96.025000  103.125000 96.195000  103.295000 ;
      RECT 96.275000  100.045000 96.445000  100.215000 ;
      RECT 96.275000  100.405000 96.445000  100.575000 ;
      RECT 96.275000  100.765000 96.445000  100.935000 ;
      RECT 96.275000  101.125000 96.445000  101.295000 ;
      RECT 96.275000  101.485000 96.445000  101.655000 ;
      RECT 96.275000  101.845000 96.445000  102.015000 ;
      RECT 96.275000  102.205000 96.445000  102.375000 ;
      RECT 96.275000  102.565000 96.445000  102.735000 ;
      RECT 96.385000  103.125000 96.555000  103.295000 ;
      RECT 96.705000  100.045000 96.875000  100.215000 ;
      RECT 96.705000  100.405000 96.875000  100.575000 ;
      RECT 96.705000  100.765000 96.875000  100.935000 ;
      RECT 96.705000  101.125000 96.875000  101.295000 ;
      RECT 96.705000  101.485000 96.875000  101.655000 ;
      RECT 96.705000  101.845000 96.875000  102.015000 ;
      RECT 96.705000  102.205000 96.875000  102.375000 ;
      RECT 96.705000  102.565000 96.875000  102.735000 ;
      RECT 96.745000  103.125000 96.915000  103.295000 ;
      RECT 97.105000  103.125000 97.275000  103.295000 ;
      RECT 97.135000  100.045000 97.305000  100.215000 ;
      RECT 97.135000  100.405000 97.305000  100.575000 ;
      RECT 97.135000  100.765000 97.305000  100.935000 ;
      RECT 97.135000  101.125000 97.305000  101.295000 ;
      RECT 97.135000  101.485000 97.305000  101.655000 ;
      RECT 97.135000  101.845000 97.305000  102.015000 ;
      RECT 97.135000  102.205000 97.305000  102.375000 ;
      RECT 97.135000  102.565000 97.305000  102.735000 ;
      RECT 97.565000  100.045000 97.735000  100.215000 ;
      RECT 97.565000  100.405000 97.735000  100.575000 ;
      RECT 97.565000  100.765000 97.735000  100.935000 ;
      RECT 97.565000  101.125000 97.735000  101.295000 ;
      RECT 97.565000  101.485000 97.735000  101.655000 ;
      RECT 97.565000  101.845000 97.735000  102.015000 ;
      RECT 97.565000  102.205000 97.735000  102.375000 ;
      RECT 97.565000  102.565000 97.735000  102.735000 ;
    LAYER met1 ;
      RECT 68.470000 -125.255000 68.730000 -124.565000 ;
      RECT 69.460000   99.965000 69.720000  100.310000 ;
      RECT 72.320000 -125.330000 72.580000 -123.660000 ;
      RECT 74.580000   99.965000 74.840000  100.655000 ;
      RECT 76.230000 -125.255000 76.490000 -123.725000 ;
      RECT 77.090000 -125.255000 77.350000 -123.725000 ;
      RECT 77.300000   99.965000 77.560000  100.655000 ;
      RECT 78.160000   99.965000 78.420000  100.655000 ;
      RECT 80.515000   99.965000 80.775000  100.655000 ;
      RECT 81.375000   99.965000 81.635000  100.655000 ;
      RECT 82.235000   99.965000 82.495000  100.655000 ;
      RECT 82.365000 -125.255000 82.625000 -122.405000 ;
      RECT 83.095000   99.965000 83.355000  100.655000 ;
      RECT 86.780000 -125.290000 87.040000 -120.300000 ;
      RECT 87.020000   99.965000 87.280000  102.815000 ;
      RECT 90.510000   99.965000 90.770000  102.815000 ;
      RECT 91.370000   99.965000 91.630000  102.815000 ;
      RECT 94.510000   99.965000 94.770000  102.815000 ;
      RECT 95.370000   99.965000 95.630000  102.815000 ;
      RECT 96.230000   99.965000 96.490000  102.815000 ;
      RECT 97.090000   99.965000 97.350000  102.815000 ;
    LAYER met2 ;
      RECT 66.635000 -125.230000 71.490000 -124.590000 ;
      RECT 68.260000   99.965000 76.300000  100.310000 ;
      RECT 71.125000 -124.590000 71.490000 -124.305000 ;
      RECT 71.125000 -124.305000 75.085000 -123.665000 ;
      RECT 74.580000  100.310000 74.840000  100.630000 ;
      RECT 76.195000 -124.455000 76.525000 -123.685000 ;
      RECT 77.055000 -124.455000 77.385000 -123.685000 ;
      RECT 77.265000   99.915000 77.595000  100.685000 ;
      RECT 78.125000   99.915000 78.455000  100.685000 ;
      RECT 80.340000 -124.310000 80.885000 -123.070000 ;
      RECT 80.340000 -123.070000 85.850000 -122.430000 ;
      RECT 80.480000   99.915000 80.810000  100.685000 ;
      RECT 81.340000   99.915000 81.670000  100.685000 ;
      RECT 82.200000   99.915000 82.530000  100.685000 ;
      RECT 83.060000   99.915000 83.390000  100.685000 ;
      RECT 85.305000 -122.430000 85.850000 -120.950000 ;
      RECT 85.305000 -120.950000 87.040000 -120.310000 ;
      RECT 85.830000  102.150000 89.290000  102.875000 ;
      RECT 90.475000  102.075000 90.805000  102.845000 ;
      RECT 91.335000  102.075000 91.665000  102.845000 ;
      RECT 94.475000  102.075000 94.805000  102.845000 ;
      RECT 95.335000  102.075000 95.665000  102.845000 ;
      RECT 96.195000  102.075000 96.525000  102.845000 ;
      RECT 97.055000  102.075000 97.385000  102.845000 ;
    LAYER via ;
      RECT 68.470000 -125.200000 68.730000 -124.940000 ;
      RECT 68.470000 -124.880000 68.730000 -124.620000 ;
      RECT 69.460000  100.020000 69.720000  100.280000 ;
      RECT 72.320000 -124.275000 72.580000 -124.015000 ;
      RECT 72.320000 -123.955000 72.580000 -123.695000 ;
      RECT 74.580000  100.020000 74.840000  100.280000 ;
      RECT 74.580000  100.340000 74.840000  100.600000 ;
      RECT 76.230000 -124.360000 76.490000 -124.100000 ;
      RECT 76.230000 -124.040000 76.490000 -123.780000 ;
      RECT 77.090000 -124.360000 77.350000 -124.100000 ;
      RECT 77.090000 -124.040000 77.350000 -123.780000 ;
      RECT 77.300000  100.005000 77.560000  100.265000 ;
      RECT 77.300000  100.325000 77.560000  100.585000 ;
      RECT 78.160000  100.005000 78.420000  100.265000 ;
      RECT 78.160000  100.325000 78.420000  100.585000 ;
      RECT 80.515000  100.020000 80.775000  100.280000 ;
      RECT 80.515000  100.340000 80.775000  100.600000 ;
      RECT 81.375000  100.010000 81.635000  100.270000 ;
      RECT 81.375000  100.330000 81.635000  100.590000 ;
      RECT 82.235000  100.010000 82.495000  100.270000 ;
      RECT 82.235000  100.330000 82.495000  100.590000 ;
      RECT 82.365000 -123.040000 82.625000 -122.780000 ;
      RECT 82.365000 -122.720000 82.625000 -122.460000 ;
      RECT 83.095000  100.010000 83.355000  100.270000 ;
      RECT 83.095000  100.330000 83.355000  100.590000 ;
      RECT 86.780000 -120.920000 87.040000 -120.660000 ;
      RECT 86.780000 -120.600000 87.040000 -120.340000 ;
      RECT 87.020000  102.180000 87.280000  102.440000 ;
      RECT 87.020000  102.500000 87.280000  102.760000 ;
      RECT 90.510000  102.165000 90.770000  102.425000 ;
      RECT 90.510000  102.485000 90.770000  102.745000 ;
      RECT 91.370000  102.165000 91.630000  102.425000 ;
      RECT 91.370000  102.485000 91.630000  102.745000 ;
      RECT 94.510000  102.170000 94.770000  102.430000 ;
      RECT 94.510000  102.490000 94.770000  102.750000 ;
      RECT 95.370000  102.170000 95.630000  102.430000 ;
      RECT 95.370000  102.490000 95.630000  102.750000 ;
      RECT 96.230000  102.170000 96.490000  102.430000 ;
      RECT 96.230000  102.490000 96.490000  102.750000 ;
      RECT 97.090000  102.170000 97.350000  102.430000 ;
      RECT 97.090000  102.490000 97.350000  102.750000 ;
    LAYER via2 ;
      RECT 74.565000 -124.155000 74.845000 -123.875000 ;
      RECT 75.945000  100.000000 76.225000  100.280000 ;
      RECT 76.220000 -124.410000 76.500000 -124.130000 ;
      RECT 76.220000 -124.010000 76.500000 -123.730000 ;
      RECT 77.080000 -124.410000 77.360000 -124.130000 ;
      RECT 77.080000 -124.010000 77.360000 -123.730000 ;
      RECT 77.290000   99.960000 77.570000  100.240000 ;
      RECT 77.290000  100.360000 77.570000  100.640000 ;
      RECT 78.150000   99.960000 78.430000  100.240000 ;
      RECT 78.150000  100.360000 78.430000  100.640000 ;
      RECT 80.490000 -124.155000 80.770000 -123.875000 ;
      RECT 80.505000   99.960000 80.785000  100.240000 ;
      RECT 80.505000  100.360000 80.785000  100.640000 ;
      RECT 81.365000   99.960000 81.645000  100.240000 ;
      RECT 81.365000  100.360000 81.645000  100.640000 ;
      RECT 82.225000   99.960000 82.505000  100.240000 ;
      RECT 82.225000  100.360000 82.505000  100.640000 ;
      RECT 83.085000   99.960000 83.365000  100.240000 ;
      RECT 83.085000  100.360000 83.365000  100.640000 ;
      RECT 85.885000  102.530000 86.165000  102.810000 ;
      RECT 88.885000  102.375000 89.165000  102.655000 ;
      RECT 90.500000  102.120000 90.780000  102.400000 ;
      RECT 90.500000  102.520000 90.780000  102.800000 ;
      RECT 91.360000  102.120000 91.640000  102.400000 ;
      RECT 91.360000  102.520000 91.640000  102.800000 ;
      RECT 94.500000  102.120000 94.780000  102.400000 ;
      RECT 94.500000  102.520000 94.780000  102.800000 ;
      RECT 95.360000  102.120000 95.640000  102.400000 ;
      RECT 95.360000  102.520000 95.640000  102.800000 ;
      RECT 96.220000  102.120000 96.500000  102.400000 ;
      RECT 96.220000  102.520000 96.500000  102.800000 ;
      RECT 97.080000  102.120000 97.360000  102.400000 ;
      RECT 97.080000  102.520000 97.360000  102.800000 ;
  END
END sky130_fd_pr__rf_aura_lvs_drc
END LIBRARY
