* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0








.subckt sky130_fd_pr__rf_aura_drc_flag_check B_P NWELL VGND
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_1/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_1/SOURCE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_1/GATE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_1/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_1/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_1/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_2 sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_2/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_2/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_2/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_0 sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_0/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_0/GATE sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_0/SOURCE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_1 sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_1/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_2/GATE sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_1/SOURCE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_3 sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_3/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_3/GATE sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_3/SOURCE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_0 sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_0/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_0/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_1/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_2 sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_2/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_2/GATE sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_2/SOURCE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_1 sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_1/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_1/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_1/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_1/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_4/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_1/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_2 sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_2/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_3/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_2/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_3 sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_3/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_3/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_3/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_2 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_2/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_2/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_2/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_3 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_3/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_2/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_3/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_1 sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_1/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_1/SOURCE sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_3/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_0 sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_0/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_2/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_0/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_4 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_4/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_4/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_4/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_2 sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_2/DRAIN
+ sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_2/SOURCE sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_2/GATE
+ B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_5 sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_5/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_5/GATE sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_5/SOURCE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_0/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_0/SOURCE sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_1/GATE
+ SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15
.ends
