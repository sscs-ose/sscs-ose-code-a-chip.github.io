# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p25 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  4.270000 BY  3.540000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.895000 4.340000 2.535000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.650000 ;
    PORT
      LAYER li1 ;
        RECT 1.240000 0.000000 3.170000 0.695000 ;
        RECT 1.240000 2.845000 3.170000 3.540000 ;
      LAYER mcon ;
        RECT 1.400000 0.095000 3.010000 0.625000 ;
        RECT 1.400000 2.915000 3.010000 3.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.320000 0.000000 3.090000 0.685000 ;
        RECT 1.320000 2.855000 3.090000 3.540000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.005000 4.340000 1.645000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.072500 ;
    ANTENNAGATEAREA  0.247500 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.005000 0.500000 2.535000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.910000 1.005000 4.205000 2.535000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 0.800000 2.615000 ;
      RECT 0.600000 0.485000 0.930000 0.815000 ;
      RECT 0.600000 0.815000 0.800000 0.925000 ;
      RECT 0.600000 2.615000 0.800000 2.725000 ;
      RECT 0.600000 2.725000 0.930000 3.055000 ;
      RECT 1.060000 0.925000 1.230000 2.615000 ;
      RECT 1.590000 0.925000 1.760000 2.615000 ;
      RECT 2.120000 0.925000 2.290000 2.615000 ;
      RECT 2.650000 0.925000 2.820000 2.615000 ;
      RECT 3.180000 0.925000 3.350000 2.615000 ;
      RECT 3.480000 0.485000 3.810000 0.815000 ;
      RECT 3.480000 2.725000 3.810000 3.055000 ;
      RECT 3.610000 0.815000 3.810000 0.925000 ;
      RECT 3.610000 0.925000 4.205000 2.615000 ;
      RECT 3.610000 2.615000 3.810000 2.725000 ;
    LAYER mcon ;
      RECT 0.300000 1.145000 0.470000 1.315000 ;
      RECT 0.300000 1.505000 0.470000 1.675000 ;
      RECT 0.300000 1.865000 0.470000 2.035000 ;
      RECT 0.300000 2.225000 0.470000 2.395000 ;
      RECT 1.060000 1.145000 1.230000 1.315000 ;
      RECT 1.060000 1.505000 1.230000 1.675000 ;
      RECT 1.060000 1.865000 1.230000 2.035000 ;
      RECT 1.060000 2.225000 1.230000 2.395000 ;
      RECT 1.590000 1.145000 1.760000 1.315000 ;
      RECT 1.590000 1.505000 1.760000 1.675000 ;
      RECT 1.590000 1.865000 1.760000 2.035000 ;
      RECT 1.590000 2.225000 1.760000 2.395000 ;
      RECT 2.120000 1.145000 2.290000 1.315000 ;
      RECT 2.120000 1.505000 2.290000 1.675000 ;
      RECT 2.120000 1.865000 2.290000 2.035000 ;
      RECT 2.120000 2.225000 2.290000 2.395000 ;
      RECT 2.650000 1.145000 2.820000 1.315000 ;
      RECT 2.650000 1.505000 2.820000 1.675000 ;
      RECT 2.650000 1.865000 2.820000 2.035000 ;
      RECT 2.650000 2.225000 2.820000 2.395000 ;
      RECT 3.180000 1.145000 3.350000 1.315000 ;
      RECT 3.180000 1.505000 3.350000 1.675000 ;
      RECT 3.180000 1.865000 3.350000 2.035000 ;
      RECT 3.180000 2.225000 3.350000 2.395000 ;
      RECT 3.940000 1.145000 4.110000 1.315000 ;
      RECT 3.940000 1.505000 4.110000 1.675000 ;
      RECT 3.940000 1.865000 4.110000 2.035000 ;
      RECT 3.940000 2.225000 4.110000 2.395000 ;
    LAYER met1 ;
      RECT 1.015000 1.005000 1.275000 2.535000 ;
      RECT 1.545000 1.005000 1.805000 2.535000 ;
      RECT 2.075000 1.005000 2.335000 2.535000 ;
      RECT 2.605000 1.005000 2.865000 2.535000 ;
      RECT 3.135000 1.005000 3.395000 2.535000 ;
    LAYER via ;
      RECT 1.015000 1.035000 1.275000 1.295000 ;
      RECT 1.015000 1.355000 1.275000 1.615000 ;
      RECT 1.545000 1.925000 1.805000 2.185000 ;
      RECT 1.545000 2.245000 1.805000 2.505000 ;
      RECT 2.075000 1.035000 2.335000 1.295000 ;
      RECT 2.075000 1.355000 2.335000 1.615000 ;
      RECT 2.605000 1.925000 2.865000 2.185000 ;
      RECT 2.605000 2.245000 2.865000 2.505000 ;
      RECT 3.135000 1.035000 3.395000 1.295000 ;
      RECT 3.135000 1.355000 3.395000 1.615000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p25
END LIBRARY
