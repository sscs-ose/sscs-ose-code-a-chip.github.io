# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_aura_drc_flag_check
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_aura_drc_flag_check ;
  ORIGIN  0.000000  213.9700 ;
  SIZE  1555.530 BY  412.1700 ;
  PIN B_P
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 -205.320000 11.985000 -202.345000 ;
    END
  END B_P
  PIN NWELL
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 8.650000 11.985000 11.625000 ;
    END
  END NWELL
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 60.140000 90.690000 62.950000 93.665000 ;
    END
  END VGND
  OBS
    LAYER li1 ;
      RECT  64.430000  103.905000  64.600000  104.235000 ;
      RECT  64.610000  104.405000  65.280000  104.735000 ;
      RECT  64.860000  103.905000  65.030000  104.235000 ;
      RECT  65.290000  103.905000  65.460000  104.235000 ;
      RECT  65.930000  103.905000  66.100000  104.235000 ;
      RECT  66.110000  104.405000  66.780000  104.735000 ;
      RECT  66.360000  103.905000  66.530000  104.235000 ;
      RECT  66.790000  103.905000  66.960000  104.235000 ;
      RECT  68.460000 -125.255000  68.630000 -124.565000 ;
      RECT  68.640000 -124.335000  69.310000 -123.995000 ;
      RECT  68.890000 -125.255000  69.060000 -124.565000 ;
      RECT  69.320000 -125.255000  69.490000 -124.565000 ;
      RECT  69.960000 -125.255000  70.130000 -124.565000 ;
      RECT  70.140000 -124.335000  70.810000 -123.995000 ;
      RECT  70.390000 -125.255000  70.560000 -124.565000 ;
      RECT  70.820000 -125.255000  70.990000 -124.565000 ;
      RECT  72.455000  101.200000  72.625000  104.050000 ;
      RECT  72.885000  101.200000  73.055000  104.050000 ;
      RECT  72.905000  100.640000  75.615000  100.970000 ;
      RECT  73.315000  101.200000  73.485000  104.050000 ;
      RECT  73.745000  101.200000  73.915000  104.050000 ;
      RECT  74.175000  101.200000  74.345000  104.050000 ;
      RECT  74.605000  101.200000  74.775000  104.050000 ;
      RECT  75.035000  101.200000  75.205000  104.050000 ;
      RECT  75.465000  101.200000  75.635000  104.050000 ;
      RECT  75.895000  101.200000  76.065000  104.050000 ;
      RECT  76.535000  101.200000  76.705000  104.050000 ;
      RECT  76.630000 -125.330000  76.800000 -120.340000 ;
      RECT  76.810000 -120.170000  77.480000 -119.840000 ;
      RECT  76.965000  101.200000  77.135000  104.050000 ;
      RECT  76.985000  100.640000  79.695000  100.970000 ;
      RECT  77.060000 -125.330000  77.230000 -120.340000 ;
      RECT  77.395000  101.200000  77.565000  104.050000 ;
      RECT  77.490000 -125.330000  77.660000 -120.340000 ;
      RECT  77.825000  101.200000  77.995000  104.050000 ;
      RECT  78.100000 -125.330000  78.270000 -120.340000 ;
      RECT  78.255000  101.200000  78.425000  104.050000 ;
      RECT  78.280000 -120.170000  78.950000 -119.840000 ;
      RECT  78.530000 -125.330000  78.700000 -120.340000 ;
      RECT  78.685000  101.200000  78.855000  104.050000 ;
      RECT  78.960000 -125.330000  79.130000 -120.340000 ;
      RECT  79.115000  101.200000  79.285000  104.050000 ;
      RECT  79.545000  101.200000  79.715000  104.050000 ;
      RECT  79.975000  101.200000  80.145000  104.050000 ;
      RECT  99.085000  102.355000  99.255000  102.685000 ;
      RECT  99.265000  102.855000  99.935000  103.185000 ;
      RECT  99.515000  102.355000  99.685000  102.685000 ;
      RECT  99.945000  102.355000 100.115000  102.685000 ;
      RECT 100.495000  102.355000 100.665000  102.685000 ;
      RECT 100.495000  103.355000 100.665000  103.685000 ;
      RECT 100.675000  102.855000 101.345000  103.185000 ;
      RECT 100.925000  102.355000 101.095000  102.685000 ;
      RECT 100.925000  103.355000 101.095000  103.685000 ;
      RECT 100.930000 -125.255000 101.100000 -124.565000 ;
      RECT 100.930000 -123.755000 101.100000 -123.065000 ;
      RECT 101.110000 -124.335000 101.780000 -123.985000 ;
      RECT 101.355000  102.355000 101.525000  102.685000 ;
      RECT 101.355000  103.355000 101.525000  103.685000 ;
      RECT 101.360000 -125.255000 101.530000 -124.565000 ;
      RECT 101.360000 -123.755000 101.530000 -123.065000 ;
      RECT 101.790000 -125.255000 101.960000 -124.565000 ;
      RECT 101.790000 -123.755000 101.960000 -123.065000 ;
      RECT 104.960000  102.355000 105.130000  103.045000 ;
      RECT 104.960000  103.835000 105.130000  104.525000 ;
      RECT 105.230000  103.275000 106.580000  103.605000 ;
      RECT 105.390000  102.355000 105.560000  103.045000 ;
      RECT 105.390000  103.835000 105.560000  104.525000 ;
      RECT 105.820000  102.355000 105.990000  103.045000 ;
      RECT 105.820000  103.835000 105.990000  104.525000 ;
      RECT 106.250000  102.355000 106.420000  103.045000 ;
      RECT 106.250000  103.835000 106.420000  104.525000 ;
      RECT 106.680000  102.355000 106.850000  103.045000 ;
      RECT 106.680000  103.835000 106.850000  104.525000 ;
      RECT 107.745000 -125.255000 107.915000 -123.725000 ;
      RECT 107.745000 -122.915000 107.915000 -121.385000 ;
      RECT 108.015000 -123.495000 109.365000 -123.145000 ;
      RECT 108.175000 -125.255000 108.345000 -123.725000 ;
      RECT 108.175000 -122.915000 108.345000 -121.385000 ;
      RECT 108.605000 -125.255000 108.775000 -123.725000 ;
      RECT 108.605000 -122.915000 108.775000 -121.385000 ;
      RECT 109.035000 -125.255000 109.205000 -123.725000 ;
      RECT 109.035000 -122.915000 109.205000 -121.385000 ;
      RECT 109.465000 -125.255000 109.635000 -123.725000 ;
      RECT 109.465000 -122.915000 109.635000 -121.385000 ;
      RECT 109.985000 -125.255000 110.155000 -123.725000 ;
      RECT 110.255000 -123.495000 111.605000 -123.155000 ;
      RECT 110.415000 -125.255000 110.585000 -123.725000 ;
      RECT 110.845000 -125.255000 111.015000 -123.725000 ;
      RECT 111.275000 -125.255000 111.445000 -123.725000 ;
      RECT 111.705000 -125.255000 111.875000 -123.725000 ;
      RECT 113.205000  103.490000 113.375000  106.340000 ;
      RECT 113.635000  103.490000 113.805000  106.340000 ;
      RECT 113.655000  102.930000 116.365000  103.260000 ;
      RECT 114.065000  103.490000 114.235000  106.340000 ;
      RECT 114.495000  102.430000 114.665000  102.760000 ;
      RECT 114.495000  103.490000 114.665000  106.340000 ;
      RECT 114.925000  102.430000 115.095000  102.760000 ;
      RECT 114.925000  103.490000 115.095000  106.340000 ;
      RECT 115.355000  102.430000 115.525000  102.760000 ;
      RECT 115.355000  103.490000 115.525000  106.340000 ;
      RECT 115.785000  103.490000 115.955000  106.340000 ;
      RECT 116.215000  103.490000 116.385000  106.340000 ;
      RECT 116.645000  103.490000 116.815000  106.340000 ;
      RECT 116.855000 -122.915000 117.025000 -121.385000 ;
      RECT 117.125000 -123.485000 118.475000 -123.145000 ;
      RECT 117.285000 -128.645000 117.455000 -123.655000 ;
      RECT 117.285000 -122.915000 117.455000 -121.385000 ;
      RECT 117.715000 -128.645000 117.885000 -123.655000 ;
      RECT 117.715000 -122.915000 117.885000 -121.385000 ;
      RECT 118.145000 -128.645000 118.315000 -123.655000 ;
      RECT 118.145000 -122.915000 118.315000 -121.385000 ;
      RECT 118.575000 -122.915000 118.745000 -121.385000 ;
    LAYER mcon ;
      RECT  64.430000  103.985000  64.600000  104.155000 ;
      RECT  64.680000  104.485000  64.850000  104.655000 ;
      RECT  64.860000  103.985000  65.030000  104.155000 ;
      RECT  65.040000  104.485000  65.210000  104.655000 ;
      RECT  65.290000  103.985000  65.460000  104.155000 ;
      RECT  65.930000  103.985000  66.100000  104.155000 ;
      RECT  66.180000  104.485000  66.350000  104.655000 ;
      RECT  66.360000  103.985000  66.530000  104.155000 ;
      RECT  66.540000  104.485000  66.710000  104.655000 ;
      RECT  66.790000  103.985000  66.960000  104.155000 ;
      RECT  68.460000 -125.175000  68.630000 -125.005000 ;
      RECT  68.460000 -124.815000  68.630000 -124.645000 ;
      RECT  68.710000 -124.245000  68.880000 -124.075000 ;
      RECT  68.890000 -125.175000  69.060000 -125.005000 ;
      RECT  68.890000 -124.815000  69.060000 -124.645000 ;
      RECT  69.070000 -124.245000  69.240000 -124.075000 ;
      RECT  69.320000 -125.175000  69.490000 -125.005000 ;
      RECT  69.320000 -124.815000  69.490000 -124.645000 ;
      RECT  69.960000 -125.175000  70.130000 -125.005000 ;
      RECT  69.960000 -124.815000  70.130000 -124.645000 ;
      RECT  70.210000 -124.245000  70.380000 -124.075000 ;
      RECT  70.390000 -125.175000  70.560000 -125.005000 ;
      RECT  70.390000 -124.815000  70.560000 -124.645000 ;
      RECT  70.570000 -124.245000  70.740000 -124.075000 ;
      RECT  70.820000 -125.175000  70.990000 -125.005000 ;
      RECT  70.820000 -124.815000  70.990000 -124.645000 ;
      RECT  72.455000  101.280000  72.625000  101.450000 ;
      RECT  72.455000  101.640000  72.625000  101.810000 ;
      RECT  72.455000  102.000000  72.625000  102.170000 ;
      RECT  72.455000  102.360000  72.625000  102.530000 ;
      RECT  72.455000  102.720000  72.625000  102.890000 ;
      RECT  72.455000  103.080000  72.625000  103.250000 ;
      RECT  72.455000  103.440000  72.625000  103.610000 ;
      RECT  72.455000  103.800000  72.625000  103.970000 ;
      RECT  72.885000  101.280000  73.055000  101.450000 ;
      RECT  72.885000  101.640000  73.055000  101.810000 ;
      RECT  72.885000  102.000000  73.055000  102.170000 ;
      RECT  72.885000  102.360000  73.055000  102.530000 ;
      RECT  72.885000  102.720000  73.055000  102.890000 ;
      RECT  72.885000  103.080000  73.055000  103.250000 ;
      RECT  72.885000  103.440000  73.055000  103.610000 ;
      RECT  72.885000  103.800000  73.055000  103.970000 ;
      RECT  72.915000  100.720000  73.085000  100.890000 ;
      RECT  73.275000  100.720000  73.445000  100.890000 ;
      RECT  73.315000  101.280000  73.485000  101.450000 ;
      RECT  73.315000  101.640000  73.485000  101.810000 ;
      RECT  73.315000  102.000000  73.485000  102.170000 ;
      RECT  73.315000  102.360000  73.485000  102.530000 ;
      RECT  73.315000  102.720000  73.485000  102.890000 ;
      RECT  73.315000  103.080000  73.485000  103.250000 ;
      RECT  73.315000  103.440000  73.485000  103.610000 ;
      RECT  73.315000  103.800000  73.485000  103.970000 ;
      RECT  73.635000  100.720000  73.805000  100.890000 ;
      RECT  73.745000  101.280000  73.915000  101.450000 ;
      RECT  73.745000  101.640000  73.915000  101.810000 ;
      RECT  73.745000  102.000000  73.915000  102.170000 ;
      RECT  73.745000  102.360000  73.915000  102.530000 ;
      RECT  73.745000  102.720000  73.915000  102.890000 ;
      RECT  73.745000  103.080000  73.915000  103.250000 ;
      RECT  73.745000  103.440000  73.915000  103.610000 ;
      RECT  73.745000  103.800000  73.915000  103.970000 ;
      RECT  73.995000  100.720000  74.165000  100.890000 ;
      RECT  74.175000  101.280000  74.345000  101.450000 ;
      RECT  74.175000  101.640000  74.345000  101.810000 ;
      RECT  74.175000  102.000000  74.345000  102.170000 ;
      RECT  74.175000  102.360000  74.345000  102.530000 ;
      RECT  74.175000  102.720000  74.345000  102.890000 ;
      RECT  74.175000  103.080000  74.345000  103.250000 ;
      RECT  74.175000  103.440000  74.345000  103.610000 ;
      RECT  74.175000  103.800000  74.345000  103.970000 ;
      RECT  74.355000  100.720000  74.525000  100.890000 ;
      RECT  74.605000  101.280000  74.775000  101.450000 ;
      RECT  74.605000  101.640000  74.775000  101.810000 ;
      RECT  74.605000  102.000000  74.775000  102.170000 ;
      RECT  74.605000  102.360000  74.775000  102.530000 ;
      RECT  74.605000  102.720000  74.775000  102.890000 ;
      RECT  74.605000  103.080000  74.775000  103.250000 ;
      RECT  74.605000  103.440000  74.775000  103.610000 ;
      RECT  74.605000  103.800000  74.775000  103.970000 ;
      RECT  74.715000  100.720000  74.885000  100.890000 ;
      RECT  75.035000  101.280000  75.205000  101.450000 ;
      RECT  75.035000  101.640000  75.205000  101.810000 ;
      RECT  75.035000  102.000000  75.205000  102.170000 ;
      RECT  75.035000  102.360000  75.205000  102.530000 ;
      RECT  75.035000  102.720000  75.205000  102.890000 ;
      RECT  75.035000  103.080000  75.205000  103.250000 ;
      RECT  75.035000  103.440000  75.205000  103.610000 ;
      RECT  75.035000  103.800000  75.205000  103.970000 ;
      RECT  75.075000  100.720000  75.245000  100.890000 ;
      RECT  75.435000  100.720000  75.605000  100.890000 ;
      RECT  75.465000  101.280000  75.635000  101.450000 ;
      RECT  75.465000  101.640000  75.635000  101.810000 ;
      RECT  75.465000  102.000000  75.635000  102.170000 ;
      RECT  75.465000  102.360000  75.635000  102.530000 ;
      RECT  75.465000  102.720000  75.635000  102.890000 ;
      RECT  75.465000  103.080000  75.635000  103.250000 ;
      RECT  75.465000  103.440000  75.635000  103.610000 ;
      RECT  75.465000  103.800000  75.635000  103.970000 ;
      RECT  75.895000  101.280000  76.065000  101.450000 ;
      RECT  75.895000  101.640000  76.065000  101.810000 ;
      RECT  75.895000  102.000000  76.065000  102.170000 ;
      RECT  75.895000  102.360000  76.065000  102.530000 ;
      RECT  75.895000  102.720000  76.065000  102.890000 ;
      RECT  75.895000  103.080000  76.065000  103.250000 ;
      RECT  75.895000  103.440000  76.065000  103.610000 ;
      RECT  75.895000  103.800000  76.065000  103.970000 ;
      RECT  76.535000  101.280000  76.705000  101.450000 ;
      RECT  76.535000  101.640000  76.705000  101.810000 ;
      RECT  76.535000  102.000000  76.705000  102.170000 ;
      RECT  76.535000  102.360000  76.705000  102.530000 ;
      RECT  76.535000  102.720000  76.705000  102.890000 ;
      RECT  76.535000  103.080000  76.705000  103.250000 ;
      RECT  76.535000  103.440000  76.705000  103.610000 ;
      RECT  76.535000  103.800000  76.705000  103.970000 ;
      RECT  76.630000 -125.075000  76.800000 -124.905000 ;
      RECT  76.630000 -124.715000  76.800000 -124.545000 ;
      RECT  76.630000 -124.355000  76.800000 -124.185000 ;
      RECT  76.630000 -123.995000  76.800000 -123.825000 ;
      RECT  76.630000 -123.635000  76.800000 -123.465000 ;
      RECT  76.630000 -123.275000  76.800000 -123.105000 ;
      RECT  76.630000 -122.915000  76.800000 -122.745000 ;
      RECT  76.630000 -122.555000  76.800000 -122.385000 ;
      RECT  76.630000 -122.195000  76.800000 -122.025000 ;
      RECT  76.630000 -121.835000  76.800000 -121.665000 ;
      RECT  76.630000 -121.475000  76.800000 -121.305000 ;
      RECT  76.630000 -121.115000  76.800000 -120.945000 ;
      RECT  76.630000 -120.755000  76.800000 -120.585000 ;
      RECT  76.880000 -120.090000  77.050000 -119.920000 ;
      RECT  76.965000  101.280000  77.135000  101.450000 ;
      RECT  76.965000  101.640000  77.135000  101.810000 ;
      RECT  76.965000  102.000000  77.135000  102.170000 ;
      RECT  76.965000  102.360000  77.135000  102.530000 ;
      RECT  76.965000  102.720000  77.135000  102.890000 ;
      RECT  76.965000  103.080000  77.135000  103.250000 ;
      RECT  76.965000  103.440000  77.135000  103.610000 ;
      RECT  76.965000  103.800000  77.135000  103.970000 ;
      RECT  76.995000  100.720000  77.165000  100.890000 ;
      RECT  77.060000 -125.075000  77.230000 -124.905000 ;
      RECT  77.060000 -124.715000  77.230000 -124.545000 ;
      RECT  77.060000 -124.355000  77.230000 -124.185000 ;
      RECT  77.060000 -123.995000  77.230000 -123.825000 ;
      RECT  77.060000 -123.635000  77.230000 -123.465000 ;
      RECT  77.060000 -123.275000  77.230000 -123.105000 ;
      RECT  77.060000 -122.915000  77.230000 -122.745000 ;
      RECT  77.060000 -122.555000  77.230000 -122.385000 ;
      RECT  77.060000 -122.195000  77.230000 -122.025000 ;
      RECT  77.060000 -121.835000  77.230000 -121.665000 ;
      RECT  77.060000 -121.475000  77.230000 -121.305000 ;
      RECT  77.060000 -121.115000  77.230000 -120.945000 ;
      RECT  77.060000 -120.755000  77.230000 -120.585000 ;
      RECT  77.240000 -120.090000  77.410000 -119.920000 ;
      RECT  77.355000  100.720000  77.525000  100.890000 ;
      RECT  77.395000  101.280000  77.565000  101.450000 ;
      RECT  77.395000  101.640000  77.565000  101.810000 ;
      RECT  77.395000  102.000000  77.565000  102.170000 ;
      RECT  77.395000  102.360000  77.565000  102.530000 ;
      RECT  77.395000  102.720000  77.565000  102.890000 ;
      RECT  77.395000  103.080000  77.565000  103.250000 ;
      RECT  77.395000  103.440000  77.565000  103.610000 ;
      RECT  77.395000  103.800000  77.565000  103.970000 ;
      RECT  77.490000 -125.075000  77.660000 -124.905000 ;
      RECT  77.490000 -124.715000  77.660000 -124.545000 ;
      RECT  77.490000 -124.355000  77.660000 -124.185000 ;
      RECT  77.490000 -123.995000  77.660000 -123.825000 ;
      RECT  77.490000 -123.635000  77.660000 -123.465000 ;
      RECT  77.490000 -123.275000  77.660000 -123.105000 ;
      RECT  77.490000 -122.915000  77.660000 -122.745000 ;
      RECT  77.490000 -122.555000  77.660000 -122.385000 ;
      RECT  77.490000 -122.195000  77.660000 -122.025000 ;
      RECT  77.490000 -121.835000  77.660000 -121.665000 ;
      RECT  77.490000 -121.475000  77.660000 -121.305000 ;
      RECT  77.490000 -121.115000  77.660000 -120.945000 ;
      RECT  77.490000 -120.755000  77.660000 -120.585000 ;
      RECT  77.715000  100.720000  77.885000  100.890000 ;
      RECT  77.825000  101.280000  77.995000  101.450000 ;
      RECT  77.825000  101.640000  77.995000  101.810000 ;
      RECT  77.825000  102.000000  77.995000  102.170000 ;
      RECT  77.825000  102.360000  77.995000  102.530000 ;
      RECT  77.825000  102.720000  77.995000  102.890000 ;
      RECT  77.825000  103.080000  77.995000  103.250000 ;
      RECT  77.825000  103.440000  77.995000  103.610000 ;
      RECT  77.825000  103.800000  77.995000  103.970000 ;
      RECT  78.075000  100.720000  78.245000  100.890000 ;
      RECT  78.100000 -125.075000  78.270000 -124.905000 ;
      RECT  78.100000 -124.715000  78.270000 -124.545000 ;
      RECT  78.100000 -124.355000  78.270000 -124.185000 ;
      RECT  78.100000 -123.995000  78.270000 -123.825000 ;
      RECT  78.100000 -123.635000  78.270000 -123.465000 ;
      RECT  78.100000 -123.275000  78.270000 -123.105000 ;
      RECT  78.100000 -122.915000  78.270000 -122.745000 ;
      RECT  78.100000 -122.555000  78.270000 -122.385000 ;
      RECT  78.100000 -122.195000  78.270000 -122.025000 ;
      RECT  78.100000 -121.835000  78.270000 -121.665000 ;
      RECT  78.100000 -121.475000  78.270000 -121.305000 ;
      RECT  78.100000 -121.115000  78.270000 -120.945000 ;
      RECT  78.100000 -120.755000  78.270000 -120.585000 ;
      RECT  78.255000  101.280000  78.425000  101.450000 ;
      RECT  78.255000  101.640000  78.425000  101.810000 ;
      RECT  78.255000  102.000000  78.425000  102.170000 ;
      RECT  78.255000  102.360000  78.425000  102.530000 ;
      RECT  78.255000  102.720000  78.425000  102.890000 ;
      RECT  78.255000  103.080000  78.425000  103.250000 ;
      RECT  78.255000  103.440000  78.425000  103.610000 ;
      RECT  78.255000  103.800000  78.425000  103.970000 ;
      RECT  78.350000 -120.090000  78.520000 -119.920000 ;
      RECT  78.435000  100.720000  78.605000  100.890000 ;
      RECT  78.530000 -125.075000  78.700000 -124.905000 ;
      RECT  78.530000 -124.715000  78.700000 -124.545000 ;
      RECT  78.530000 -124.355000  78.700000 -124.185000 ;
      RECT  78.530000 -123.995000  78.700000 -123.825000 ;
      RECT  78.530000 -123.635000  78.700000 -123.465000 ;
      RECT  78.530000 -123.275000  78.700000 -123.105000 ;
      RECT  78.530000 -122.915000  78.700000 -122.745000 ;
      RECT  78.530000 -122.555000  78.700000 -122.385000 ;
      RECT  78.530000 -122.195000  78.700000 -122.025000 ;
      RECT  78.530000 -121.835000  78.700000 -121.665000 ;
      RECT  78.530000 -121.475000  78.700000 -121.305000 ;
      RECT  78.530000 -121.115000  78.700000 -120.945000 ;
      RECT  78.530000 -120.755000  78.700000 -120.585000 ;
      RECT  78.685000  101.280000  78.855000  101.450000 ;
      RECT  78.685000  101.640000  78.855000  101.810000 ;
      RECT  78.685000  102.000000  78.855000  102.170000 ;
      RECT  78.685000  102.360000  78.855000  102.530000 ;
      RECT  78.685000  102.720000  78.855000  102.890000 ;
      RECT  78.685000  103.080000  78.855000  103.250000 ;
      RECT  78.685000  103.440000  78.855000  103.610000 ;
      RECT  78.685000  103.800000  78.855000  103.970000 ;
      RECT  78.710000 -120.090000  78.880000 -119.920000 ;
      RECT  78.795000  100.720000  78.965000  100.890000 ;
      RECT  78.960000 -125.075000  79.130000 -124.905000 ;
      RECT  78.960000 -124.715000  79.130000 -124.545000 ;
      RECT  78.960000 -124.355000  79.130000 -124.185000 ;
      RECT  78.960000 -123.995000  79.130000 -123.825000 ;
      RECT  78.960000 -123.635000  79.130000 -123.465000 ;
      RECT  78.960000 -123.275000  79.130000 -123.105000 ;
      RECT  78.960000 -122.915000  79.130000 -122.745000 ;
      RECT  78.960000 -122.555000  79.130000 -122.385000 ;
      RECT  78.960000 -122.195000  79.130000 -122.025000 ;
      RECT  78.960000 -121.835000  79.130000 -121.665000 ;
      RECT  78.960000 -121.475000  79.130000 -121.305000 ;
      RECT  78.960000 -121.115000  79.130000 -120.945000 ;
      RECT  78.960000 -120.755000  79.130000 -120.585000 ;
      RECT  79.115000  101.280000  79.285000  101.450000 ;
      RECT  79.115000  101.640000  79.285000  101.810000 ;
      RECT  79.115000  102.000000  79.285000  102.170000 ;
      RECT  79.115000  102.360000  79.285000  102.530000 ;
      RECT  79.115000  102.720000  79.285000  102.890000 ;
      RECT  79.115000  103.080000  79.285000  103.250000 ;
      RECT  79.115000  103.440000  79.285000  103.610000 ;
      RECT  79.115000  103.800000  79.285000  103.970000 ;
      RECT  79.155000  100.720000  79.325000  100.890000 ;
      RECT  79.515000  100.720000  79.685000  100.890000 ;
      RECT  79.545000  101.280000  79.715000  101.450000 ;
      RECT  79.545000  101.640000  79.715000  101.810000 ;
      RECT  79.545000  102.000000  79.715000  102.170000 ;
      RECT  79.545000  102.360000  79.715000  102.530000 ;
      RECT  79.545000  102.720000  79.715000  102.890000 ;
      RECT  79.545000  103.080000  79.715000  103.250000 ;
      RECT  79.545000  103.440000  79.715000  103.610000 ;
      RECT  79.545000  103.800000  79.715000  103.970000 ;
      RECT  79.975000  101.280000  80.145000  101.450000 ;
      RECT  79.975000  101.640000  80.145000  101.810000 ;
      RECT  79.975000  102.000000  80.145000  102.170000 ;
      RECT  79.975000  102.360000  80.145000  102.530000 ;
      RECT  79.975000  102.720000  80.145000  102.890000 ;
      RECT  79.975000  103.080000  80.145000  103.250000 ;
      RECT  79.975000  103.440000  80.145000  103.610000 ;
      RECT  79.975000  103.800000  80.145000  103.970000 ;
      RECT  99.085000  102.435000  99.255000  102.605000 ;
      RECT  99.335000  102.935000  99.505000  103.105000 ;
      RECT  99.515000  102.435000  99.685000  102.605000 ;
      RECT  99.695000  102.935000  99.865000  103.105000 ;
      RECT  99.945000  102.435000 100.115000  102.605000 ;
      RECT 100.495000  102.435000 100.665000  102.605000 ;
      RECT 100.495000  103.435000 100.665000  103.605000 ;
      RECT 100.745000  102.935000 100.915000  103.105000 ;
      RECT 100.925000  102.435000 101.095000  102.605000 ;
      RECT 100.925000  103.435000 101.095000  103.605000 ;
      RECT 100.930000 -125.175000 101.100000 -125.005000 ;
      RECT 100.930000 -124.815000 101.100000 -124.645000 ;
      RECT 100.930000 -123.675000 101.100000 -123.505000 ;
      RECT 100.930000 -123.315000 101.100000 -123.145000 ;
      RECT 101.105000  102.935000 101.275000  103.105000 ;
      RECT 101.180000 -124.245000 101.350000 -124.075000 ;
      RECT 101.355000  102.435000 101.525000  102.605000 ;
      RECT 101.355000  103.435000 101.525000  103.605000 ;
      RECT 101.360000 -125.175000 101.530000 -125.005000 ;
      RECT 101.360000 -124.815000 101.530000 -124.645000 ;
      RECT 101.360000 -123.675000 101.530000 -123.505000 ;
      RECT 101.360000 -123.315000 101.530000 -123.145000 ;
      RECT 101.540000 -124.245000 101.710000 -124.075000 ;
      RECT 101.790000 -125.175000 101.960000 -125.005000 ;
      RECT 101.790000 -124.815000 101.960000 -124.645000 ;
      RECT 101.790000 -123.675000 101.960000 -123.505000 ;
      RECT 101.790000 -123.315000 101.960000 -123.145000 ;
      RECT 104.960000  102.435000 105.130000  102.605000 ;
      RECT 104.960000  102.795000 105.130000  102.965000 ;
      RECT 104.960000  103.915000 105.130000  104.085000 ;
      RECT 104.960000  104.275000 105.130000  104.445000 ;
      RECT 105.280000  103.355000 105.450000  103.525000 ;
      RECT 105.390000  102.435000 105.560000  102.605000 ;
      RECT 105.390000  102.795000 105.560000  102.965000 ;
      RECT 105.390000  103.915000 105.560000  104.085000 ;
      RECT 105.390000  104.275000 105.560000  104.445000 ;
      RECT 105.640000  103.355000 105.810000  103.525000 ;
      RECT 105.820000  102.435000 105.990000  102.605000 ;
      RECT 105.820000  102.795000 105.990000  102.965000 ;
      RECT 105.820000  103.915000 105.990000  104.085000 ;
      RECT 105.820000  104.275000 105.990000  104.445000 ;
      RECT 106.000000  103.355000 106.170000  103.525000 ;
      RECT 106.250000  102.435000 106.420000  102.605000 ;
      RECT 106.250000  102.795000 106.420000  102.965000 ;
      RECT 106.250000  103.915000 106.420000  104.085000 ;
      RECT 106.250000  104.275000 106.420000  104.445000 ;
      RECT 106.360000  103.355000 106.530000  103.525000 ;
      RECT 106.680000  102.435000 106.850000  102.605000 ;
      RECT 106.680000  102.795000 106.850000  102.965000 ;
      RECT 106.680000  103.915000 106.850000  104.085000 ;
      RECT 106.680000  104.275000 106.850000  104.445000 ;
      RECT 107.745000 -125.115000 107.915000 -124.945000 ;
      RECT 107.745000 -124.755000 107.915000 -124.585000 ;
      RECT 107.745000 -124.395000 107.915000 -124.225000 ;
      RECT 107.745000 -124.035000 107.915000 -123.865000 ;
      RECT 107.745000 -122.775000 107.915000 -122.605000 ;
      RECT 107.745000 -122.415000 107.915000 -122.245000 ;
      RECT 107.745000 -122.055000 107.915000 -121.885000 ;
      RECT 107.745000 -121.695000 107.915000 -121.525000 ;
      RECT 108.065000 -123.405000 108.235000 -123.235000 ;
      RECT 108.175000 -125.115000 108.345000 -124.945000 ;
      RECT 108.175000 -124.755000 108.345000 -124.585000 ;
      RECT 108.175000 -124.395000 108.345000 -124.225000 ;
      RECT 108.175000 -124.035000 108.345000 -123.865000 ;
      RECT 108.175000 -122.775000 108.345000 -122.605000 ;
      RECT 108.175000 -122.415000 108.345000 -122.245000 ;
      RECT 108.175000 -122.055000 108.345000 -121.885000 ;
      RECT 108.175000 -121.695000 108.345000 -121.525000 ;
      RECT 108.425000 -123.405000 108.595000 -123.235000 ;
      RECT 108.605000 -125.115000 108.775000 -124.945000 ;
      RECT 108.605000 -124.755000 108.775000 -124.585000 ;
      RECT 108.605000 -124.395000 108.775000 -124.225000 ;
      RECT 108.605000 -124.035000 108.775000 -123.865000 ;
      RECT 108.605000 -122.775000 108.775000 -122.605000 ;
      RECT 108.605000 -122.415000 108.775000 -122.245000 ;
      RECT 108.605000 -122.055000 108.775000 -121.885000 ;
      RECT 108.605000 -121.695000 108.775000 -121.525000 ;
      RECT 108.785000 -123.405000 108.955000 -123.235000 ;
      RECT 109.035000 -125.115000 109.205000 -124.945000 ;
      RECT 109.035000 -124.755000 109.205000 -124.585000 ;
      RECT 109.035000 -124.395000 109.205000 -124.225000 ;
      RECT 109.035000 -124.035000 109.205000 -123.865000 ;
      RECT 109.035000 -122.775000 109.205000 -122.605000 ;
      RECT 109.035000 -122.415000 109.205000 -122.245000 ;
      RECT 109.035000 -122.055000 109.205000 -121.885000 ;
      RECT 109.035000 -121.695000 109.205000 -121.525000 ;
      RECT 109.145000 -123.405000 109.315000 -123.235000 ;
      RECT 109.465000 -125.115000 109.635000 -124.945000 ;
      RECT 109.465000 -124.755000 109.635000 -124.585000 ;
      RECT 109.465000 -124.395000 109.635000 -124.225000 ;
      RECT 109.465000 -124.035000 109.635000 -123.865000 ;
      RECT 109.465000 -122.775000 109.635000 -122.605000 ;
      RECT 109.465000 -122.415000 109.635000 -122.245000 ;
      RECT 109.465000 -122.055000 109.635000 -121.885000 ;
      RECT 109.465000 -121.695000 109.635000 -121.525000 ;
      RECT 109.985000 -125.115000 110.155000 -124.945000 ;
      RECT 109.985000 -124.755000 110.155000 -124.585000 ;
      RECT 109.985000 -124.395000 110.155000 -124.225000 ;
      RECT 109.985000 -124.035000 110.155000 -123.865000 ;
      RECT 110.305000 -123.405000 110.475000 -123.235000 ;
      RECT 110.415000 -125.115000 110.585000 -124.945000 ;
      RECT 110.415000 -124.755000 110.585000 -124.585000 ;
      RECT 110.415000 -124.395000 110.585000 -124.225000 ;
      RECT 110.415000 -124.035000 110.585000 -123.865000 ;
      RECT 110.665000 -123.405000 110.835000 -123.235000 ;
      RECT 110.845000 -125.115000 111.015000 -124.945000 ;
      RECT 110.845000 -124.755000 111.015000 -124.585000 ;
      RECT 110.845000 -124.395000 111.015000 -124.225000 ;
      RECT 110.845000 -124.035000 111.015000 -123.865000 ;
      RECT 111.025000 -123.405000 111.195000 -123.235000 ;
      RECT 111.275000 -125.115000 111.445000 -124.945000 ;
      RECT 111.275000 -124.755000 111.445000 -124.585000 ;
      RECT 111.275000 -124.395000 111.445000 -124.225000 ;
      RECT 111.275000 -124.035000 111.445000 -123.865000 ;
      RECT 111.385000 -123.405000 111.555000 -123.235000 ;
      RECT 111.705000 -125.115000 111.875000 -124.945000 ;
      RECT 111.705000 -124.755000 111.875000 -124.585000 ;
      RECT 111.705000 -124.395000 111.875000 -124.225000 ;
      RECT 111.705000 -124.035000 111.875000 -123.865000 ;
      RECT 113.205000  103.570000 113.375000  103.740000 ;
      RECT 113.205000  103.930000 113.375000  104.100000 ;
      RECT 113.205000  104.290000 113.375000  104.460000 ;
      RECT 113.205000  104.650000 113.375000  104.820000 ;
      RECT 113.205000  105.010000 113.375000  105.180000 ;
      RECT 113.205000  105.370000 113.375000  105.540000 ;
      RECT 113.205000  105.730000 113.375000  105.900000 ;
      RECT 113.205000  106.090000 113.375000  106.260000 ;
      RECT 113.635000  103.570000 113.805000  103.740000 ;
      RECT 113.635000  103.930000 113.805000  104.100000 ;
      RECT 113.635000  104.290000 113.805000  104.460000 ;
      RECT 113.635000  104.650000 113.805000  104.820000 ;
      RECT 113.635000  105.010000 113.805000  105.180000 ;
      RECT 113.635000  105.370000 113.805000  105.540000 ;
      RECT 113.635000  105.730000 113.805000  105.900000 ;
      RECT 113.635000  106.090000 113.805000  106.260000 ;
      RECT 113.665000  103.010000 113.835000  103.180000 ;
      RECT 114.025000  103.010000 114.195000  103.180000 ;
      RECT 114.065000  103.570000 114.235000  103.740000 ;
      RECT 114.065000  103.930000 114.235000  104.100000 ;
      RECT 114.065000  104.290000 114.235000  104.460000 ;
      RECT 114.065000  104.650000 114.235000  104.820000 ;
      RECT 114.065000  105.010000 114.235000  105.180000 ;
      RECT 114.065000  105.370000 114.235000  105.540000 ;
      RECT 114.065000  105.730000 114.235000  105.900000 ;
      RECT 114.065000  106.090000 114.235000  106.260000 ;
      RECT 114.385000  103.010000 114.555000  103.180000 ;
      RECT 114.495000  102.510000 114.665000  102.680000 ;
      RECT 114.495000  103.570000 114.665000  103.740000 ;
      RECT 114.495000  103.930000 114.665000  104.100000 ;
      RECT 114.495000  104.290000 114.665000  104.460000 ;
      RECT 114.495000  104.650000 114.665000  104.820000 ;
      RECT 114.495000  105.010000 114.665000  105.180000 ;
      RECT 114.495000  105.370000 114.665000  105.540000 ;
      RECT 114.495000  105.730000 114.665000  105.900000 ;
      RECT 114.495000  106.090000 114.665000  106.260000 ;
      RECT 114.745000  103.010000 114.915000  103.180000 ;
      RECT 114.925000  102.510000 115.095000  102.680000 ;
      RECT 114.925000  103.570000 115.095000  103.740000 ;
      RECT 114.925000  103.930000 115.095000  104.100000 ;
      RECT 114.925000  104.290000 115.095000  104.460000 ;
      RECT 114.925000  104.650000 115.095000  104.820000 ;
      RECT 114.925000  105.010000 115.095000  105.180000 ;
      RECT 114.925000  105.370000 115.095000  105.540000 ;
      RECT 114.925000  105.730000 115.095000  105.900000 ;
      RECT 114.925000  106.090000 115.095000  106.260000 ;
      RECT 115.105000  103.010000 115.275000  103.180000 ;
      RECT 115.355000  102.510000 115.525000  102.680000 ;
      RECT 115.355000  103.570000 115.525000  103.740000 ;
      RECT 115.355000  103.930000 115.525000  104.100000 ;
      RECT 115.355000  104.290000 115.525000  104.460000 ;
      RECT 115.355000  104.650000 115.525000  104.820000 ;
      RECT 115.355000  105.010000 115.525000  105.180000 ;
      RECT 115.355000  105.370000 115.525000  105.540000 ;
      RECT 115.355000  105.730000 115.525000  105.900000 ;
      RECT 115.355000  106.090000 115.525000  106.260000 ;
      RECT 115.465000  103.010000 115.635000  103.180000 ;
      RECT 115.785000  103.570000 115.955000  103.740000 ;
      RECT 115.785000  103.930000 115.955000  104.100000 ;
      RECT 115.785000  104.290000 115.955000  104.460000 ;
      RECT 115.785000  104.650000 115.955000  104.820000 ;
      RECT 115.785000  105.010000 115.955000  105.180000 ;
      RECT 115.785000  105.370000 115.955000  105.540000 ;
      RECT 115.785000  105.730000 115.955000  105.900000 ;
      RECT 115.785000  106.090000 115.955000  106.260000 ;
      RECT 115.825000  103.010000 115.995000  103.180000 ;
      RECT 116.185000  103.010000 116.355000  103.180000 ;
      RECT 116.215000  103.570000 116.385000  103.740000 ;
      RECT 116.215000  103.930000 116.385000  104.100000 ;
      RECT 116.215000  104.290000 116.385000  104.460000 ;
      RECT 116.215000  104.650000 116.385000  104.820000 ;
      RECT 116.215000  105.010000 116.385000  105.180000 ;
      RECT 116.215000  105.370000 116.385000  105.540000 ;
      RECT 116.215000  105.730000 116.385000  105.900000 ;
      RECT 116.215000  106.090000 116.385000  106.260000 ;
      RECT 116.645000  103.570000 116.815000  103.740000 ;
      RECT 116.645000  103.930000 116.815000  104.100000 ;
      RECT 116.645000  104.290000 116.815000  104.460000 ;
      RECT 116.645000  104.650000 116.815000  104.820000 ;
      RECT 116.645000  105.010000 116.815000  105.180000 ;
      RECT 116.645000  105.370000 116.815000  105.540000 ;
      RECT 116.645000  105.730000 116.815000  105.900000 ;
      RECT 116.645000  106.090000 116.815000  106.260000 ;
      RECT 116.855000 -122.775000 117.025000 -122.605000 ;
      RECT 116.855000 -122.415000 117.025000 -122.245000 ;
      RECT 116.855000 -122.055000 117.025000 -121.885000 ;
      RECT 116.855000 -121.695000 117.025000 -121.525000 ;
      RECT 117.175000 -123.405000 117.345000 -123.235000 ;
      RECT 117.285000 -128.390000 117.455000 -128.220000 ;
      RECT 117.285000 -128.030000 117.455000 -127.860000 ;
      RECT 117.285000 -127.670000 117.455000 -127.500000 ;
      RECT 117.285000 -127.310000 117.455000 -127.140000 ;
      RECT 117.285000 -126.950000 117.455000 -126.780000 ;
      RECT 117.285000 -126.590000 117.455000 -126.420000 ;
      RECT 117.285000 -126.230000 117.455000 -126.060000 ;
      RECT 117.285000 -125.870000 117.455000 -125.700000 ;
      RECT 117.285000 -125.510000 117.455000 -125.340000 ;
      RECT 117.285000 -125.150000 117.455000 -124.980000 ;
      RECT 117.285000 -124.790000 117.455000 -124.620000 ;
      RECT 117.285000 -124.430000 117.455000 -124.260000 ;
      RECT 117.285000 -124.070000 117.455000 -123.900000 ;
      RECT 117.285000 -122.775000 117.455000 -122.605000 ;
      RECT 117.285000 -122.415000 117.455000 -122.245000 ;
      RECT 117.285000 -122.055000 117.455000 -121.885000 ;
      RECT 117.285000 -121.695000 117.455000 -121.525000 ;
      RECT 117.535000 -123.405000 117.705000 -123.235000 ;
      RECT 117.715000 -128.390000 117.885000 -128.220000 ;
      RECT 117.715000 -128.030000 117.885000 -127.860000 ;
      RECT 117.715000 -127.670000 117.885000 -127.500000 ;
      RECT 117.715000 -127.310000 117.885000 -127.140000 ;
      RECT 117.715000 -126.950000 117.885000 -126.780000 ;
      RECT 117.715000 -126.590000 117.885000 -126.420000 ;
      RECT 117.715000 -126.230000 117.885000 -126.060000 ;
      RECT 117.715000 -125.870000 117.885000 -125.700000 ;
      RECT 117.715000 -125.510000 117.885000 -125.340000 ;
      RECT 117.715000 -125.150000 117.885000 -124.980000 ;
      RECT 117.715000 -124.790000 117.885000 -124.620000 ;
      RECT 117.715000 -124.430000 117.885000 -124.260000 ;
      RECT 117.715000 -124.070000 117.885000 -123.900000 ;
      RECT 117.715000 -122.775000 117.885000 -122.605000 ;
      RECT 117.715000 -122.415000 117.885000 -122.245000 ;
      RECT 117.715000 -122.055000 117.885000 -121.885000 ;
      RECT 117.715000 -121.695000 117.885000 -121.525000 ;
      RECT 117.895000 -123.405000 118.065000 -123.235000 ;
      RECT 118.145000 -128.390000 118.315000 -128.220000 ;
      RECT 118.145000 -128.030000 118.315000 -127.860000 ;
      RECT 118.145000 -127.670000 118.315000 -127.500000 ;
      RECT 118.145000 -127.310000 118.315000 -127.140000 ;
      RECT 118.145000 -126.950000 118.315000 -126.780000 ;
      RECT 118.145000 -126.590000 118.315000 -126.420000 ;
      RECT 118.145000 -126.230000 118.315000 -126.060000 ;
      RECT 118.145000 -125.870000 118.315000 -125.700000 ;
      RECT 118.145000 -125.510000 118.315000 -125.340000 ;
      RECT 118.145000 -125.150000 118.315000 -124.980000 ;
      RECT 118.145000 -124.790000 118.315000 -124.620000 ;
      RECT 118.145000 -124.430000 118.315000 -124.260000 ;
      RECT 118.145000 -124.070000 118.315000 -123.900000 ;
      RECT 118.145000 -122.775000 118.315000 -122.605000 ;
      RECT 118.145000 -122.415000 118.315000 -122.245000 ;
      RECT 118.145000 -122.055000 118.315000 -121.885000 ;
      RECT 118.145000 -121.695000 118.315000 -121.525000 ;
      RECT 118.255000 -123.405000 118.425000 -123.235000 ;
      RECT 118.575000 -122.775000 118.745000 -122.605000 ;
      RECT 118.575000 -122.415000 118.745000 -122.245000 ;
      RECT 118.575000 -122.055000 118.745000 -121.885000 ;
      RECT 118.575000 -121.695000 118.745000 -121.525000 ;
    LAYER met1 ;
      RECT  64.400000  103.205000  65.490000  103.505000 ;
      RECT  64.400000  103.505000  64.630000  104.250000 ;
      RECT  64.620000  104.425000  65.270000  104.715000 ;
      RECT  64.815000  103.905000  65.075000  104.250000 ;
      RECT  65.260000  103.505000  65.490000  104.250000 ;
      RECT  65.900000  103.205000  66.990000  103.505000 ;
      RECT  65.900000  103.505000  66.130000  104.250000 ;
      RECT  66.120000  104.425000  66.770000  104.715000 ;
      RECT  66.315000  103.905000  66.575000  104.250000 ;
      RECT  66.760000  103.505000  66.990000  104.250000 ;
      RECT  68.430000 -125.955000  69.520000 -125.655000 ;
      RECT  68.430000 -125.655000  68.660000 -124.565000 ;
      RECT  68.650000 -124.305000  69.300000 -124.015000 ;
      RECT  68.845000 -125.255000  69.105000 -124.565000 ;
      RECT  69.290000 -125.655000  69.520000 -124.565000 ;
      RECT  69.930000 -125.955000  71.020000 -125.655000 ;
      RECT  69.930000 -125.655000  70.160000 -124.565000 ;
      RECT  70.150000 -124.305000  70.800000 -124.015000 ;
      RECT  70.345000 -125.255000  70.605000 -124.565000 ;
      RECT  70.790000 -125.655000  71.020000 -124.565000 ;
      RECT  72.425000  101.200000  72.655000  104.450000 ;
      RECT  72.425000  104.450000  76.095000  104.750000 ;
      RECT  72.840000  101.200000  73.100000  104.050000 ;
      RECT  72.855000  100.660000  75.665000  100.950000 ;
      RECT  73.285000  101.200000  73.515000  104.450000 ;
      RECT  73.700000  101.200000  73.960000  104.050000 ;
      RECT  74.145000  101.200000  74.375000  104.450000 ;
      RECT  74.560000  101.200000  74.820000  104.050000 ;
      RECT  75.005000  101.200000  75.235000  104.450000 ;
      RECT  75.420000  101.200000  75.680000  104.050000 ;
      RECT  75.865000  101.200000  76.095000  104.450000 ;
      RECT  76.505000  101.200000  76.735000  104.450000 ;
      RECT  76.505000  104.450000  80.175000  104.750000 ;
      RECT  76.600000 -125.995000  77.690000 -125.735000 ;
      RECT  76.600000 -125.735000  76.830000 -120.340000 ;
      RECT  76.820000 -120.150000  77.470000 -119.860000 ;
      RECT  76.920000  101.200000  77.180000  104.050000 ;
      RECT  76.935000  100.660000  79.745000  100.950000 ;
      RECT  77.015000 -125.330000  77.275000 -120.340000 ;
      RECT  77.365000  101.200000  77.595000  104.450000 ;
      RECT  77.460000 -125.735000  77.690000 -120.340000 ;
      RECT  77.780000  101.200000  78.040000  104.050000 ;
      RECT  78.070000 -125.995000  79.160000 -125.735000 ;
      RECT  78.070000 -125.735000  78.300000 -120.340000 ;
      RECT  78.225000  101.200000  78.455000  104.450000 ;
      RECT  78.290000 -120.150000  78.940000 -119.860000 ;
      RECT  78.485000 -125.330000  78.745000 -120.340000 ;
      RECT  78.640000  101.200000  78.900000  104.050000 ;
      RECT  78.930000 -125.735000  79.160000 -120.340000 ;
      RECT  79.085000  101.200000  79.315000  104.450000 ;
      RECT  79.500000  101.200000  79.760000  104.050000 ;
      RECT  79.945000  101.200000  80.175000  104.450000 ;
      RECT  99.055000  101.655000 100.145000  101.955000 ;
      RECT  99.055000  101.955000  99.285000  102.700000 ;
      RECT  99.275000  102.875000  99.925000  103.165000 ;
      RECT  99.470000  102.355000  99.730000  102.700000 ;
      RECT  99.915000  101.955000 100.145000  102.700000 ;
      RECT 100.465000  101.655000 101.555000  101.955000 ;
      RECT 100.465000  101.955000 100.695000  102.700000 ;
      RECT 100.465000  103.340000 100.695000  104.085000 ;
      RECT 100.465000  104.085000 101.555000  104.385000 ;
      RECT 100.685000  102.875000 101.335000  103.165000 ;
      RECT 100.880000  102.355000 101.140000  102.700000 ;
      RECT 100.880000  103.340000 101.140000  103.685000 ;
      RECT 100.900000 -125.955000 101.990000 -125.655000 ;
      RECT 100.900000 -125.655000 101.130000 -124.565000 ;
      RECT 100.900000 -123.755000 101.130000 -122.665000 ;
      RECT 100.900000 -122.665000 101.990000 -122.365000 ;
      RECT 101.120000 -124.305000 101.770000 -124.015000 ;
      RECT 101.315000 -125.255000 101.575000 -124.565000 ;
      RECT 101.315000 -123.755000 101.575000 -123.065000 ;
      RECT 101.325000  101.955000 101.555000  102.700000 ;
      RECT 101.325000  103.340000 101.555000  104.085000 ;
      RECT 101.760000 -125.655000 101.990000 -124.565000 ;
      RECT 101.760000 -123.755000 101.990000 -122.665000 ;
      RECT 104.930000  101.655000 106.880000  101.955000 ;
      RECT 104.930000  101.955000 105.160000  103.045000 ;
      RECT 104.930000  103.835000 105.160000  104.925000 ;
      RECT 104.930000  104.925000 106.880000  105.225000 ;
      RECT 105.220000  103.295000 106.590000  103.585000 ;
      RECT 105.345000  102.355000 105.605000  103.045000 ;
      RECT 105.345000  103.835000 105.605000  104.525000 ;
      RECT 105.790000  101.955000 106.020000  103.045000 ;
      RECT 105.790000  103.835000 106.020000  104.925000 ;
      RECT 106.205000  102.355000 106.465000  103.045000 ;
      RECT 106.205000  103.835000 106.465000  104.525000 ;
      RECT 106.650000  101.955000 106.880000  103.045000 ;
      RECT 106.650000  103.835000 106.880000  104.925000 ;
      RECT 107.715000 -125.955000 109.665000 -125.655000 ;
      RECT 107.715000 -125.655000 107.945000 -123.725000 ;
      RECT 107.715000 -122.915000 107.945000 -120.985000 ;
      RECT 107.715000 -120.985000 109.665000 -120.685000 ;
      RECT 108.005000 -123.465000 109.375000 -123.175000 ;
      RECT 108.130000 -125.255000 108.390000 -123.725000 ;
      RECT 108.130000 -122.915000 108.390000 -121.385000 ;
      RECT 108.575000 -125.655000 108.805000 -123.725000 ;
      RECT 108.575000 -122.915000 108.805000 -120.985000 ;
      RECT 108.990000 -125.255000 109.250000 -123.725000 ;
      RECT 108.990000 -122.915000 109.250000 -121.385000 ;
      RECT 109.435000 -125.655000 109.665000 -123.725000 ;
      RECT 109.435000 -122.915000 109.665000 -120.985000 ;
      RECT 109.955000 -125.955000 111.905000 -125.655000 ;
      RECT 109.955000 -125.655000 110.185000 -123.725000 ;
      RECT 110.245000 -123.465000 111.615000 -123.175000 ;
      RECT 110.370000 -125.255000 110.630000 -123.725000 ;
      RECT 110.815000 -125.655000 111.045000 -123.725000 ;
      RECT 111.230000 -125.255000 111.490000 -123.725000 ;
      RECT 111.675000 -125.655000 111.905000 -123.725000 ;
      RECT 113.175000  103.490000 113.405000  106.740000 ;
      RECT 113.175000  106.740000 116.845000  107.040000 ;
      RECT 113.590000  103.490000 113.850000  106.340000 ;
      RECT 113.605000  102.950000 116.415000  103.240000 ;
      RECT 114.035000  103.490000 114.265000  106.740000 ;
      RECT 114.450000  103.490000 114.710000  106.340000 ;
      RECT 114.465000  101.730000 115.555000  102.030000 ;
      RECT 114.465000  102.030000 114.695000  102.775000 ;
      RECT 114.880000  102.430000 115.140000  102.775000 ;
      RECT 114.895000  103.490000 115.125000  106.740000 ;
      RECT 115.310000  103.490000 115.570000  106.340000 ;
      RECT 115.325000  102.030000 115.555000  102.775000 ;
      RECT 115.755000  103.490000 115.985000  106.740000 ;
      RECT 116.170000  103.490000 116.430000  106.340000 ;
      RECT 116.615000  103.490000 116.845000  106.740000 ;
      RECT 116.825000 -122.915000 117.055000 -120.985000 ;
      RECT 116.825000 -120.985000 118.775000 -120.685000 ;
      RECT 117.115000 -123.465000 118.485000 -123.175000 ;
      RECT 117.240000 -122.915000 117.500000 -121.385000 ;
      RECT 117.255000 -129.310000 118.345000 -129.050000 ;
      RECT 117.255000 -129.050000 117.485000 -123.655000 ;
      RECT 117.670000 -128.645000 117.930000 -123.655000 ;
      RECT 117.685000 -122.915000 117.915000 -120.985000 ;
      RECT 118.100000 -122.915000 118.360000 -121.385000 ;
      RECT 118.115000 -129.050000 118.345000 -123.655000 ;
      RECT 118.545000 -122.915000 118.775000 -120.985000 ;
    LAYER met2 ;
      RECT  64.815000  103.905000  65.075000  104.250000 ;
      RECT  66.315000  103.905000  66.575000  104.250000 ;
      RECT  68.845000 -125.230000  69.105000 -124.590000 ;
      RECT  70.345000 -125.230000  70.605000 -124.590000 ;
      RECT  72.805000  101.170000  73.135000  101.940000 ;
      RECT  73.665000  101.170000  73.995000  101.940000 ;
      RECT  74.525000  101.170000  74.855000  101.940000 ;
      RECT  75.385000  101.170000  75.715000  101.940000 ;
      RECT  76.885000  101.170000  77.215000  101.940000 ;
      RECT  77.015000 -120.990000  77.275000 -120.350000 ;
      RECT  77.745000  101.170000  78.075000  101.940000 ;
      RECT  78.485000 -120.990000  78.745000 -120.350000 ;
      RECT  78.605000  101.170000  78.935000  101.940000 ;
      RECT  79.465000  101.170000  79.795000  101.940000 ;
      RECT  99.470000  102.355000  99.730000  102.700000 ;
      RECT 100.880000  102.355000 101.140000  102.700000 ;
      RECT 100.880000  103.340000 101.140000  103.685000 ;
      RECT 101.315000 -125.230000 101.575000 -124.590000 ;
      RECT 101.315000 -123.730000 101.575000 -123.090000 ;
      RECT 105.310000  102.305000 105.640000  103.075000 ;
      RECT 105.310000  103.805000 105.640000  104.575000 ;
      RECT 106.170000  102.305000 106.500000  103.075000 ;
      RECT 106.170000  103.805000 106.500000  104.575000 ;
      RECT 108.095000 -124.455000 108.425000 -123.685000 ;
      RECT 108.095000 -122.955000 108.425000 -122.185000 ;
      RECT 108.955000 -124.455000 109.285000 -123.685000 ;
      RECT 108.955000 -122.955000 109.285000 -122.185000 ;
      RECT 110.335000 -124.455000 110.665000 -123.685000 ;
      RECT 111.195000 -124.455000 111.525000 -123.685000 ;
      RECT 113.555000  103.460000 113.885000  104.230000 ;
      RECT 114.415000  103.460000 114.745000  104.230000 ;
      RECT 114.880000  102.430000 115.140000  102.775000 ;
      RECT 115.275000  103.460000 115.605000  104.230000 ;
      RECT 116.135000  103.460000 116.465000  104.230000 ;
      RECT 117.205000 -122.955000 117.535000 -122.185000 ;
      RECT 117.670000 -124.305000 117.930000 -123.665000 ;
      RECT 118.065000 -122.955000 118.395000 -122.185000 ;
    LAYER met3 ;
      RECT  72.805000  101.170000  75.715000  101.500000 ;
      RECT  72.805000  101.500000  73.135000  101.940000 ;
      RECT  73.665000  101.500000  73.995000  101.940000 ;
      RECT  74.525000  101.500000  74.855000  101.940000 ;
      RECT  75.385000  101.500000  75.715000  101.940000 ;
      RECT  76.885000  101.170000  79.795000  101.500000 ;
      RECT  76.885000  101.500000  77.215000  101.940000 ;
      RECT  77.745000  101.500000  78.075000  101.940000 ;
      RECT  78.605000  101.500000  78.935000  101.940000 ;
      RECT  79.465000  101.500000  79.795000  101.940000 ;
      RECT 105.310000  102.305000 105.640000  102.745000 ;
      RECT 105.310000  102.745000 106.500000  103.075000 ;
      RECT 105.310000  103.805000 106.500000  104.135000 ;
      RECT 105.310000  104.135000 105.640000  104.575000 ;
      RECT 106.170000  102.305000 106.500000  102.745000 ;
      RECT 106.170000  104.135000 106.500000  104.575000 ;
      RECT 108.095000 -124.455000 108.425000 -124.015000 ;
      RECT 108.095000 -124.015000 109.285000 -123.685000 ;
      RECT 108.095000 -122.955000 109.285000 -122.625000 ;
      RECT 108.095000 -122.625000 108.425000 -122.185000 ;
      RECT 108.955000 -124.455000 109.285000 -124.015000 ;
      RECT 108.955000 -122.625000 109.285000 -122.185000 ;
      RECT 110.335000 -124.455000 110.665000 -124.015000 ;
      RECT 110.335000 -124.015000 111.525000 -123.685000 ;
      RECT 111.195000 -124.455000 111.525000 -124.015000 ;
      RECT 113.555000  103.460000 116.465000  103.790000 ;
      RECT 113.555000  103.790000 113.885000  104.230000 ;
      RECT 114.415000  103.790000 114.745000  104.230000 ;
      RECT 115.275000  103.790000 115.605000  104.230000 ;
      RECT 116.135000  103.790000 116.465000  104.230000 ;
      RECT 117.205000 -122.955000 118.395000 -122.625000 ;
      RECT 117.205000 -122.625000 117.535000 -122.185000 ;
      RECT 118.065000 -122.625000 118.395000 -122.185000 ;
    LAYER via ;
      RECT  64.815000  103.960000  65.075000  104.220000 ;
      RECT  66.315000  103.960000  66.575000  104.220000 ;
      RECT  68.845000 -125.200000  69.105000 -124.940000 ;
      RECT  68.845000 -124.880000  69.105000 -124.620000 ;
      RECT  70.345000 -125.200000  70.605000 -124.940000 ;
      RECT  70.345000 -124.880000  70.605000 -124.620000 ;
      RECT  72.840000  101.265000  73.100000  101.525000 ;
      RECT  72.840000  101.585000  73.100000  101.845000 ;
      RECT  73.700000  101.265000  73.960000  101.525000 ;
      RECT  73.700000  101.585000  73.960000  101.845000 ;
      RECT  74.560000  101.265000  74.820000  101.525000 ;
      RECT  74.560000  101.585000  74.820000  101.845000 ;
      RECT  75.420000  101.265000  75.680000  101.525000 ;
      RECT  75.420000  101.585000  75.680000  101.845000 ;
      RECT  76.920000  101.265000  77.180000  101.525000 ;
      RECT  76.920000  101.585000  77.180000  101.845000 ;
      RECT  77.015000 -120.960000  77.275000 -120.700000 ;
      RECT  77.015000 -120.640000  77.275000 -120.380000 ;
      RECT  77.780000  101.265000  78.040000  101.525000 ;
      RECT  77.780000  101.585000  78.040000  101.845000 ;
      RECT  78.485000 -120.960000  78.745000 -120.700000 ;
      RECT  78.485000 -120.640000  78.745000 -120.380000 ;
      RECT  78.640000  101.265000  78.900000  101.525000 ;
      RECT  78.640000  101.585000  78.900000  101.845000 ;
      RECT  79.500000  101.265000  79.760000  101.525000 ;
      RECT  79.500000  101.585000  79.760000  101.845000 ;
      RECT  99.470000  102.410000  99.730000  102.670000 ;
      RECT 100.880000  102.410000 101.140000  102.670000 ;
      RECT 100.880000  103.370000 101.140000  103.630000 ;
      RECT 101.315000 -125.200000 101.575000 -124.940000 ;
      RECT 101.315000 -124.880000 101.575000 -124.620000 ;
      RECT 101.315000 -123.700000 101.575000 -123.440000 ;
      RECT 101.315000 -123.380000 101.575000 -123.120000 ;
      RECT 105.345000  102.395000 105.605000  102.655000 ;
      RECT 105.345000  102.715000 105.605000  102.975000 ;
      RECT 105.345000  103.905000 105.605000  104.165000 ;
      RECT 105.345000  104.225000 105.605000  104.485000 ;
      RECT 106.205000  102.395000 106.465000  102.655000 ;
      RECT 106.205000  102.715000 106.465000  102.975000 ;
      RECT 106.205000  103.905000 106.465000  104.165000 ;
      RECT 106.205000  104.225000 106.465000  104.485000 ;
      RECT 108.130000 -124.360000 108.390000 -124.100000 ;
      RECT 108.130000 -124.040000 108.390000 -123.780000 ;
      RECT 108.130000 -122.860000 108.390000 -122.600000 ;
      RECT 108.130000 -122.540000 108.390000 -122.280000 ;
      RECT 108.990000 -124.360000 109.250000 -124.100000 ;
      RECT 108.990000 -124.040000 109.250000 -123.780000 ;
      RECT 108.990000 -122.860000 109.250000 -122.600000 ;
      RECT 108.990000 -122.540000 109.250000 -122.280000 ;
      RECT 110.370000 -124.360000 110.630000 -124.100000 ;
      RECT 110.370000 -124.040000 110.630000 -123.780000 ;
      RECT 111.230000 -124.360000 111.490000 -124.100000 ;
      RECT 111.230000 -124.040000 111.490000 -123.780000 ;
      RECT 113.590000  103.555000 113.850000  103.815000 ;
      RECT 113.590000  103.875000 113.850000  104.135000 ;
      RECT 114.450000  103.555000 114.710000  103.815000 ;
      RECT 114.450000  103.875000 114.710000  104.135000 ;
      RECT 114.880000  102.485000 115.140000  102.745000 ;
      RECT 115.310000  103.555000 115.570000  103.815000 ;
      RECT 115.310000  103.875000 115.570000  104.135000 ;
      RECT 116.170000  103.555000 116.430000  103.815000 ;
      RECT 116.170000  103.875000 116.430000  104.135000 ;
      RECT 117.240000 -122.860000 117.500000 -122.600000 ;
      RECT 117.240000 -122.540000 117.500000 -122.280000 ;
      RECT 117.670000 -124.275000 117.930000 -124.015000 ;
      RECT 117.670000 -123.955000 117.930000 -123.695000 ;
      RECT 118.100000 -122.860000 118.360000 -122.600000 ;
      RECT 118.100000 -122.540000 118.360000 -122.280000 ;
    LAYER via2 ;
      RECT  72.830000  101.215000  73.110000  101.495000 ;
      RECT  72.830000  101.615000  73.110000  101.895000 ;
      RECT  73.690000  101.215000  73.970000  101.495000 ;
      RECT  73.690000  101.615000  73.970000  101.895000 ;
      RECT  74.550000  101.215000  74.830000  101.495000 ;
      RECT  74.550000  101.615000  74.830000  101.895000 ;
      RECT  75.410000  101.215000  75.690000  101.495000 ;
      RECT  75.410000  101.615000  75.690000  101.895000 ;
      RECT  76.910000  101.215000  77.190000  101.495000 ;
      RECT  76.910000  101.615000  77.190000  101.895000 ;
      RECT  77.770000  101.215000  78.050000  101.495000 ;
      RECT  77.770000  101.615000  78.050000  101.895000 ;
      RECT  78.630000  101.215000  78.910000  101.495000 ;
      RECT  78.630000  101.615000  78.910000  101.895000 ;
      RECT  79.490000  101.215000  79.770000  101.495000 ;
      RECT  79.490000  101.615000  79.770000  101.895000 ;
      RECT 105.335000  102.350000 105.615000  102.630000 ;
      RECT 105.335000  102.750000 105.615000  103.030000 ;
      RECT 105.335000  103.850000 105.615000  104.130000 ;
      RECT 105.335000  104.250000 105.615000  104.530000 ;
      RECT 106.195000  102.350000 106.475000  102.630000 ;
      RECT 106.195000  102.750000 106.475000  103.030000 ;
      RECT 106.195000  103.850000 106.475000  104.130000 ;
      RECT 106.195000  104.250000 106.475000  104.530000 ;
      RECT 108.120000 -124.410000 108.400000 -124.130000 ;
      RECT 108.120000 -124.010000 108.400000 -123.730000 ;
      RECT 108.120000 -122.910000 108.400000 -122.630000 ;
      RECT 108.120000 -122.510000 108.400000 -122.230000 ;
      RECT 108.980000 -124.410000 109.260000 -124.130000 ;
      RECT 108.980000 -124.010000 109.260000 -123.730000 ;
      RECT 108.980000 -122.910000 109.260000 -122.630000 ;
      RECT 108.980000 -122.510000 109.260000 -122.230000 ;
      RECT 110.360000 -124.410000 110.640000 -124.130000 ;
      RECT 110.360000 -124.010000 110.640000 -123.730000 ;
      RECT 111.220000 -124.410000 111.500000 -124.130000 ;
      RECT 111.220000 -124.010000 111.500000 -123.730000 ;
      RECT 113.580000  103.505000 113.860000  103.785000 ;
      RECT 113.580000  103.905000 113.860000  104.185000 ;
      RECT 114.440000  103.505000 114.720000  103.785000 ;
      RECT 114.440000  103.905000 114.720000  104.185000 ;
      RECT 115.300000  103.505000 115.580000  103.785000 ;
      RECT 115.300000  103.905000 115.580000  104.185000 ;
      RECT 116.160000  103.505000 116.440000  103.785000 ;
      RECT 116.160000  103.905000 116.440000  104.185000 ;
      RECT 117.230000 -122.910000 117.510000 -122.630000 ;
      RECT 117.230000 -122.510000 117.510000 -122.230000 ;
      RECT 118.090000 -122.910000 118.370000 -122.630000 ;
      RECT 118.090000 -122.510000 118.370000 -122.230000 ;
  END
END sky130_fd_pr__rf_aura_drc_flag_check
END LIBRARY
