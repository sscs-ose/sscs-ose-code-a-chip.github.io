# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.850000 BY  6.100000 ;
  PIN C0
    PORT
      LAYER met4 ;
        RECT 0.000000 0.330000 0.330000 6.100000 ;
        RECT 1.260000 0.330000 1.590000 6.100000 ;
        RECT 2.520000 0.330000 2.850000 6.100000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met4 ;
        RECT 0.630000 0.000000 0.960000 5.770000 ;
        RECT 1.890000 0.000000 2.220000 5.770000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 1.330000 2.820000 1.435000 3.065000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.080000 0.000000 0.250000 6.100000 ;
      RECT 2.600000 0.000000 2.770000 6.100000 ;
    LAYER met1 ;
      RECT 0.080000 0.630000 0.250000 5.770000 ;
      RECT 0.080000 5.770000 2.770000 6.100000 ;
      RECT 0.330000 0.000000 2.520000 0.330000 ;
      RECT 0.390000 0.330000 0.570000 5.470000 ;
      RECT 0.710000 0.630000 0.880000 5.770000 ;
      RECT 1.020000 0.330000 1.200000 5.470000 ;
      RECT 1.340000 0.630000 1.510000 5.770000 ;
      RECT 1.650000 0.330000 1.830000 5.470000 ;
      RECT 1.970000 0.630000 2.140000 5.770000 ;
      RECT 2.280000 0.330000 2.460000 5.470000 ;
      RECT 2.600000 0.630000 2.770000 5.770000 ;
    LAYER met2 ;
      RECT 0.080000 0.630000 0.250000 5.770000 ;
      RECT 0.080000 5.770000 2.770000 6.100000 ;
      RECT 0.330000 0.000000 2.520000 0.330000 ;
      RECT 0.390000 0.330000 0.570000 5.470000 ;
      RECT 0.710000 0.630000 0.880000 5.770000 ;
      RECT 1.020000 0.330000 1.200000 5.470000 ;
      RECT 1.340000 0.630000 1.510000 5.770000 ;
      RECT 1.650000 0.330000 1.830000 5.470000 ;
      RECT 1.970000 0.630000 2.140000 5.770000 ;
      RECT 2.280000 0.330000 2.460000 5.470000 ;
      RECT 2.600000 0.630000 2.770000 5.770000 ;
    LAYER met3 ;
      RECT 0.000000 0.630000 0.330000 5.770000 ;
      RECT 0.000000 5.770000 2.850000 6.100000 ;
      RECT 0.330000 0.000000 2.520000 0.330000 ;
      RECT 0.630000 0.330000 0.960000 5.470000 ;
      RECT 1.260000 0.630000 1.590000 5.770000 ;
      RECT 1.890000 0.330000 2.220000 5.470000 ;
      RECT 2.520000 0.630000 2.850000 5.770000 ;
    LAYER via ;
      RECT 0.295000 5.805000 0.555000 6.065000 ;
      RECT 0.495000 0.035000 0.755000 0.295000 ;
      RECT 0.695000 5.805000 0.955000 6.065000 ;
      RECT 0.895000 0.035000 1.155000 0.295000 ;
      RECT 1.095000 5.805000 1.355000 6.065000 ;
      RECT 1.295000 0.035000 1.555000 0.295000 ;
      RECT 1.495000 5.805000 1.755000 6.065000 ;
      RECT 1.695000 0.035000 1.955000 0.295000 ;
      RECT 1.895000 5.805000 2.155000 6.065000 ;
      RECT 2.095000 0.035000 2.355000 0.295000 ;
      RECT 2.295000 5.805000 2.555000 6.065000 ;
    LAYER via2 ;
      RECT 0.285000 5.795000 0.565000 6.075000 ;
      RECT 0.485000 0.025000 0.765000 0.305000 ;
      RECT 0.685000 5.795000 0.965000 6.075000 ;
      RECT 0.885000 0.025000 1.165000 0.305000 ;
      RECT 1.085000 5.795000 1.365000 6.075000 ;
      RECT 1.285000 0.025000 1.565000 0.305000 ;
      RECT 1.485000 5.795000 1.765000 6.075000 ;
      RECT 1.685000 0.025000 1.965000 0.305000 ;
      RECT 1.885000 5.795000 2.165000 6.075000 ;
      RECT 2.085000 0.025000 2.365000 0.305000 ;
      RECT 2.285000 5.795000 2.565000 6.075000 ;
    LAYER via3 ;
      RECT 0.005000 0.975000 0.325000 1.295000 ;
      RECT 0.005000 1.605000 0.325000 1.925000 ;
      RECT 0.005000 2.235000 0.325000 2.555000 ;
      RECT 0.005000 2.865000 0.325000 3.185000 ;
      RECT 0.005000 3.495000 0.325000 3.815000 ;
      RECT 0.005000 4.125000 0.325000 4.445000 ;
      RECT 0.005000 4.755000 0.325000 5.075000 ;
      RECT 0.005000 5.385000 0.325000 5.705000 ;
      RECT 0.635000 0.660000 0.955000 0.980000 ;
      RECT 0.635000 1.290000 0.955000 1.610000 ;
      RECT 0.635000 1.920000 0.955000 2.240000 ;
      RECT 0.635000 2.550000 0.955000 2.870000 ;
      RECT 0.635000 3.180000 0.955000 3.500000 ;
      RECT 0.635000 3.810000 0.955000 4.130000 ;
      RECT 0.635000 4.440000 0.955000 4.760000 ;
      RECT 0.635000 5.070000 0.955000 5.390000 ;
      RECT 1.265000 0.975000 1.585000 1.295000 ;
      RECT 1.265000 1.605000 1.585000 1.925000 ;
      RECT 1.265000 2.235000 1.585000 2.555000 ;
      RECT 1.265000 2.865000 1.585000 3.185000 ;
      RECT 1.265000 3.495000 1.585000 3.815000 ;
      RECT 1.265000 4.125000 1.585000 4.445000 ;
      RECT 1.265000 4.755000 1.585000 5.075000 ;
      RECT 1.265000 5.385000 1.585000 5.705000 ;
      RECT 1.895000 0.660000 2.215000 0.980000 ;
      RECT 1.895000 1.290000 2.215000 1.610000 ;
      RECT 1.895000 1.920000 2.215000 2.240000 ;
      RECT 1.895000 2.550000 2.215000 2.870000 ;
      RECT 1.895000 3.180000 2.215000 3.500000 ;
      RECT 1.895000 3.810000 2.215000 4.130000 ;
      RECT 1.895000 4.440000 2.215000 4.760000 ;
      RECT 1.895000 5.070000 2.215000 5.390000 ;
      RECT 2.525000 0.975000 2.845000 1.295000 ;
      RECT 2.525000 1.605000 2.845000 1.925000 ;
      RECT 2.525000 2.235000 2.845000 2.555000 ;
      RECT 2.525000 2.865000 2.845000 3.185000 ;
      RECT 2.525000 3.495000 2.845000 3.815000 ;
      RECT 2.525000 4.125000 2.845000 4.445000 ;
      RECT 2.525000 4.755000 2.845000 5.075000 ;
      RECT 2.525000 5.385000 2.845000 5.705000 ;
  END
END sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2
END LIBRARY
