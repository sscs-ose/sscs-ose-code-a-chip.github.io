# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.380000 BY  3.930000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2.090000 3.380000 3.370000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.806000 ;
    PORT
      LAYER li1 ;
        RECT 0.845000 0.100000 2.535000 0.270000 ;
        RECT 0.845000 3.660000 2.535000 3.830000 ;
      LAYER mcon ;
        RECT 0.885000 0.100000 1.055000 0.270000 ;
        RECT 0.885000 3.660000 1.055000 3.830000 ;
        RECT 1.245000 0.100000 1.415000 0.270000 ;
        RECT 1.245000 3.660000 1.415000 3.830000 ;
        RECT 1.605000 0.100000 1.775000 0.270000 ;
        RECT 1.605000 3.660000 1.775000 3.830000 ;
        RECT 1.965000 0.100000 2.135000 0.270000 ;
        RECT 1.965000 3.660000 2.135000 3.830000 ;
        RECT 2.325000 0.100000 2.495000 0.270000 ;
        RECT 2.325000 3.660000 2.495000 3.830000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.825000 0.000000 2.555000 0.330000 ;
        RECT 0.825000 3.600000 2.555000 3.930000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.528400 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.560000 3.380000 1.840000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.872900 ;
    PORT
      LAYER met1 ;
        RECT 0.130000 0.560000 0.420000 3.370000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.960000 0.560000 3.250000 3.370000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.190000 0.610000 0.360000 3.320000 ;
      RECT 0.745000 0.440000 0.915000 3.490000 ;
      RECT 1.175000 0.440000 1.345000 3.490000 ;
      RECT 1.605000 0.440000 1.775000 3.490000 ;
      RECT 2.035000 0.440000 2.205000 3.490000 ;
      RECT 2.465000 0.440000 2.635000 3.490000 ;
      RECT 3.020000 0.610000 3.190000 3.320000 ;
    LAYER mcon ;
      RECT 0.190000 0.620000 0.360000 0.790000 ;
      RECT 0.190000 0.980000 0.360000 1.150000 ;
      RECT 0.190000 1.340000 0.360000 1.510000 ;
      RECT 0.190000 1.700000 0.360000 1.870000 ;
      RECT 0.190000 2.060000 0.360000 2.230000 ;
      RECT 0.190000 2.420000 0.360000 2.590000 ;
      RECT 0.190000 2.780000 0.360000 2.950000 ;
      RECT 0.190000 3.140000 0.360000 3.310000 ;
      RECT 0.745000 0.620000 0.915000 0.790000 ;
      RECT 0.745000 0.980000 0.915000 1.150000 ;
      RECT 0.745000 1.340000 0.915000 1.510000 ;
      RECT 0.745000 1.700000 0.915000 1.870000 ;
      RECT 0.745000 2.060000 0.915000 2.230000 ;
      RECT 0.745000 2.420000 0.915000 2.590000 ;
      RECT 0.745000 2.780000 0.915000 2.950000 ;
      RECT 0.745000 3.140000 0.915000 3.310000 ;
      RECT 1.175000 0.620000 1.345000 0.790000 ;
      RECT 1.175000 0.980000 1.345000 1.150000 ;
      RECT 1.175000 1.340000 1.345000 1.510000 ;
      RECT 1.175000 1.700000 1.345000 1.870000 ;
      RECT 1.175000 2.060000 1.345000 2.230000 ;
      RECT 1.175000 2.420000 1.345000 2.590000 ;
      RECT 1.175000 2.780000 1.345000 2.950000 ;
      RECT 1.175000 3.140000 1.345000 3.310000 ;
      RECT 1.605000 0.620000 1.775000 0.790000 ;
      RECT 1.605000 0.980000 1.775000 1.150000 ;
      RECT 1.605000 1.340000 1.775000 1.510000 ;
      RECT 1.605000 1.700000 1.775000 1.870000 ;
      RECT 1.605000 2.060000 1.775000 2.230000 ;
      RECT 1.605000 2.420000 1.775000 2.590000 ;
      RECT 1.605000 2.780000 1.775000 2.950000 ;
      RECT 1.605000 3.140000 1.775000 3.310000 ;
      RECT 2.035000 0.620000 2.205000 0.790000 ;
      RECT 2.035000 0.980000 2.205000 1.150000 ;
      RECT 2.035000 1.340000 2.205000 1.510000 ;
      RECT 2.035000 1.700000 2.205000 1.870000 ;
      RECT 2.035000 2.060000 2.205000 2.230000 ;
      RECT 2.035000 2.420000 2.205000 2.590000 ;
      RECT 2.035000 2.780000 2.205000 2.950000 ;
      RECT 2.035000 3.140000 2.205000 3.310000 ;
      RECT 2.465000 0.620000 2.635000 0.790000 ;
      RECT 2.465000 0.980000 2.635000 1.150000 ;
      RECT 2.465000 1.340000 2.635000 1.510000 ;
      RECT 2.465000 1.700000 2.635000 1.870000 ;
      RECT 2.465000 2.060000 2.635000 2.230000 ;
      RECT 2.465000 2.420000 2.635000 2.590000 ;
      RECT 2.465000 2.780000 2.635000 2.950000 ;
      RECT 2.465000 3.140000 2.635000 3.310000 ;
      RECT 3.020000 0.620000 3.190000 0.790000 ;
      RECT 3.020000 0.980000 3.190000 1.150000 ;
      RECT 3.020000 1.340000 3.190000 1.510000 ;
      RECT 3.020000 1.700000 3.190000 1.870000 ;
      RECT 3.020000 2.060000 3.190000 2.230000 ;
      RECT 3.020000 2.420000 3.190000 2.590000 ;
      RECT 3.020000 2.780000 3.190000 2.950000 ;
      RECT 3.020000 3.140000 3.190000 3.310000 ;
    LAYER met1 ;
      RECT 0.700000 0.560000 0.960000 3.370000 ;
      RECT 1.130000 0.560000 1.390000 3.370000 ;
      RECT 1.560000 0.560000 1.820000 3.370000 ;
      RECT 1.990000 0.560000 2.250000 3.370000 ;
      RECT 2.420000 0.560000 2.680000 3.370000 ;
    LAYER via ;
      RECT 0.700000 0.590000 0.960000 0.850000 ;
      RECT 0.700000 0.910000 0.960000 1.170000 ;
      RECT 0.700000 1.230000 0.960000 1.490000 ;
      RECT 0.700000 1.550000 0.960000 1.810000 ;
      RECT 1.130000 2.120000 1.390000 2.380000 ;
      RECT 1.130000 2.440000 1.390000 2.700000 ;
      RECT 1.130000 2.760000 1.390000 3.020000 ;
      RECT 1.130000 3.080000 1.390000 3.340000 ;
      RECT 1.560000 0.590000 1.820000 0.850000 ;
      RECT 1.560000 0.910000 1.820000 1.170000 ;
      RECT 1.560000 1.230000 1.820000 1.490000 ;
      RECT 1.560000 1.550000 1.820000 1.810000 ;
      RECT 1.990000 2.120000 2.250000 2.380000 ;
      RECT 1.990000 2.440000 2.250000 2.700000 ;
      RECT 1.990000 2.760000 2.250000 3.020000 ;
      RECT 1.990000 3.080000 2.250000 3.340000 ;
      RECT 2.420000 0.590000 2.680000 0.850000 ;
      RECT 2.420000 0.910000 2.680000 1.170000 ;
      RECT 2.420000 1.230000 2.680000 1.490000 ;
      RECT 2.420000 1.550000 2.680000 1.810000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15
END LIBRARY
