# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15 ;
  ORIGIN  0.050000  0.000000 ;
  SIZE  4.515000 BY  6.460000 ;
  PIN DRAIN
    ANTENNADIFFAREA  6.262000 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2.110000 4.420000 4.350000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.030000 ;
    PORT
      LAYER met1 ;
        RECT 0.910000 0.170000 3.720000 0.460000 ;
        RECT 0.910000 6.000000 3.720000 6.290000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  6.034750 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.690000 4.420000 1.970000 ;
        RECT 0.000000 4.490000 4.420000 5.775000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.190000 0.805000 0.360000 5.655000 ;
      RECT 0.745000 0.685000 0.915000 5.775000 ;
      RECT 0.970000 0.230000 3.680000 0.400000 ;
      RECT 0.970000 6.060000 3.680000 6.230000 ;
      RECT 1.165000 0.685000 1.695000 5.775000 ;
      RECT 1.935000 0.685000 2.465000 5.775000 ;
      RECT 2.705000 0.685000 3.235000 5.775000 ;
      RECT 3.485000 0.685000 3.655000 5.775000 ;
      RECT 4.055000 0.805000 4.225000 5.655000 ;
    LAYER mcon ;
      RECT 0.190000 1.165000 0.360000 1.335000 ;
      RECT 0.190000 1.525000 0.360000 1.695000 ;
      RECT 0.190000 1.885000 0.360000 2.055000 ;
      RECT 0.190000 2.245000 0.360000 2.415000 ;
      RECT 0.190000 2.605000 0.360000 2.775000 ;
      RECT 0.190000 2.965000 0.360000 3.135000 ;
      RECT 0.190000 3.325000 0.360000 3.495000 ;
      RECT 0.190000 3.685000 0.360000 3.855000 ;
      RECT 0.190000 4.045000 0.360000 4.215000 ;
      RECT 0.190000 4.405000 0.360000 4.575000 ;
      RECT 0.190000 4.765000 0.360000 4.935000 ;
      RECT 0.190000 5.125000 0.360000 5.295000 ;
      RECT 0.190000 5.485000 0.360000 5.655000 ;
      RECT 0.745000 0.805000 0.915000 0.975000 ;
      RECT 0.745000 1.165000 0.915000 1.335000 ;
      RECT 0.745000 1.525000 0.915000 1.695000 ;
      RECT 0.745000 1.885000 0.915000 2.055000 ;
      RECT 0.745000 2.245000 0.915000 2.415000 ;
      RECT 0.745000 2.605000 0.915000 2.775000 ;
      RECT 0.745000 2.965000 0.915000 3.135000 ;
      RECT 0.745000 3.325000 0.915000 3.495000 ;
      RECT 0.745000 3.685000 0.915000 3.855000 ;
      RECT 0.745000 4.045000 0.915000 4.215000 ;
      RECT 0.745000 4.405000 0.915000 4.575000 ;
      RECT 0.745000 4.765000 0.915000 4.935000 ;
      RECT 0.745000 5.125000 0.915000 5.295000 ;
      RECT 0.745000 5.485000 0.915000 5.655000 ;
      RECT 0.970000 0.230000 1.140000 0.400000 ;
      RECT 0.970000 6.060000 1.140000 6.230000 ;
      RECT 1.165000 0.805000 1.695000 5.655000 ;
      RECT 1.330000 0.230000 1.500000 0.400000 ;
      RECT 1.330000 6.060000 1.500000 6.230000 ;
      RECT 1.690000 0.230000 1.860000 0.400000 ;
      RECT 1.690000 6.060000 1.860000 6.230000 ;
      RECT 1.935000 0.805000 2.465000 5.655000 ;
      RECT 2.050000 0.230000 2.220000 0.400000 ;
      RECT 2.050000 6.060000 2.220000 6.230000 ;
      RECT 2.410000 0.230000 2.580000 0.400000 ;
      RECT 2.410000 6.060000 2.580000 6.230000 ;
      RECT 2.705000 0.805000 3.235000 5.655000 ;
      RECT 2.770000 0.230000 2.940000 0.400000 ;
      RECT 2.770000 6.060000 2.940000 6.230000 ;
      RECT 3.130000 0.230000 3.300000 0.400000 ;
      RECT 3.130000 6.060000 3.300000 6.230000 ;
      RECT 3.485000 0.805000 3.655000 0.975000 ;
      RECT 3.485000 1.165000 3.655000 1.335000 ;
      RECT 3.485000 1.525000 3.655000 1.695000 ;
      RECT 3.485000 1.885000 3.655000 2.055000 ;
      RECT 3.485000 2.245000 3.655000 2.415000 ;
      RECT 3.485000 2.605000 3.655000 2.775000 ;
      RECT 3.485000 2.965000 3.655000 3.135000 ;
      RECT 3.485000 3.325000 3.655000 3.495000 ;
      RECT 3.485000 3.685000 3.655000 3.855000 ;
      RECT 3.485000 4.045000 3.655000 4.215000 ;
      RECT 3.485000 4.405000 3.655000 4.575000 ;
      RECT 3.485000 4.765000 3.655000 4.935000 ;
      RECT 3.485000 5.125000 3.655000 5.295000 ;
      RECT 3.485000 5.485000 3.655000 5.655000 ;
      RECT 3.490000 0.230000 3.660000 0.400000 ;
      RECT 3.490000 6.060000 3.660000 6.230000 ;
      RECT 4.055000 1.165000 4.225000 1.335000 ;
      RECT 4.055000 1.525000 4.225000 1.695000 ;
      RECT 4.055000 1.885000 4.225000 2.055000 ;
      RECT 4.055000 2.245000 4.225000 2.415000 ;
      RECT 4.055000 2.605000 4.225000 2.775000 ;
      RECT 4.055000 2.965000 4.225000 3.135000 ;
      RECT 4.055000 3.325000 4.225000 3.495000 ;
      RECT 4.055000 3.685000 4.225000 3.855000 ;
      RECT 4.055000 4.045000 4.225000 4.215000 ;
      RECT 4.055000 4.405000 4.225000 4.575000 ;
      RECT 4.055000 4.765000 4.225000 4.935000 ;
      RECT 4.055000 5.125000 4.225000 5.295000 ;
      RECT 4.055000 5.485000 4.225000 5.655000 ;
    LAYER met1 ;
      RECT 0.130000 0.745000 0.420000 5.715000 ;
      RECT 0.700000 0.690000 0.960000 0.745000 ;
      RECT 0.700000 0.745000 0.975000 5.715000 ;
      RECT 0.700000 5.715000 0.960000 5.770000 ;
      RECT 1.115000 0.745000 1.745000 5.715000 ;
      RECT 1.885000 0.745000 2.515000 5.715000 ;
      RECT 1.910000 5.715000 2.490000 5.775000 ;
      RECT 2.655000 0.745000 3.285000 5.715000 ;
      RECT 3.425000 0.745000 3.715000 5.715000 ;
      RECT 3.440000 0.690000 3.700000 0.745000 ;
      RECT 3.440000 5.715000 3.700000 5.775000 ;
      RECT 3.995000 0.745000 4.285000 5.715000 ;
    LAYER via ;
      RECT 0.700000 0.720000 0.960000 0.980000 ;
      RECT 0.700000 1.040000 0.960000 1.300000 ;
      RECT 0.700000 1.360000 0.960000 1.620000 ;
      RECT 0.700000 1.680000 0.960000 1.940000 ;
      RECT 0.700000 4.520000 0.960000 4.780000 ;
      RECT 0.700000 4.840000 0.960000 5.100000 ;
      RECT 0.700000 5.160000 0.960000 5.420000 ;
      RECT 0.700000 5.480000 0.960000 5.740000 ;
      RECT 1.140000 2.140000 1.720000 4.320000 ;
      RECT 1.910000 4.525000 2.490000 5.745000 ;
      RECT 2.680000 2.140000 3.260000 4.320000 ;
      RECT 3.440000 0.720000 3.700000 0.980000 ;
      RECT 3.440000 1.040000 3.700000 1.300000 ;
      RECT 3.440000 1.360000 3.700000 1.620000 ;
      RECT 3.440000 1.680000 3.700000 1.940000 ;
      RECT 3.440000 4.525000 3.700000 4.785000 ;
      RECT 3.440000 4.845000 3.700000 5.105000 ;
      RECT 3.440000 5.165000 3.700000 5.425000 ;
      RECT 3.440000 5.485000 3.700000 5.745000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15
END LIBRARY
