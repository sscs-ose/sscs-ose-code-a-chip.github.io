# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_npn_05v5_W2p00L2p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_npn_05v5_W2p00L2p00 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  10.70000 BY  10.70000 ;
  OBS
    LAYER li1 ;
      RECT  0.170000  0.170000 10.790000  0.500000 ;
      RECT  0.170000  0.500000  0.500000 10.460000 ;
      RECT  0.170000 10.460000 10.790000 10.790000 ;
      RECT  1.300000  1.300000  9.660000  1.630000 ;
      RECT  1.300000  1.630000  1.630000  9.330000 ;
      RECT  1.300000  9.330000  9.660000  9.660000 ;
      RECT  3.310000  3.310000  7.650000  3.640000 ;
      RECT  3.310000  3.640000  3.640000  7.320000 ;
      RECT  3.310000  7.320000  7.650000  7.650000 ;
      RECT  4.465000  4.465000  6.495000  6.495000 ;
      RECT  7.320000  3.640000  7.650000  7.320000 ;
      RECT  9.330000  1.630000  9.660000  9.330000 ;
      RECT 10.460000  0.500000 10.790000 10.460000 ;
    LAYER mcon ;
      RECT  0.250000  0.250000  0.420000  0.420000 ;
      RECT  0.250000  0.715000  0.420000  0.885000 ;
      RECT  0.250000  1.075000  0.420000  1.245000 ;
      RECT  0.250000  1.435000  0.420000  1.605000 ;
      RECT  0.250000  1.795000  0.420000  1.965000 ;
      RECT  0.250000  2.155000  0.420000  2.325000 ;
      RECT  0.250000  2.515000  0.420000  2.685000 ;
      RECT  0.250000  2.875000  0.420000  3.045000 ;
      RECT  0.250000  3.235000  0.420000  3.405000 ;
      RECT  0.250000  3.595000  0.420000  3.765000 ;
      RECT  0.250000  3.955000  0.420000  4.125000 ;
      RECT  0.250000  4.315000  0.420000  4.485000 ;
      RECT  0.250000  4.675000  0.420000  4.845000 ;
      RECT  0.250000  5.035000  0.420000  5.205000 ;
      RECT  0.250000  5.395000  0.420000  5.565000 ;
      RECT  0.250000  5.755000  0.420000  5.925000 ;
      RECT  0.250000  6.115000  0.420000  6.285000 ;
      RECT  0.250000  6.475000  0.420000  6.645000 ;
      RECT  0.250000  6.835000  0.420000  7.005000 ;
      RECT  0.250000  7.195000  0.420000  7.365000 ;
      RECT  0.250000  7.555000  0.420000  7.725000 ;
      RECT  0.250000  7.915000  0.420000  8.085000 ;
      RECT  0.250000  8.275000  0.420000  8.445000 ;
      RECT  0.250000  8.635000  0.420000  8.805000 ;
      RECT  0.250000  8.995000  0.420000  9.165000 ;
      RECT  0.250000  9.355000  0.420000  9.525000 ;
      RECT  0.250000  9.715000  0.420000  9.885000 ;
      RECT  0.250000 10.075000  0.420000 10.245000 ;
      RECT  0.250000 10.540000  0.420000 10.710000 ;
      RECT  0.715000  0.250000  0.885000  0.420000 ;
      RECT  0.715000 10.540000  0.885000 10.710000 ;
      RECT  1.075000  0.250000  1.245000  0.420000 ;
      RECT  1.075000 10.540000  1.245000 10.710000 ;
      RECT  1.380000  1.380000  1.550000  1.550000 ;
      RECT  1.380000  1.795000  1.550000  1.965000 ;
      RECT  1.380000  2.155000  1.550000  2.325000 ;
      RECT  1.380000  2.515000  1.550000  2.685000 ;
      RECT  1.380000  2.875000  1.550000  3.045000 ;
      RECT  1.380000  3.235000  1.550000  3.405000 ;
      RECT  1.380000  3.595000  1.550000  3.765000 ;
      RECT  1.380000  3.955000  1.550000  4.125000 ;
      RECT  1.380000  4.315000  1.550000  4.485000 ;
      RECT  1.380000  4.675000  1.550000  4.845000 ;
      RECT  1.380000  5.035000  1.550000  5.205000 ;
      RECT  1.380000  5.395000  1.550000  5.565000 ;
      RECT  1.380000  5.755000  1.550000  5.925000 ;
      RECT  1.380000  6.115000  1.550000  6.285000 ;
      RECT  1.380000  6.475000  1.550000  6.645000 ;
      RECT  1.380000  6.835000  1.550000  7.005000 ;
      RECT  1.380000  7.195000  1.550000  7.365000 ;
      RECT  1.380000  7.555000  1.550000  7.725000 ;
      RECT  1.380000  7.915000  1.550000  8.085000 ;
      RECT  1.380000  8.275000  1.550000  8.445000 ;
      RECT  1.380000  8.635000  1.550000  8.805000 ;
      RECT  1.380000  8.995000  1.550000  9.165000 ;
      RECT  1.380000  9.410000  1.550000  9.580000 ;
      RECT  1.435000  0.250000  1.605000  0.420000 ;
      RECT  1.435000 10.540000  1.605000 10.710000 ;
      RECT  1.795000  0.250000  1.965000  0.420000 ;
      RECT  1.795000  1.380000  1.965000  1.550000 ;
      RECT  1.795000  9.410000  1.965000  9.580000 ;
      RECT  1.795000 10.540000  1.965000 10.710000 ;
      RECT  2.155000  0.250000  2.325000  0.420000 ;
      RECT  2.155000  1.380000  2.325000  1.550000 ;
      RECT  2.155000  9.410000  2.325000  9.580000 ;
      RECT  2.155000 10.540000  2.325000 10.710000 ;
      RECT  2.515000  0.250000  2.685000  0.420000 ;
      RECT  2.515000  1.380000  2.685000  1.550000 ;
      RECT  2.515000  9.410000  2.685000  9.580000 ;
      RECT  2.515000 10.540000  2.685000 10.710000 ;
      RECT  2.875000  0.250000  3.045000  0.420000 ;
      RECT  2.875000  1.380000  3.045000  1.550000 ;
      RECT  2.875000  9.410000  3.045000  9.580000 ;
      RECT  2.875000 10.540000  3.045000 10.710000 ;
      RECT  3.235000  0.250000  3.405000  0.420000 ;
      RECT  3.235000  1.380000  3.405000  1.550000 ;
      RECT  3.235000  9.410000  3.405000  9.580000 ;
      RECT  3.235000 10.540000  3.405000 10.710000 ;
      RECT  3.390000  3.390000  3.560000  3.560000 ;
      RECT  3.390000  3.775000  3.560000  3.945000 ;
      RECT  3.390000  4.135000  3.560000  4.305000 ;
      RECT  3.390000  4.495000  3.560000  4.665000 ;
      RECT  3.390000  4.855000  3.560000  5.025000 ;
      RECT  3.390000  5.215000  3.560000  5.385000 ;
      RECT  3.390000  5.575000  3.560000  5.745000 ;
      RECT  3.390000  5.935000  3.560000  6.105000 ;
      RECT  3.390000  6.295000  3.560000  6.465000 ;
      RECT  3.390000  6.655000  3.560000  6.825000 ;
      RECT  3.390000  7.015000  3.560000  7.185000 ;
      RECT  3.390000  7.400000  3.560000  7.570000 ;
      RECT  3.595000  0.250000  3.765000  0.420000 ;
      RECT  3.595000  1.380000  3.765000  1.550000 ;
      RECT  3.595000  9.410000  3.765000  9.580000 ;
      RECT  3.595000 10.540000  3.765000 10.710000 ;
      RECT  3.775000  3.390000  3.945000  3.560000 ;
      RECT  3.775000  7.400000  3.945000  7.570000 ;
      RECT  3.955000  0.250000  4.125000  0.420000 ;
      RECT  3.955000  1.380000  4.125000  1.550000 ;
      RECT  3.955000  9.410000  4.125000  9.580000 ;
      RECT  3.955000 10.540000  4.125000 10.710000 ;
      RECT  4.135000  3.390000  4.305000  3.560000 ;
      RECT  4.135000  7.400000  4.305000  7.570000 ;
      RECT  4.315000  0.250000  4.485000  0.420000 ;
      RECT  4.315000  1.380000  4.485000  1.550000 ;
      RECT  4.315000  9.410000  4.485000  9.580000 ;
      RECT  4.315000 10.540000  4.485000 10.710000 ;
      RECT  4.495000  3.390000  4.665000  3.560000 ;
      RECT  4.495000  7.400000  4.665000  7.570000 ;
      RECT  4.675000  0.250000  4.845000  0.420000 ;
      RECT  4.675000  1.380000  4.845000  1.550000 ;
      RECT  4.675000  4.675000  6.285000  6.285000 ;
      RECT  4.675000  9.410000  4.845000  9.580000 ;
      RECT  4.675000 10.540000  4.845000 10.710000 ;
      RECT  4.855000  3.390000  5.025000  3.560000 ;
      RECT  4.855000  7.400000  5.025000  7.570000 ;
      RECT  5.035000  0.250000  5.205000  0.420000 ;
      RECT  5.035000  1.380000  5.205000  1.550000 ;
      RECT  5.035000  9.410000  5.205000  9.580000 ;
      RECT  5.035000 10.540000  5.205000 10.710000 ;
      RECT  5.215000  3.390000  5.385000  3.560000 ;
      RECT  5.215000  7.400000  5.385000  7.570000 ;
      RECT  5.395000  0.250000  5.565000  0.420000 ;
      RECT  5.395000  1.380000  5.565000  1.550000 ;
      RECT  5.395000  9.410000  5.565000  9.580000 ;
      RECT  5.395000 10.540000  5.565000 10.710000 ;
      RECT  5.575000  3.390000  5.745000  3.560000 ;
      RECT  5.575000  7.400000  5.745000  7.570000 ;
      RECT  5.755000  0.250000  5.925000  0.420000 ;
      RECT  5.755000  1.380000  5.925000  1.550000 ;
      RECT  5.755000  9.410000  5.925000  9.580000 ;
      RECT  5.755000 10.540000  5.925000 10.710000 ;
      RECT  5.935000  3.390000  6.105000  3.560000 ;
      RECT  5.935000  7.400000  6.105000  7.570000 ;
      RECT  6.115000  0.250000  6.285000  0.420000 ;
      RECT  6.115000  1.380000  6.285000  1.550000 ;
      RECT  6.115000  9.410000  6.285000  9.580000 ;
      RECT  6.115000 10.540000  6.285000 10.710000 ;
      RECT  6.295000  3.390000  6.465000  3.560000 ;
      RECT  6.295000  7.400000  6.465000  7.570000 ;
      RECT  6.475000  0.250000  6.645000  0.420000 ;
      RECT  6.475000  1.380000  6.645000  1.550000 ;
      RECT  6.475000  9.410000  6.645000  9.580000 ;
      RECT  6.475000 10.540000  6.645000 10.710000 ;
      RECT  6.655000  3.390000  6.825000  3.560000 ;
      RECT  6.655000  7.400000  6.825000  7.570000 ;
      RECT  6.835000  0.250000  7.005000  0.420000 ;
      RECT  6.835000  1.380000  7.005000  1.550000 ;
      RECT  6.835000  9.410000  7.005000  9.580000 ;
      RECT  6.835000 10.540000  7.005000 10.710000 ;
      RECT  7.015000  3.390000  7.185000  3.560000 ;
      RECT  7.015000  7.400000  7.185000  7.570000 ;
      RECT  7.195000  0.250000  7.365000  0.420000 ;
      RECT  7.195000  1.380000  7.365000  1.550000 ;
      RECT  7.195000  9.410000  7.365000  9.580000 ;
      RECT  7.195000 10.540000  7.365000 10.710000 ;
      RECT  7.400000  3.390000  7.570000  3.560000 ;
      RECT  7.400000  3.775000  7.570000  3.945000 ;
      RECT  7.400000  4.135000  7.570000  4.305000 ;
      RECT  7.400000  4.495000  7.570000  4.665000 ;
      RECT  7.400000  4.855000  7.570000  5.025000 ;
      RECT  7.400000  5.215000  7.570000  5.385000 ;
      RECT  7.400000  5.575000  7.570000  5.745000 ;
      RECT  7.400000  5.935000  7.570000  6.105000 ;
      RECT  7.400000  6.295000  7.570000  6.465000 ;
      RECT  7.400000  6.655000  7.570000  6.825000 ;
      RECT  7.400000  7.015000  7.570000  7.185000 ;
      RECT  7.400000  7.400000  7.570000  7.570000 ;
      RECT  7.555000  0.250000  7.725000  0.420000 ;
      RECT  7.555000  1.380000  7.725000  1.550000 ;
      RECT  7.555000  9.410000  7.725000  9.580000 ;
      RECT  7.555000 10.540000  7.725000 10.710000 ;
      RECT  7.915000  0.250000  8.085000  0.420000 ;
      RECT  7.915000  1.380000  8.085000  1.550000 ;
      RECT  7.915000  9.410000  8.085000  9.580000 ;
      RECT  7.915000 10.540000  8.085000 10.710000 ;
      RECT  8.275000  0.250000  8.445000  0.420000 ;
      RECT  8.275000  1.380000  8.445000  1.550000 ;
      RECT  8.275000  9.410000  8.445000  9.580000 ;
      RECT  8.275000 10.540000  8.445000 10.710000 ;
      RECT  8.635000  0.250000  8.805000  0.420000 ;
      RECT  8.635000  1.380000  8.805000  1.550000 ;
      RECT  8.635000  9.410000  8.805000  9.580000 ;
      RECT  8.635000 10.540000  8.805000 10.710000 ;
      RECT  8.995000  0.250000  9.165000  0.420000 ;
      RECT  8.995000  1.380000  9.165000  1.550000 ;
      RECT  8.995000  9.410000  9.165000  9.580000 ;
      RECT  8.995000 10.540000  9.165000 10.710000 ;
      RECT  9.355000  0.250000  9.525000  0.420000 ;
      RECT  9.355000 10.540000  9.525000 10.710000 ;
      RECT  9.410000  1.380000  9.580000  1.550000 ;
      RECT  9.410000  1.795000  9.580000  1.965000 ;
      RECT  9.410000  2.155000  9.580000  2.325000 ;
      RECT  9.410000  2.515000  9.580000  2.685000 ;
      RECT  9.410000  2.875000  9.580000  3.045000 ;
      RECT  9.410000  3.235000  9.580000  3.405000 ;
      RECT  9.410000  3.595000  9.580000  3.765000 ;
      RECT  9.410000  3.955000  9.580000  4.125000 ;
      RECT  9.410000  4.315000  9.580000  4.485000 ;
      RECT  9.410000  4.675000  9.580000  4.845000 ;
      RECT  9.410000  5.035000  9.580000  5.205000 ;
      RECT  9.410000  5.395000  9.580000  5.565000 ;
      RECT  9.410000  5.755000  9.580000  5.925000 ;
      RECT  9.410000  6.115000  9.580000  6.285000 ;
      RECT  9.410000  6.475000  9.580000  6.645000 ;
      RECT  9.410000  6.835000  9.580000  7.005000 ;
      RECT  9.410000  7.195000  9.580000  7.365000 ;
      RECT  9.410000  7.555000  9.580000  7.725000 ;
      RECT  9.410000  7.915000  9.580000  8.085000 ;
      RECT  9.410000  8.275000  9.580000  8.445000 ;
      RECT  9.410000  8.635000  9.580000  8.805000 ;
      RECT  9.410000  8.995000  9.580000  9.165000 ;
      RECT  9.410000  9.410000  9.580000  9.580000 ;
      RECT  9.715000  0.250000  9.885000  0.420000 ;
      RECT  9.715000 10.540000  9.885000 10.710000 ;
      RECT 10.075000  0.250000 10.245000  0.420000 ;
      RECT 10.075000 10.540000 10.245000 10.710000 ;
      RECT 10.540000  0.250000 10.710000  0.420000 ;
      RECT 10.540000  0.715000 10.710000  0.885000 ;
      RECT 10.540000  1.075000 10.710000  1.245000 ;
      RECT 10.540000  1.435000 10.710000  1.605000 ;
      RECT 10.540000  1.795000 10.710000  1.965000 ;
      RECT 10.540000  2.155000 10.710000  2.325000 ;
      RECT 10.540000  2.515000 10.710000  2.685000 ;
      RECT 10.540000  2.875000 10.710000  3.045000 ;
      RECT 10.540000  3.235000 10.710000  3.405000 ;
      RECT 10.540000  3.595000 10.710000  3.765000 ;
      RECT 10.540000  3.955000 10.710000  4.125000 ;
      RECT 10.540000  4.315000 10.710000  4.485000 ;
      RECT 10.540000  4.675000 10.710000  4.845000 ;
      RECT 10.540000  5.035000 10.710000  5.205000 ;
      RECT 10.540000  5.395000 10.710000  5.565000 ;
      RECT 10.540000  5.755000 10.710000  5.925000 ;
      RECT 10.540000  6.115000 10.710000  6.285000 ;
      RECT 10.540000  6.475000 10.710000  6.645000 ;
      RECT 10.540000  6.835000 10.710000  7.005000 ;
      RECT 10.540000  7.195000 10.710000  7.365000 ;
      RECT 10.540000  7.555000 10.710000  7.725000 ;
      RECT 10.540000  7.915000 10.710000  8.085000 ;
      RECT 10.540000  8.275000 10.710000  8.445000 ;
      RECT 10.540000  8.635000 10.710000  8.805000 ;
      RECT 10.540000  8.995000 10.710000  9.165000 ;
      RECT 10.540000  9.355000 10.710000  9.525000 ;
      RECT 10.540000  9.715000 10.710000  9.885000 ;
      RECT 10.540000 10.075000 10.710000 10.245000 ;
      RECT 10.540000 10.540000 10.710000 10.710000 ;
    LAYER met1 ;
      RECT  0.190000  0.190000 10.770000  0.480000 ;
      RECT  0.190000  0.480000  0.480000 10.480000 ;
      RECT  0.190000 10.480000 10.770000 10.770000 ;
      RECT  1.320000  1.320000  9.640000  1.610000 ;
      RECT  1.320000  1.610000  1.610000  9.350000 ;
      RECT  1.320000  9.350000  9.640000  9.640000 ;
      RECT  3.330000  3.330000  7.630000  3.620000 ;
      RECT  3.330000  3.620000  3.620000  7.340000 ;
      RECT  3.330000  7.340000  7.630000  7.630000 ;
      RECT  4.615000  4.615000  6.345000  6.345000 ;
      RECT  7.340000  3.620000  7.630000  7.340000 ;
      RECT  9.350000  1.610000  9.640000  9.350000 ;
      RECT 10.480000  0.480000 10.770000 10.480000 ;
  END
END sky130_fd_pr__rf_npn_05v5_W2p00L2p00
END LIBRARY
