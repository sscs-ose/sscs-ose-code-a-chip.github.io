.param w1_2=7.49
.param w3_4=2.64
.param w5_6=59.49
.param w7_8=21.0
.param w9_10=14.98
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=65u
.param iref_post_layout=70u
