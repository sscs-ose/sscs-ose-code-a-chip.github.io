# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50 ;
  ORIGIN -0.050000  0.000000 ;
  SIZE  9.700000 BY  8.010000 ;
  PIN DRAIN
    ANTENNADIFFAREA  9.926000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.405000 9.750000 5.605000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  35.450001 ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.100000 8.805000 0.270000 ;
        RECT 0.995000 7.740000 8.805000 7.910000 ;
      LAYER mcon ;
        RECT 1.035000 0.100000 1.205000 0.270000 ;
        RECT 1.035000 7.740000 1.205000 7.910000 ;
        RECT 1.395000 0.100000 1.565000 0.270000 ;
        RECT 1.395000 7.740000 1.565000 7.910000 ;
        RECT 1.755000 0.100000 1.925000 0.270000 ;
        RECT 1.755000 7.740000 1.925000 7.910000 ;
        RECT 2.115000 0.100000 2.285000 0.270000 ;
        RECT 2.115000 7.740000 2.285000 7.910000 ;
        RECT 2.475000 0.100000 2.645000 0.270000 ;
        RECT 2.475000 7.740000 2.645000 7.910000 ;
        RECT 2.835000 0.100000 3.005000 0.270000 ;
        RECT 2.835000 7.740000 3.005000 7.910000 ;
        RECT 3.195000 0.100000 3.365000 0.270000 ;
        RECT 3.195000 7.740000 3.365000 7.910000 ;
        RECT 3.555000 0.100000 3.725000 0.270000 ;
        RECT 3.555000 7.740000 3.725000 7.910000 ;
        RECT 3.915000 0.100000 4.085000 0.270000 ;
        RECT 3.915000 7.740000 4.085000 7.910000 ;
        RECT 4.275000 0.100000 4.445000 0.270000 ;
        RECT 4.275000 7.740000 4.445000 7.910000 ;
        RECT 4.635000 0.100000 4.805000 0.270000 ;
        RECT 4.635000 7.740000 4.805000 7.910000 ;
        RECT 4.995000 0.100000 5.165000 0.270000 ;
        RECT 4.995000 7.740000 5.165000 7.910000 ;
        RECT 5.355000 0.100000 5.525000 0.270000 ;
        RECT 5.355000 7.740000 5.525000 7.910000 ;
        RECT 5.715000 0.100000 5.885000 0.270000 ;
        RECT 5.715000 7.740000 5.885000 7.910000 ;
        RECT 6.075000 0.100000 6.245000 0.270000 ;
        RECT 6.075000 7.740000 6.245000 7.910000 ;
        RECT 6.435000 0.100000 6.605000 0.270000 ;
        RECT 6.435000 7.740000 6.605000 7.910000 ;
        RECT 6.795000 0.100000 6.965000 0.270000 ;
        RECT 6.795000 7.740000 6.965000 7.910000 ;
        RECT 7.155000 0.100000 7.325000 0.270000 ;
        RECT 7.155000 7.740000 7.325000 7.910000 ;
        RECT 7.515000 0.100000 7.685000 0.270000 ;
        RECT 7.515000 7.740000 7.685000 7.910000 ;
        RECT 7.875000 0.100000 8.045000 0.270000 ;
        RECT 7.875000 7.740000 8.045000 7.910000 ;
        RECT 8.235000 0.100000 8.405000 0.270000 ;
        RECT 8.235000 7.740000 8.405000 7.910000 ;
        RECT 8.595000 0.100000 8.765000 0.270000 ;
        RECT 8.595000 7.740000 8.765000 7.910000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.975000 0.000000 8.825000 0.330000 ;
        RECT 0.975000 7.680000 8.825000 8.010000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  11.91120 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.525000 9.750000 2.125000 ;
        RECT 0.050000 5.885000 9.750000 7.485000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  2.056100 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.525000 0.470000 7.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.330000 0.525000 9.620000 7.485000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.440000 0.410000 7.570000 ;
      RECT 0.915000 0.440000 1.085000 7.570000 ;
      RECT 1.695000 0.440000 1.865000 7.570000 ;
      RECT 2.475000 0.440000 2.645000 7.570000 ;
      RECT 3.255000 0.440000 3.425000 7.570000 ;
      RECT 4.035000 0.440000 4.205000 7.570000 ;
      RECT 4.815000 0.440000 4.985000 7.570000 ;
      RECT 5.595000 0.440000 5.765000 7.570000 ;
      RECT 6.375000 0.440000 6.545000 7.570000 ;
      RECT 7.155000 0.440000 7.325000 7.570000 ;
      RECT 7.935000 0.440000 8.105000 7.570000 ;
      RECT 8.715000 0.440000 8.885000 7.570000 ;
      RECT 9.390000 0.440000 9.560000 7.570000 ;
    LAYER mcon ;
      RECT 0.240000 0.680000 0.410000 0.850000 ;
      RECT 0.240000 1.040000 0.410000 1.210000 ;
      RECT 0.240000 1.400000 0.410000 1.570000 ;
      RECT 0.240000 1.760000 0.410000 1.930000 ;
      RECT 0.240000 2.120000 0.410000 2.290000 ;
      RECT 0.240000 2.480000 0.410000 2.650000 ;
      RECT 0.240000 2.840000 0.410000 3.010000 ;
      RECT 0.240000 3.200000 0.410000 3.370000 ;
      RECT 0.240000 3.560000 0.410000 3.730000 ;
      RECT 0.240000 3.920000 0.410000 4.090000 ;
      RECT 0.240000 4.280000 0.410000 4.450000 ;
      RECT 0.240000 4.640000 0.410000 4.810000 ;
      RECT 0.240000 5.000000 0.410000 5.170000 ;
      RECT 0.240000 5.360000 0.410000 5.530000 ;
      RECT 0.240000 5.720000 0.410000 5.890000 ;
      RECT 0.240000 6.080000 0.410000 6.250000 ;
      RECT 0.240000 6.440000 0.410000 6.610000 ;
      RECT 0.240000 6.800000 0.410000 6.970000 ;
      RECT 0.240000 7.160000 0.410000 7.330000 ;
      RECT 0.915000 0.680000 1.085000 0.850000 ;
      RECT 0.915000 1.040000 1.085000 1.210000 ;
      RECT 0.915000 1.400000 1.085000 1.570000 ;
      RECT 0.915000 1.760000 1.085000 1.930000 ;
      RECT 0.915000 2.120000 1.085000 2.290000 ;
      RECT 0.915000 2.480000 1.085000 2.650000 ;
      RECT 0.915000 2.840000 1.085000 3.010000 ;
      RECT 0.915000 3.200000 1.085000 3.370000 ;
      RECT 0.915000 3.560000 1.085000 3.730000 ;
      RECT 0.915000 3.920000 1.085000 4.090000 ;
      RECT 0.915000 4.280000 1.085000 4.450000 ;
      RECT 0.915000 4.640000 1.085000 4.810000 ;
      RECT 0.915000 5.000000 1.085000 5.170000 ;
      RECT 0.915000 5.360000 1.085000 5.530000 ;
      RECT 0.915000 5.720000 1.085000 5.890000 ;
      RECT 0.915000 6.080000 1.085000 6.250000 ;
      RECT 0.915000 6.440000 1.085000 6.610000 ;
      RECT 0.915000 6.800000 1.085000 6.970000 ;
      RECT 0.915000 7.160000 1.085000 7.330000 ;
      RECT 1.695000 0.680000 1.865000 0.850000 ;
      RECT 1.695000 1.040000 1.865000 1.210000 ;
      RECT 1.695000 1.400000 1.865000 1.570000 ;
      RECT 1.695000 1.760000 1.865000 1.930000 ;
      RECT 1.695000 2.120000 1.865000 2.290000 ;
      RECT 1.695000 2.480000 1.865000 2.650000 ;
      RECT 1.695000 2.840000 1.865000 3.010000 ;
      RECT 1.695000 3.200000 1.865000 3.370000 ;
      RECT 1.695000 3.560000 1.865000 3.730000 ;
      RECT 1.695000 3.920000 1.865000 4.090000 ;
      RECT 1.695000 4.280000 1.865000 4.450000 ;
      RECT 1.695000 4.640000 1.865000 4.810000 ;
      RECT 1.695000 5.000000 1.865000 5.170000 ;
      RECT 1.695000 5.360000 1.865000 5.530000 ;
      RECT 1.695000 5.720000 1.865000 5.890000 ;
      RECT 1.695000 6.080000 1.865000 6.250000 ;
      RECT 1.695000 6.440000 1.865000 6.610000 ;
      RECT 1.695000 6.800000 1.865000 6.970000 ;
      RECT 1.695000 7.160000 1.865000 7.330000 ;
      RECT 2.475000 0.680000 2.645000 0.850000 ;
      RECT 2.475000 1.040000 2.645000 1.210000 ;
      RECT 2.475000 1.400000 2.645000 1.570000 ;
      RECT 2.475000 1.760000 2.645000 1.930000 ;
      RECT 2.475000 2.120000 2.645000 2.290000 ;
      RECT 2.475000 2.480000 2.645000 2.650000 ;
      RECT 2.475000 2.840000 2.645000 3.010000 ;
      RECT 2.475000 3.200000 2.645000 3.370000 ;
      RECT 2.475000 3.560000 2.645000 3.730000 ;
      RECT 2.475000 3.920000 2.645000 4.090000 ;
      RECT 2.475000 4.280000 2.645000 4.450000 ;
      RECT 2.475000 4.640000 2.645000 4.810000 ;
      RECT 2.475000 5.000000 2.645000 5.170000 ;
      RECT 2.475000 5.360000 2.645000 5.530000 ;
      RECT 2.475000 5.720000 2.645000 5.890000 ;
      RECT 2.475000 6.080000 2.645000 6.250000 ;
      RECT 2.475000 6.440000 2.645000 6.610000 ;
      RECT 2.475000 6.800000 2.645000 6.970000 ;
      RECT 2.475000 7.160000 2.645000 7.330000 ;
      RECT 3.255000 0.680000 3.425000 0.850000 ;
      RECT 3.255000 1.040000 3.425000 1.210000 ;
      RECT 3.255000 1.400000 3.425000 1.570000 ;
      RECT 3.255000 1.760000 3.425000 1.930000 ;
      RECT 3.255000 2.120000 3.425000 2.290000 ;
      RECT 3.255000 2.480000 3.425000 2.650000 ;
      RECT 3.255000 2.840000 3.425000 3.010000 ;
      RECT 3.255000 3.200000 3.425000 3.370000 ;
      RECT 3.255000 3.560000 3.425000 3.730000 ;
      RECT 3.255000 3.920000 3.425000 4.090000 ;
      RECT 3.255000 4.280000 3.425000 4.450000 ;
      RECT 3.255000 4.640000 3.425000 4.810000 ;
      RECT 3.255000 5.000000 3.425000 5.170000 ;
      RECT 3.255000 5.360000 3.425000 5.530000 ;
      RECT 3.255000 5.720000 3.425000 5.890000 ;
      RECT 3.255000 6.080000 3.425000 6.250000 ;
      RECT 3.255000 6.440000 3.425000 6.610000 ;
      RECT 3.255000 6.800000 3.425000 6.970000 ;
      RECT 3.255000 7.160000 3.425000 7.330000 ;
      RECT 4.035000 0.680000 4.205000 0.850000 ;
      RECT 4.035000 1.040000 4.205000 1.210000 ;
      RECT 4.035000 1.400000 4.205000 1.570000 ;
      RECT 4.035000 1.760000 4.205000 1.930000 ;
      RECT 4.035000 2.120000 4.205000 2.290000 ;
      RECT 4.035000 2.480000 4.205000 2.650000 ;
      RECT 4.035000 2.840000 4.205000 3.010000 ;
      RECT 4.035000 3.200000 4.205000 3.370000 ;
      RECT 4.035000 3.560000 4.205000 3.730000 ;
      RECT 4.035000 3.920000 4.205000 4.090000 ;
      RECT 4.035000 4.280000 4.205000 4.450000 ;
      RECT 4.035000 4.640000 4.205000 4.810000 ;
      RECT 4.035000 5.000000 4.205000 5.170000 ;
      RECT 4.035000 5.360000 4.205000 5.530000 ;
      RECT 4.035000 5.720000 4.205000 5.890000 ;
      RECT 4.035000 6.080000 4.205000 6.250000 ;
      RECT 4.035000 6.440000 4.205000 6.610000 ;
      RECT 4.035000 6.800000 4.205000 6.970000 ;
      RECT 4.035000 7.160000 4.205000 7.330000 ;
      RECT 4.815000 0.680000 4.985000 0.850000 ;
      RECT 4.815000 1.040000 4.985000 1.210000 ;
      RECT 4.815000 1.400000 4.985000 1.570000 ;
      RECT 4.815000 1.760000 4.985000 1.930000 ;
      RECT 4.815000 2.120000 4.985000 2.290000 ;
      RECT 4.815000 2.480000 4.985000 2.650000 ;
      RECT 4.815000 2.840000 4.985000 3.010000 ;
      RECT 4.815000 3.200000 4.985000 3.370000 ;
      RECT 4.815000 3.560000 4.985000 3.730000 ;
      RECT 4.815000 3.920000 4.985000 4.090000 ;
      RECT 4.815000 4.280000 4.985000 4.450000 ;
      RECT 4.815000 4.640000 4.985000 4.810000 ;
      RECT 4.815000 5.000000 4.985000 5.170000 ;
      RECT 4.815000 5.360000 4.985000 5.530000 ;
      RECT 4.815000 5.720000 4.985000 5.890000 ;
      RECT 4.815000 6.080000 4.985000 6.250000 ;
      RECT 4.815000 6.440000 4.985000 6.610000 ;
      RECT 4.815000 6.800000 4.985000 6.970000 ;
      RECT 4.815000 7.160000 4.985000 7.330000 ;
      RECT 5.595000 0.680000 5.765000 0.850000 ;
      RECT 5.595000 1.040000 5.765000 1.210000 ;
      RECT 5.595000 1.400000 5.765000 1.570000 ;
      RECT 5.595000 1.760000 5.765000 1.930000 ;
      RECT 5.595000 2.120000 5.765000 2.290000 ;
      RECT 5.595000 2.480000 5.765000 2.650000 ;
      RECT 5.595000 2.840000 5.765000 3.010000 ;
      RECT 5.595000 3.200000 5.765000 3.370000 ;
      RECT 5.595000 3.560000 5.765000 3.730000 ;
      RECT 5.595000 3.920000 5.765000 4.090000 ;
      RECT 5.595000 4.280000 5.765000 4.450000 ;
      RECT 5.595000 4.640000 5.765000 4.810000 ;
      RECT 5.595000 5.000000 5.765000 5.170000 ;
      RECT 5.595000 5.360000 5.765000 5.530000 ;
      RECT 5.595000 5.720000 5.765000 5.890000 ;
      RECT 5.595000 6.080000 5.765000 6.250000 ;
      RECT 5.595000 6.440000 5.765000 6.610000 ;
      RECT 5.595000 6.800000 5.765000 6.970000 ;
      RECT 5.595000 7.160000 5.765000 7.330000 ;
      RECT 6.375000 0.680000 6.545000 0.850000 ;
      RECT 6.375000 1.040000 6.545000 1.210000 ;
      RECT 6.375000 1.400000 6.545000 1.570000 ;
      RECT 6.375000 1.760000 6.545000 1.930000 ;
      RECT 6.375000 2.120000 6.545000 2.290000 ;
      RECT 6.375000 2.480000 6.545000 2.650000 ;
      RECT 6.375000 2.840000 6.545000 3.010000 ;
      RECT 6.375000 3.200000 6.545000 3.370000 ;
      RECT 6.375000 3.560000 6.545000 3.730000 ;
      RECT 6.375000 3.920000 6.545000 4.090000 ;
      RECT 6.375000 4.280000 6.545000 4.450000 ;
      RECT 6.375000 4.640000 6.545000 4.810000 ;
      RECT 6.375000 5.000000 6.545000 5.170000 ;
      RECT 6.375000 5.360000 6.545000 5.530000 ;
      RECT 6.375000 5.720000 6.545000 5.890000 ;
      RECT 6.375000 6.080000 6.545000 6.250000 ;
      RECT 6.375000 6.440000 6.545000 6.610000 ;
      RECT 6.375000 6.800000 6.545000 6.970000 ;
      RECT 6.375000 7.160000 6.545000 7.330000 ;
      RECT 7.155000 0.680000 7.325000 0.850000 ;
      RECT 7.155000 1.040000 7.325000 1.210000 ;
      RECT 7.155000 1.400000 7.325000 1.570000 ;
      RECT 7.155000 1.760000 7.325000 1.930000 ;
      RECT 7.155000 2.120000 7.325000 2.290000 ;
      RECT 7.155000 2.480000 7.325000 2.650000 ;
      RECT 7.155000 2.840000 7.325000 3.010000 ;
      RECT 7.155000 3.200000 7.325000 3.370000 ;
      RECT 7.155000 3.560000 7.325000 3.730000 ;
      RECT 7.155000 3.920000 7.325000 4.090000 ;
      RECT 7.155000 4.280000 7.325000 4.450000 ;
      RECT 7.155000 4.640000 7.325000 4.810000 ;
      RECT 7.155000 5.000000 7.325000 5.170000 ;
      RECT 7.155000 5.360000 7.325000 5.530000 ;
      RECT 7.155000 5.720000 7.325000 5.890000 ;
      RECT 7.155000 6.080000 7.325000 6.250000 ;
      RECT 7.155000 6.440000 7.325000 6.610000 ;
      RECT 7.155000 6.800000 7.325000 6.970000 ;
      RECT 7.155000 7.160000 7.325000 7.330000 ;
      RECT 7.935000 0.680000 8.105000 0.850000 ;
      RECT 7.935000 1.040000 8.105000 1.210000 ;
      RECT 7.935000 1.400000 8.105000 1.570000 ;
      RECT 7.935000 1.760000 8.105000 1.930000 ;
      RECT 7.935000 2.120000 8.105000 2.290000 ;
      RECT 7.935000 2.480000 8.105000 2.650000 ;
      RECT 7.935000 2.840000 8.105000 3.010000 ;
      RECT 7.935000 3.200000 8.105000 3.370000 ;
      RECT 7.935000 3.560000 8.105000 3.730000 ;
      RECT 7.935000 3.920000 8.105000 4.090000 ;
      RECT 7.935000 4.280000 8.105000 4.450000 ;
      RECT 7.935000 4.640000 8.105000 4.810000 ;
      RECT 7.935000 5.000000 8.105000 5.170000 ;
      RECT 7.935000 5.360000 8.105000 5.530000 ;
      RECT 7.935000 5.720000 8.105000 5.890000 ;
      RECT 7.935000 6.080000 8.105000 6.250000 ;
      RECT 7.935000 6.440000 8.105000 6.610000 ;
      RECT 7.935000 6.800000 8.105000 6.970000 ;
      RECT 7.935000 7.160000 8.105000 7.330000 ;
      RECT 8.715000 0.680000 8.885000 0.850000 ;
      RECT 8.715000 1.040000 8.885000 1.210000 ;
      RECT 8.715000 1.400000 8.885000 1.570000 ;
      RECT 8.715000 1.760000 8.885000 1.930000 ;
      RECT 8.715000 2.120000 8.885000 2.290000 ;
      RECT 8.715000 2.480000 8.885000 2.650000 ;
      RECT 8.715000 2.840000 8.885000 3.010000 ;
      RECT 8.715000 3.200000 8.885000 3.370000 ;
      RECT 8.715000 3.560000 8.885000 3.730000 ;
      RECT 8.715000 3.920000 8.885000 4.090000 ;
      RECT 8.715000 4.280000 8.885000 4.450000 ;
      RECT 8.715000 4.640000 8.885000 4.810000 ;
      RECT 8.715000 5.000000 8.885000 5.170000 ;
      RECT 8.715000 5.360000 8.885000 5.530000 ;
      RECT 8.715000 5.720000 8.885000 5.890000 ;
      RECT 8.715000 6.080000 8.885000 6.250000 ;
      RECT 8.715000 6.440000 8.885000 6.610000 ;
      RECT 8.715000 6.800000 8.885000 6.970000 ;
      RECT 8.715000 7.160000 8.885000 7.330000 ;
      RECT 9.390000 0.680000 9.560000 0.850000 ;
      RECT 9.390000 1.040000 9.560000 1.210000 ;
      RECT 9.390000 1.400000 9.560000 1.570000 ;
      RECT 9.390000 1.760000 9.560000 1.930000 ;
      RECT 9.390000 2.120000 9.560000 2.290000 ;
      RECT 9.390000 2.480000 9.560000 2.650000 ;
      RECT 9.390000 2.840000 9.560000 3.010000 ;
      RECT 9.390000 3.200000 9.560000 3.370000 ;
      RECT 9.390000 3.560000 9.560000 3.730000 ;
      RECT 9.390000 3.920000 9.560000 4.090000 ;
      RECT 9.390000 4.280000 9.560000 4.450000 ;
      RECT 9.390000 4.640000 9.560000 4.810000 ;
      RECT 9.390000 5.000000 9.560000 5.170000 ;
      RECT 9.390000 5.360000 9.560000 5.530000 ;
      RECT 9.390000 5.720000 9.560000 5.890000 ;
      RECT 9.390000 6.080000 9.560000 6.250000 ;
      RECT 9.390000 6.440000 9.560000 6.610000 ;
      RECT 9.390000 6.800000 9.560000 6.970000 ;
      RECT 9.390000 7.160000 9.560000 7.330000 ;
    LAYER met1 ;
      RECT 0.870000 0.525000 1.130000 7.485000 ;
      RECT 1.650000 0.525000 1.910000 7.485000 ;
      RECT 2.430000 0.525000 2.690000 7.485000 ;
      RECT 3.210000 0.525000 3.470000 7.485000 ;
      RECT 3.990000 0.525000 4.250000 7.485000 ;
      RECT 4.770000 0.525000 5.030000 7.485000 ;
      RECT 5.550000 0.525000 5.810000 7.485000 ;
      RECT 6.330000 0.525000 6.590000 7.485000 ;
      RECT 7.110000 0.525000 7.370000 7.485000 ;
      RECT 7.890000 0.525000 8.150000 7.485000 ;
      RECT 8.670000 0.525000 8.930000 7.485000 ;
    LAYER via ;
      RECT 0.870000 0.555000 1.130000 0.815000 ;
      RECT 0.870000 0.875000 1.130000 1.135000 ;
      RECT 0.870000 1.195000 1.130000 1.455000 ;
      RECT 0.870000 1.515000 1.130000 1.775000 ;
      RECT 0.870000 1.835000 1.130000 2.095000 ;
      RECT 0.870000 5.915000 1.130000 6.175000 ;
      RECT 0.870000 6.235000 1.130000 6.495000 ;
      RECT 0.870000 6.555000 1.130000 6.815000 ;
      RECT 0.870000 6.875000 1.130000 7.135000 ;
      RECT 0.870000 7.195000 1.130000 7.455000 ;
      RECT 1.650000 2.435000 1.910000 2.695000 ;
      RECT 1.650000 2.755000 1.910000 3.015000 ;
      RECT 1.650000 3.075000 1.910000 3.335000 ;
      RECT 1.650000 3.395000 1.910000 3.655000 ;
      RECT 1.650000 3.715000 1.910000 3.975000 ;
      RECT 1.650000 4.035000 1.910000 4.295000 ;
      RECT 1.650000 4.355000 1.910000 4.615000 ;
      RECT 1.650000 4.675000 1.910000 4.935000 ;
      RECT 1.650000 4.995000 1.910000 5.255000 ;
      RECT 1.650000 5.315000 1.910000 5.575000 ;
      RECT 2.430000 0.555000 2.690000 0.815000 ;
      RECT 2.430000 0.875000 2.690000 1.135000 ;
      RECT 2.430000 1.195000 2.690000 1.455000 ;
      RECT 2.430000 1.515000 2.690000 1.775000 ;
      RECT 2.430000 1.835000 2.690000 2.095000 ;
      RECT 2.430000 5.915000 2.690000 6.175000 ;
      RECT 2.430000 6.235000 2.690000 6.495000 ;
      RECT 2.430000 6.555000 2.690000 6.815000 ;
      RECT 2.430000 6.875000 2.690000 7.135000 ;
      RECT 2.430000 7.195000 2.690000 7.455000 ;
      RECT 3.210000 2.435000 3.470000 2.695000 ;
      RECT 3.210000 2.755000 3.470000 3.015000 ;
      RECT 3.210000 3.075000 3.470000 3.335000 ;
      RECT 3.210000 3.395000 3.470000 3.655000 ;
      RECT 3.210000 3.715000 3.470000 3.975000 ;
      RECT 3.210000 4.035000 3.470000 4.295000 ;
      RECT 3.210000 4.355000 3.470000 4.615000 ;
      RECT 3.210000 4.675000 3.470000 4.935000 ;
      RECT 3.210000 4.995000 3.470000 5.255000 ;
      RECT 3.210000 5.315000 3.470000 5.575000 ;
      RECT 3.990000 0.555000 4.250000 0.815000 ;
      RECT 3.990000 0.875000 4.250000 1.135000 ;
      RECT 3.990000 1.195000 4.250000 1.455000 ;
      RECT 3.990000 1.515000 4.250000 1.775000 ;
      RECT 3.990000 1.835000 4.250000 2.095000 ;
      RECT 3.990000 5.915000 4.250000 6.175000 ;
      RECT 3.990000 6.235000 4.250000 6.495000 ;
      RECT 3.990000 6.555000 4.250000 6.815000 ;
      RECT 3.990000 6.875000 4.250000 7.135000 ;
      RECT 3.990000 7.195000 4.250000 7.455000 ;
      RECT 4.770000 2.435000 5.030000 2.695000 ;
      RECT 4.770000 2.755000 5.030000 3.015000 ;
      RECT 4.770000 3.075000 5.030000 3.335000 ;
      RECT 4.770000 3.395000 5.030000 3.655000 ;
      RECT 4.770000 3.715000 5.030000 3.975000 ;
      RECT 4.770000 4.035000 5.030000 4.295000 ;
      RECT 4.770000 4.355000 5.030000 4.615000 ;
      RECT 4.770000 4.675000 5.030000 4.935000 ;
      RECT 4.770000 4.995000 5.030000 5.255000 ;
      RECT 4.770000 5.315000 5.030000 5.575000 ;
      RECT 5.550000 0.555000 5.810000 0.815000 ;
      RECT 5.550000 0.875000 5.810000 1.135000 ;
      RECT 5.550000 1.195000 5.810000 1.455000 ;
      RECT 5.550000 1.515000 5.810000 1.775000 ;
      RECT 5.550000 1.835000 5.810000 2.095000 ;
      RECT 5.550000 5.915000 5.810000 6.175000 ;
      RECT 5.550000 6.235000 5.810000 6.495000 ;
      RECT 5.550000 6.555000 5.810000 6.815000 ;
      RECT 5.550000 6.875000 5.810000 7.135000 ;
      RECT 5.550000 7.195000 5.810000 7.455000 ;
      RECT 6.330000 2.435000 6.590000 2.695000 ;
      RECT 6.330000 2.755000 6.590000 3.015000 ;
      RECT 6.330000 3.075000 6.590000 3.335000 ;
      RECT 6.330000 3.395000 6.590000 3.655000 ;
      RECT 6.330000 3.715000 6.590000 3.975000 ;
      RECT 6.330000 4.035000 6.590000 4.295000 ;
      RECT 6.330000 4.355000 6.590000 4.615000 ;
      RECT 6.330000 4.675000 6.590000 4.935000 ;
      RECT 6.330000 4.995000 6.590000 5.255000 ;
      RECT 6.330000 5.315000 6.590000 5.575000 ;
      RECT 7.110000 0.555000 7.370000 0.815000 ;
      RECT 7.110000 0.875000 7.370000 1.135000 ;
      RECT 7.110000 1.195000 7.370000 1.455000 ;
      RECT 7.110000 1.515000 7.370000 1.775000 ;
      RECT 7.110000 1.835000 7.370000 2.095000 ;
      RECT 7.110000 5.915000 7.370000 6.175000 ;
      RECT 7.110000 6.235000 7.370000 6.495000 ;
      RECT 7.110000 6.555000 7.370000 6.815000 ;
      RECT 7.110000 6.875000 7.370000 7.135000 ;
      RECT 7.110000 7.195000 7.370000 7.455000 ;
      RECT 7.890000 2.435000 8.150000 2.695000 ;
      RECT 7.890000 2.755000 8.150000 3.015000 ;
      RECT 7.890000 3.075000 8.150000 3.335000 ;
      RECT 7.890000 3.395000 8.150000 3.655000 ;
      RECT 7.890000 3.715000 8.150000 3.975000 ;
      RECT 7.890000 4.035000 8.150000 4.295000 ;
      RECT 7.890000 4.355000 8.150000 4.615000 ;
      RECT 7.890000 4.675000 8.150000 4.935000 ;
      RECT 7.890000 4.995000 8.150000 5.255000 ;
      RECT 7.890000 5.315000 8.150000 5.575000 ;
      RECT 8.670000 0.555000 8.930000 0.815000 ;
      RECT 8.670000 0.875000 8.930000 1.135000 ;
      RECT 8.670000 1.195000 8.930000 1.455000 ;
      RECT 8.670000 1.515000 8.930000 1.775000 ;
      RECT 8.670000 1.835000 8.930000 2.095000 ;
      RECT 8.670000 5.915000 8.930000 6.175000 ;
      RECT 8.670000 6.235000 8.930000 6.495000 ;
      RECT 8.670000 6.555000 8.930000 6.815000 ;
      RECT 8.670000 6.875000 8.930000 7.135000 ;
      RECT 8.670000 7.195000 8.930000 7.455000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50
END LIBRARY
