module approxMult_signed8x8 (A, B, OUT);
  input  [7:0] A;
  input  [7:0] B;
  output [15:0] OUT;
  wire n0, n1, n10, n11, n12, n13, n14, n15, n2, n3, n4, n5, n6, n7, n8, n9, v0_0, v100_0, v101_0, v102_0, v103_0, v104_0, v105_0, v106_0, v107_0, v108_0, v109_0, v10_0, v110_0, v111_0, v112_0, v113_0, v114_0, v115_0, v116_0, v117_0, v118_0, v119_0, v11_0, v120_0, v121_0, v122_0, v123_0, v124_0, v125_0, v126_0, v127_0, v128_0, v129_0, v12_0, v130_0, v131_0, v132_0, v133_0, v134_0, v135_0, v136_0, v137_0, v138_0, v139_0, v13_0, v140_0, v141_0, v142_0, v143_0, v144_0, v145_0, v146_0, v147_0, v148_0, v149_0, v14_0, v150_0, v151_0, v152_0, v153_0, v154_0, v155_0, v156_0, v157_0, v158_0, v159_0, v15_0, v160_0, v161_0, v162_0, v163_0, v164_0, v165_0, v166_0, v167_0, v168_0, v169_0, v16_0, v170_0, v171_0, v172_0, v173_0, v174_0, v175_0, v176_0, v177_0, v178_0, v179_0, v17_0, v180_0, v181_0, v182_0, v183_0, v184_0, v185_0, v186_0, v187_0, v188_0, v189_0, v18_0, v190_0, v191_0, v192_0, v193_0, v194_0, v195_0, v196_0, v197_0, v198_0, v199_0, v19_0, v1_0, v200_0, v201_0, v202_0, v203_0, v204_0, v205_0, v206_0, v207_0, v208_0, v209_0, v20_0, v210_0, v211_0, v212_0, v213_0, v214_0, v215_0, v216_0, v217_0, v218_0, v219_0, v21_0, v220_0, v221_0, v222_0, v223_0, v224_0, v225_0, v226_0, v227_0, v228_0, v229_0, v22_0, v230_0, v231_0, v232_0, v233_0, v234_0, v235_0, v236_0, v237_0, v238_0, v239_0, v23_0, v240_0, v241_0, v242_0, v243_0, v244_0, v245_0, v246_0, v247_0, v248_0, v249_0, v24_0, v250_0, v251_0, v252_0, v253_0, v254_0, v255_0, v256_0, v257_0, v258_0, v259_0, v25_0, v260_0, v261_0, v262_0, v263_0, v264_0, v265_0, v266_0, v267_0, v268_0, v269_0, v26_0, v270_0, v271_0, v272_0, v273_0, v274_0, v275_0, v276_0, v277_0, v278_0, v279_0, v27_0, v280_0, v281_0, v282_0, v283_0, v284_0, v285_0, v286_0, v287_0, v288_0, v289_0, v28_0, v290_0, v291_0, v292_0, v293_0, v294_0, v295_0, v296_0, v297_0, v298_0, v299_0, v29_0, v2_0, v300_0, v301_0, v302_0, v303_0, v304_0, v305_0, v306_0, v307_0, v308_0, v309_0, v30_0, v310_0, v311_0, v312_0, v313_0, v314_0, v315_0, v316_0, v317_0, v318_0, v319_0, v31_0, v320_0, v321_0, v322_0, v323_0, v324_0, v325_0, v326_0, v327_0, v328_0, v329_0, v32_0, v330_0, v331_0, v332_0, v333_0, v334_0, v335_0, v336_0, v337_0, v338_0, v339_0, v33_0, v340_0, v341_0, v342_0, v343_0, v344_0, v345_0, v346_0, v347_0, v348_0, v349_0, v34_0, v350_0, v351_0, v352_0, v353_0, v354_0, v355_0, v356_0, v357_0, v358_0, v359_0, v35_0, v360_0, v361_0, v362_0, v363_0, v364_0, v365_0, v366_0, v367_0, v368_0, v369_0, v36_0, v370_0, v371_0, v372_0, v373_0, v374_0, v375_0, v376_0, v377_0, v378_0, v379_0, v37_0, v380_0, v381_0, v382_0, v383_0, v384_0, v385_0, v386_0, v387_0, v388_0, v389_0, v38_0, v390_0, v391_0, v392_0, v393_0, v394_0, v395_0, v396_0, v397_0, v398_0, v399_0, v39_0, v3_0, v40_0, v41_0, v42_0, v43_0, v44_0, v45_0, v46_0, v47_0, v48_0, v49_0, v4_0, v50_0, v51_0, v52_0, v53_0, v54_0, v55_0, v56_0, v57_0, v58_0, v59_0, v5_0, v60_0, v61_0, v62_0, v63_0, v64_0, v65_0, v66_0, v67_0, v68_0, v69_0, v6_0, v70_0, v71_0, v72_0, v73_0, v74_0, v75_0, v76_0, v77_0, v78_0, v79_0, v7_0, v80_0, v81_0, v82_0, v83_0, v84_0, v85_0, v86_0, v87_0, v88_0, v89_0, v8_0, v90_0, v91_0, v92_0, v93_0, v94_0, v95_0, v96_0, v97_0, v98_0, v99_0, v9_0;

  // Map n0..n7 to A[0..7], n8..n15 to B[0..7]
  assign n0 = A[0];
  assign n1 = A[1];
  assign n2 = A[2];
  assign n3 = A[3];
  assign n4 = A[4];
  assign n5 = A[5];
  assign n6 = A[6];
  assign n7 = A[7];
  assign n8 = B[0];
  assign n9 = B[1];
  assign n10 = B[2];
  assign n11 = B[3];
  assign n12 = B[4];
  assign n13 = B[5];
  assign n14 = B[6];
  assign n15 = B[7];

  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0001_ (
    .A1(n12),
    .A2(n1),
    .ZN(v0_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0002_ (
    .I(v0_0),
    .ZN(v1_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0003_ (
    .I(n2),
    .ZN(v2_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0004_ (
    .A1(n8),
    .A2(n4),
    .ZN(v3_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0005_ (
    .A1(n2),
    .A2(n11),
    .ZN(v4_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0006_ (
    .I(v4_0),
    .ZN(v5_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0007_ (
    .A1(v1_0),
    .A2(v5_0),
    .ZN(v6_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0008_ (
    .A1(v0_0),
    .A2(v4_0),
    .ZN(v7_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0009_ (
    .I(v7_0),
    .ZN(v8_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0010_ (
    .A1(n13),
    .A2(n0),
    .ZN(v9_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0011_ (
    .A1(v8_0),
    .A2(v9_0),
    .Z(v10_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0012_ (
    .A1(n10),
    .A2(n3),
    .ZN(v11_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0013_ (
    .A1(n5),
    .A2(n9),
    .ZN(v12_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0014_ (
    .A1(v3_0),
    .A2(v12_0),
    .Z(v13_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0015_ (
    .I(v3_0),
    .ZN(v14_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0016_ (
    .I(v14_0),
    .ZN(v15_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0017_ (
    .A1(v8_0),
    .A2(v15_0),
    .Z(v16_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0018_ (
    .I(v16_0),
    .ZN(v17_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0019_ (
    .I(v17_0),
    .ZN(v18_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0020_ (
    .I(v18_0),
    .ZN(v19_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0021_ (
    .A1(v15_0),
    .A2(v8_0),
    .Z(v20_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0022_ (
    .I(v20_0),
    .ZN(v21_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0023_ (
    .A1(n3),
    .A2(n12),
    .ZN(v22_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0024_ (
    .I(v22_0),
    .ZN(v23_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0025_ (
    .A1(v23_0),
    .A2(v5_0),
    .ZN(v24_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0026_ (
    .A1(n2),
    .A2(n12),
    .ZN(v25_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0027_ (
    .A1(n3),
    .A2(n11),
    .ZN(v26_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0028_ (
    .A1(v25_0),
    .A2(v26_0),
    .ZN(v27_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0029_ (
    .A1(v24_0),
    .A2(v27_0),
    .ZN(v28_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0030_ (
    .A1(n1),
    .A2(n13),
    .ZN(v29_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0031_ (
    .A1(v28_0),
    .A2(v29_0),
    .Z(v30_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0032_ (
    .A1(v28_0),
    .A2(v29_0),
    .ZN(v31_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0033_ (
    .A1(v30_0),
    .A2(v31_0),
    .ZN(v32_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0034_ (
    .A1(v11_0),
    .A2(v13_0),
    .Z(v33_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0035_ (
    .A1(n8),
    .A2(n6),
    .ZN(v34_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0036_ (
    .A1(v12_0),
    .A2(v34_0),
    .ZN(v35_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0037_ (
    .A1(n4),
    .A2(n10),
    .ZN(v36_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0038_ (
    .I(v36_0),
    .ZN(v37_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0039_ (
    .A1(v35_0),
    .A2(v37_0),
    .ZN(v38_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0040_ (
    .A1(n5),
    .A2(n8),
    .Z(v39_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0041_ (
    .A1(n9),
    .A2(n6),
    .Z(v40_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0042_ (
    .A1(v39_0),
    .A2(v40_0),
    .ZN(v41_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0043_ (
    .A1(v41_0),
    .A2(v35_0),
    .ZN(v42_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0044_ (
    .A1(v42_0),
    .A2(v36_0),
    .ZN(v43_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0045_ (
    .A1(v38_0),
    .A2(v43_0),
    .ZN(v44_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0046_ (
    .A1(v33_0),
    .A2(v44_0),
    .ZN(v45_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0047_ (
    .A1(v36_0),
    .A2(v42_0),
    .Z(v46_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0048_ (
    .A1(v11_0),
    .A2(v13_0),
    .ZN(v47_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0049_ (
    .A1(v46_0),
    .A2(v47_0),
    .ZN(v48_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0050_ (
    .A1(v45_0),
    .A2(v48_0),
    .ZN(v49_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0051_ (
    .A1(v32_0),
    .A2(v49_0),
    .Z(v50_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0052_ (
    .A1(v21_0),
    .A2(v50_0),
    .Z(v51_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0053_ (
    .A1(n0),
    .A2(n14),
    .ZN(v52_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0054_ (
    .I(v52_0),
    .ZN(v53_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0055_ (
    .A1(v10_0),
    .A2(v6_0),
    .ZN(v54_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0056_ (
    .A1(v53_0),
    .A2(v54_0),
    .Z(v55_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0057_ (
    .A1(v51_0),
    .A2(v55_0),
    .ZN(v56_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0058_ (
    .A1(v50_0),
    .A2(v21_0),
    .ZN(v57_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0059_ (
    .I(v51_0),
    .ZN(v58_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0060_ (
    .I(v55_0),
    .ZN(v59_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0061_ (
    .A1(v58_0),
    .A2(v59_0),
    .ZN(v60_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0062_ (
    .A1(v56_0),
    .A2(v60_0),
    .ZN(v61_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0063_ (
    .A1(v19_0),
    .A2(v61_0),
    .ZN(v62_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0064_ (
    .I(v61_0),
    .ZN(v63_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0065_ (
    .A1(v63_0),
    .A2(v18_0),
    .ZN(v64_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0066_ (
    .A1(v62_0),
    .A2(v64_0),
    .ZN(v65_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0067_ (
    .I(v65_0),
    .ZN(v66_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0068_ (
    .A1(v56_0),
    .A2(v57_0),
    .ZN(v67_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0069_ (
    .A1(v30_0),
    .A2(v24_0),
    .ZN(v68_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0070_ (
    .A1(n1),
    .A2(n14),
    .ZN(v69_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0071_ (
    .A1(n2),
    .A2(n13),
    .ZN(v70_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0072_ (
    .A1(v69_0),
    .A2(v70_0),
    .Z(v71_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0073_ (
    .I(v71_0),
    .ZN(v72_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0074_ (
    .I(n15),
    .ZN(v73_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0075_ (
    .A1(v73_0),
    .A2(n0),
    .Z(v74_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0076_ (
    .A1(v72_0),
    .A2(v74_0),
    .Z(v75_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0077_ (
    .A1(v72_0),
    .A2(v74_0),
    .ZN(v76_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0078_ (
    .A1(v75_0),
    .A2(v76_0),
    .ZN(v77_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0079_ (
    .A1(v68_0),
    .A2(v77_0),
    .Z(v78_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0080_ (
    .I(v32_0),
    .ZN(v79_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0081_ (
    .A1(v45_0),
    .A2(v79_0),
    .ZN(v80_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0082_ (
    .A1(v80_0),
    .A2(v48_0),
    .Z(v81_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0083_ (
    .A1(n8),
    .A2(n7),
    .ZN(v82_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0084_ (
    .A1(v73_0),
    .A2(v82_0),
    .Z(v83_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0085_ (
    .A1(v83_0),
    .A2(v40_0),
    .ZN(v84_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0086_ (
    .A1(n8),
    .A2(n7),
    .Z(v85_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0087_ (
    .A1(v85_0),
    .A2(n15),
    .ZN(v86_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0088_ (
    .I(v83_0),
    .ZN(v87_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0089_ (
    .I(v40_0),
    .ZN(v88_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0090_ (
    .A1(v87_0),
    .A2(v88_0),
    .ZN(v89_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0091_ (
    .A1(v84_0),
    .A2(v89_0),
    .ZN(v90_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0092_ (
    .A1(v38_0),
    .A2(v41_0),
    .ZN(v91_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0093_ (
    .A1(v90_0),
    .A2(v91_0),
    .Z(v92_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0094_ (
    .A1(n5),
    .A2(n11),
    .ZN(v93_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0095_ (
    .A1(v36_0),
    .A2(v93_0),
    .Z(v94_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0096_ (
    .A1(n4),
    .A2(n11),
    .ZN(v95_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0097_ (
    .A1(n5),
    .A2(n10),
    .ZN(v96_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0098_ (
    .A1(v95_0),
    .A2(v96_0),
    .ZN(v97_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0099_ (
    .A1(v94_0),
    .A2(v97_0),
    .ZN(v98_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0100_ (
    .A1(v98_0),
    .A2(v22_0),
    .Z(v99_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0101_ (
    .A1(v98_0),
    .A2(v22_0),
    .ZN(v100_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0102_ (
    .I(v81_0),
    .ZN(v101_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0103_ (
    .A1(v99_0),
    .A2(v100_0),
    .ZN(v102_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0104_ (
    .A1(v92_0),
    .A2(v102_0),
    .Z(v103_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0105_ (
    .A1(v92_0),
    .A2(v102_0),
    .ZN(v104_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0106_ (
    .A1(v103_0),
    .A2(v104_0),
    .ZN(v105_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0107_ (
    .A1(v81_0),
    .A2(v105_0),
    .ZN(v106_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0108_ (
    .A1(v102_0),
    .A2(v92_0),
    .Z(v107_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0109_ (
    .A1(v107_0),
    .A2(v101_0),
    .ZN(v108_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0110_ (
    .A1(v106_0),
    .A2(v108_0),
    .ZN(v109_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0111_ (
    .A1(v78_0),
    .A2(v109_0),
    .Z(v110_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0112_ (
    .A1(v67_0),
    .A2(v110_0),
    .Z(v111_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0113_ (
    .A1(v54_0),
    .A2(v53_0),
    .ZN(v112_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0114_ (
    .I(v112_0),
    .ZN(v113_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0115_ (
    .A1(v111_0),
    .A2(v113_0),
    .ZN(v114_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0116_ (
    .A1(v110_0),
    .A2(v67_0),
    .ZN(v115_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0117_ (
    .I(v111_0),
    .ZN(v116_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0118_ (
    .A1(v116_0),
    .A2(v112_0),
    .ZN(v117_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0119_ (
    .A1(v114_0),
    .A2(v117_0),
    .ZN(v118_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0120_ (
    .A1(v64_0),
    .A2(v118_0),
    .Z(v119_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0121_ (
    .A1(v114_0),
    .A2(v115_0),
    .ZN(v120_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0122_ (
    .A1(v78_0),
    .A2(v68_0),
    .ZN(v121_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0123_ (
    .A1(v109_0),
    .A2(v78_0),
    .Z(v122_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0124_ (
    .A1(v122_0),
    .A2(v108_0),
    .ZN(v123_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0125_ (
    .A1(n5),
    .A2(n12),
    .ZN(v124_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0126_ (
    .A1(v95_0),
    .A2(v124_0),
    .Z(v125_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0127_ (
    .A1(n4),
    .A2(n12),
    .ZN(v126_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0128_ (
    .A1(v93_0),
    .A2(v126_0),
    .ZN(v127_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0129_ (
    .A1(v125_0),
    .A2(v127_0),
    .ZN(v128_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0130_ (
    .A1(n3),
    .A2(n13),
    .ZN(v129_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0131_ (
    .A1(v128_0),
    .A2(v129_0),
    .Z(v130_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0132_ (
    .A1(v128_0),
    .A2(v129_0),
    .ZN(v131_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0133_ (
    .A1(v130_0),
    .A2(v131_0),
    .ZN(v132_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0134_ (
    .A1(v84_0),
    .A2(v86_0),
    .ZN(v133_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0135_ (
    .A1(v85_0),
    .A2(n9),
    .ZN(v134_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0136_ (
    .A1(n9),
    .A2(n7),
    .ZN(v135_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0137_ (
    .A1(v82_0),
    .A2(v135_0),
    .ZN(v136_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0138_ (
    .A1(v134_0),
    .A2(v136_0),
    .ZN(v137_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0139_ (
    .A1(n10),
    .A2(n6),
    .ZN(v138_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0140_ (
    .A1(v137_0),
    .A2(v138_0),
    .Z(v139_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0141_ (
    .A1(v137_0),
    .A2(v138_0),
    .ZN(v140_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0142_ (
    .A1(v139_0),
    .A2(v140_0),
    .ZN(v141_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0143_ (
    .A1(v133_0),
    .A2(v141_0),
    .Z(v142_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0144_ (
    .A1(v132_0),
    .A2(v142_0),
    .Z(v143_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0145_ (
    .A1(v92_0),
    .A2(v91_0),
    .ZN(v144_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0146_ (
    .A1(v103_0),
    .A2(v144_0),
    .ZN(v145_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0147_ (
    .A1(v143_0),
    .A2(v145_0),
    .Z(v146_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0148_ (
    .A1(v143_0),
    .A2(v145_0),
    .ZN(v147_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0149_ (
    .A1(v146_0),
    .A2(v147_0),
    .ZN(v148_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0150_ (
    .A1(n2),
    .A2(n14),
    .ZN(v149_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0151_ (
    .A1(v29_0),
    .A2(v149_0),
    .Z(v150_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0152_ (
    .A1(v75_0),
    .A2(v150_0),
    .ZN(v151_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0153_ (
    .A1(v99_0),
    .A2(v94_0),
    .ZN(v152_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0154_ (
    .I(n1),
    .ZN(v153_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0155_ (
    .A1(v153_0),
    .A2(n15),
    .ZN(v154_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0156_ (
    .A1(v149_0),
    .A2(v154_0),
    .Z(v155_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0157_ (
    .A1(v152_0),
    .A2(v155_0),
    .Z(v156_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0158_ (
    .A1(v152_0),
    .A2(v155_0),
    .ZN(v157_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0159_ (
    .A1(v156_0),
    .A2(v157_0),
    .ZN(v158_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0160_ (
    .A1(v151_0),
    .A2(v158_0),
    .Z(v159_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0161_ (
    .A1(v148_0),
    .A2(v159_0),
    .Z(v160_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0162_ (
    .A1(v148_0),
    .A2(v159_0),
    .ZN(v161_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0163_ (
    .A1(v160_0),
    .A2(v161_0),
    .ZN(v162_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0164_ (
    .A1(v123_0),
    .A2(v162_0),
    .Z(v163_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0165_ (
    .A1(v121_0),
    .A2(v163_0),
    .Z(v164_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0166_ (
    .A1(v120_0),
    .A2(v164_0),
    .Z(v165_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0167_ (
    .A1(v118_0),
    .A2(v64_0),
    .Z(v166_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0168_ (
    .I(v166_0),
    .ZN(v167_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0169_ (
    .A1(v165_0),
    .A2(v167_0),
    .Z(v168_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0170_ (
    .A1(v156_0),
    .A2(v151_0),
    .ZN(v169_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0171_ (
    .A1(v169_0),
    .A2(v157_0),
    .ZN(v170_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0172_ (
    .I(v170_0),
    .ZN(v171_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0173_ (
    .A1(v160_0),
    .A2(v147_0),
    .ZN(v172_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0174_ (
    .A1(v142_0),
    .A2(v132_0),
    .Z(v173_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0175_ (
    .A1(v142_0),
    .A2(v133_0),
    .ZN(v174_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0176_ (
    .A1(v173_0),
    .A2(v174_0),
    .ZN(v175_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0177_ (
    .A1(n11),
    .A2(n6),
    .ZN(v176_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0178_ (
    .A1(v124_0),
    .A2(v176_0),
    .Z(v177_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0179_ (
    .I(v177_0),
    .ZN(v178_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0180_ (
    .A1(n4),
    .A2(n13),
    .ZN(v179_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0181_ (
    .A1(v178_0),
    .A2(v179_0),
    .Z(v180_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0182_ (
    .A1(v178_0),
    .A2(v179_0),
    .ZN(v181_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0183_ (
    .A1(v180_0),
    .A2(v181_0),
    .ZN(v182_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0184_ (
    .A1(n10),
    .A2(n7),
    .ZN(v183_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0185_ (
    .A1(v183_0),
    .A2(v137_0),
    .Z(v184_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0186_ (
    .A1(v139_0),
    .A2(v134_0),
    .ZN(v185_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0187_ (
    .A1(v184_0),
    .A2(v185_0),
    .Z(v186_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0188_ (
    .A1(v184_0),
    .A2(v185_0),
    .ZN(v187_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0189_ (
    .A1(v186_0),
    .A2(v187_0),
    .Z(v188_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0190_ (
    .A1(v182_0),
    .A2(v188_0),
    .Z(v189_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0191_ (
    .A1(v175_0),
    .A2(v189_0),
    .Z(v190_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0192_ (
    .A1(v154_0),
    .A2(v149_0),
    .Z(v191_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0193_ (
    .A1(n3),
    .A2(n14),
    .ZN(v192_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0194_ (
    .A1(v2_0),
    .A2(n15),
    .ZN(v193_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0195_ (
    .A1(v192_0),
    .A2(v193_0),
    .Z(v194_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0196_ (
    .A1(v130_0),
    .A2(v125_0),
    .ZN(v195_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0197_ (
    .A1(v194_0),
    .A2(v195_0),
    .Z(v196_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0198_ (
    .I(v196_0),
    .ZN(v197_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0199_ (
    .A1(v191_0),
    .A2(v197_0),
    .Z(v198_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0200_ (
    .I(v198_0),
    .ZN(v199_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0201_ (
    .A1(v190_0),
    .A2(v199_0),
    .Z(v200_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0202_ (
    .A1(v190_0),
    .A2(v199_0),
    .ZN(v201_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0203_ (
    .A1(v200_0),
    .A2(v201_0),
    .ZN(v202_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0204_ (
    .A1(v172_0),
    .A2(v202_0),
    .Z(v203_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0205_ (
    .A1(v171_0),
    .A2(v203_0),
    .Z(v204_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0206_ (
    .A1(v163_0),
    .A2(v121_0),
    .Z(v205_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0207_ (
    .A1(v163_0),
    .A2(v123_0),
    .ZN(v206_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0208_ (
    .A1(v205_0),
    .A2(v206_0),
    .ZN(v207_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0209_ (
    .A1(v204_0),
    .A2(v207_0),
    .Z(v208_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0210_ (
    .A1(v204_0),
    .A2(v207_0),
    .ZN(v209_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0211_ (
    .A1(v208_0),
    .A2(v209_0),
    .Z(v210_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0212_ (
    .A1(v167_0),
    .A2(v165_0),
    .Z(v211_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0213_ (
    .I(v211_0),
    .ZN(v212_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0214_ (
    .A1(v164_0),
    .A2(v120_0),
    .ZN(v213_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0215_ (
    .A1(v212_0),
    .A2(v213_0),
    .ZN(v214_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0216_ (
    .A1(v210_0),
    .A2(v214_0),
    .Z(v215_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0217_ (
    .A1(v203_0),
    .A2(v171_0),
    .Z(v216_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0218_ (
    .A1(v203_0),
    .A2(v172_0),
    .ZN(v217_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0219_ (
    .A1(v216_0),
    .A2(v217_0),
    .ZN(v218_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0220_ (
    .A1(v197_0),
    .A2(v191_0),
    .Z(v219_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0221_ (
    .A1(v195_0),
    .A2(v194_0),
    .ZN(v220_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0222_ (
    .A1(v219_0),
    .A2(v220_0),
    .ZN(v221_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0223_ (
    .A1(n4),
    .A2(n14),
    .ZN(v222_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0224_ (
    .I(n3),
    .ZN(v223_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0225_ (
    .A1(v223_0),
    .A2(n15),
    .ZN(v224_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0226_ (
    .A1(v222_0),
    .A2(v224_0),
    .Z(v225_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0227_ (
    .A1(n12),
    .A2(n6),
    .ZN(v226_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0228_ (
    .A1(v93_0),
    .A2(v226_0),
    .Z(v227_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0229_ (
    .A1(v180_0),
    .A2(v227_0),
    .ZN(v228_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0230_ (
    .A1(v225_0),
    .A2(v228_0),
    .Z(v229_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0231_ (
    .I(v229_0),
    .ZN(v230_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0232_ (
    .A1(v193_0),
    .A2(v192_0),
    .Z(v231_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0233_ (
    .A1(v230_0),
    .A2(v231_0),
    .Z(v232_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0234_ (
    .A1(v230_0),
    .A2(v231_0),
    .ZN(v233_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0235_ (
    .A1(v232_0),
    .A2(v233_0),
    .ZN(v234_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0236_ (
    .A1(v188_0),
    .A2(v189_0),
    .ZN(v235_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0237_ (
    .A1(v235_0),
    .A2(v187_0),
    .ZN(v236_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0238_ (
    .I(v136_0),
    .ZN(v237_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0239_ (
    .A1(v237_0),
    .A2(v183_0),
    .ZN(v238_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0240_ (
    .A1(v187_0),
    .A2(v238_0),
    .ZN(v239_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0241_ (
    .A1(n11),
    .A2(n7),
    .ZN(v240_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0242_ (
    .A1(v226_0),
    .A2(v240_0),
    .Z(v241_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0243_ (
    .I(v241_0),
    .ZN(v242_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0244_ (
    .A1(n5),
    .A2(n13),
    .ZN(v243_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0245_ (
    .A1(v242_0),
    .A2(v243_0),
    .Z(v244_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0246_ (
    .A1(v242_0),
    .A2(v243_0),
    .ZN(v245_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0247_ (
    .A1(v244_0),
    .A2(v245_0),
    .Z(v246_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0248_ (
    .I(v246_0),
    .ZN(v247_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0249_ (
    .A1(v239_0),
    .A2(v247_0),
    .Z(v248_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0250_ (
    .A1(v236_0),
    .A2(v248_0),
    .Z(v249_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0251_ (
    .A1(v236_0),
    .A2(v248_0),
    .ZN(v250_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0252_ (
    .A1(v249_0),
    .A2(v250_0),
    .ZN(v251_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0253_ (
    .A1(v234_0),
    .A2(v251_0),
    .Z(v252_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0254_ (
    .A1(v190_0),
    .A2(v175_0),
    .ZN(v253_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0255_ (
    .A1(v200_0),
    .A2(v253_0),
    .ZN(v254_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0256_ (
    .A1(v252_0),
    .A2(v254_0),
    .Z(v255_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0257_ (
    .A1(v221_0),
    .A2(v255_0),
    .Z(v256_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0258_ (
    .A1(v218_0),
    .A2(v256_0),
    .Z(v257_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0259_ (
    .A1(v211_0),
    .A2(v210_0),
    .ZN(v258_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0260_ (
    .A1(v209_0),
    .A2(v213_0),
    .ZN(v259_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0261_ (
    .A1(v259_0),
    .A2(v208_0),
    .ZN(v260_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0262_ (
    .A1(v258_0),
    .A2(v260_0),
    .ZN(v261_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0263_ (
    .A1(v257_0),
    .A2(v261_0),
    .Z(v262_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0264_ (
    .A1(v228_0),
    .A2(v225_0),
    .ZN(v263_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0265_ (
    .A1(v232_0),
    .A2(v263_0),
    .ZN(v264_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0266_ (
    .A1(v251_0),
    .A2(v234_0),
    .Z(v265_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0267_ (
    .A1(v265_0),
    .A2(v250_0),
    .ZN(v266_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0268_ (
    .A1(n5),
    .A2(n14),
    .ZN(v267_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0269_ (
    .I(n4),
    .ZN(v268_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0270_ (
    .A1(v268_0),
    .A2(n15),
    .ZN(v269_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0271_ (
    .A1(v267_0),
    .A2(v269_0),
    .Z(v270_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0272_ (
    .A1(v226_0),
    .A2(v241_0),
    .Z(v271_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0273_ (
    .A1(v244_0),
    .A2(v271_0),
    .ZN(v272_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0274_ (
    .A1(v270_0),
    .A2(v272_0),
    .Z(v273_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0275_ (
    .I(v273_0),
    .ZN(v274_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0276_ (
    .A1(v224_0),
    .A2(v222_0),
    .Z(v275_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0277_ (
    .A1(v274_0),
    .A2(v275_0),
    .Z(v276_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0278_ (
    .A1(v274_0),
    .A2(v275_0),
    .ZN(v277_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0279_ (
    .A1(v276_0),
    .A2(v277_0),
    .Z(v278_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0280_ (
    .I(v239_0),
    .ZN(v279_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0281_ (
    .A1(v279_0),
    .A2(v246_0),
    .ZN(v280_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0282_ (
    .A1(v280_0),
    .A2(v187_0),
    .ZN(v281_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0283_ (
    .I(v240_0),
    .ZN(v282_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0284_ (
    .A1(v282_0),
    .A2(n12),
    .ZN(v283_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0285_ (
    .A1(n12),
    .A2(n7),
    .ZN(v284_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0286_ (
    .A1(v240_0),
    .A2(v284_0),
    .ZN(v285_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0287_ (
    .A1(v283_0),
    .A2(v285_0),
    .ZN(v286_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0288_ (
    .A1(n13),
    .A2(n6),
    .ZN(v287_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0289_ (
    .A1(v286_0),
    .A2(v287_0),
    .Z(v288_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0290_ (
    .A1(v286_0),
    .A2(v287_0),
    .ZN(v289_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0291_ (
    .A1(v288_0),
    .A2(v289_0),
    .Z(v290_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0292_ (
    .I(v290_0),
    .ZN(v291_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0293_ (
    .A1(v291_0),
    .A2(v239_0),
    .Z(v292_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0294_ (
    .A1(v281_0),
    .A2(v292_0),
    .Z(v293_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0295_ (
    .A1(v281_0),
    .A2(v292_0),
    .ZN(v294_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0296_ (
    .A1(v293_0),
    .A2(v294_0),
    .Z(v295_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0297_ (
    .A1(v278_0),
    .A2(v295_0),
    .Z(v296_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0298_ (
    .A1(v266_0),
    .A2(v296_0),
    .Z(v297_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0299_ (
    .A1(v264_0),
    .A2(v297_0),
    .Z(v298_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0300_ (
    .A1(v255_0),
    .A2(v221_0),
    .ZN(v299_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0301_ (
    .A1(v254_0),
    .A2(v252_0),
    .ZN(v300_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0302_ (
    .A1(v299_0),
    .A2(v300_0),
    .ZN(v301_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0303_ (
    .A1(v298_0),
    .A2(v301_0),
    .Z(v302_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0304_ (
    .A1(v298_0),
    .A2(v301_0),
    .ZN(v303_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0305_ (
    .A1(v302_0),
    .A2(v303_0),
    .Z(v304_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0306_ (
    .A1(v261_0),
    .A2(v257_0),
    .ZN(v305_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0307_ (
    .A1(v256_0),
    .A2(v218_0),
    .ZN(v306_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0308_ (
    .A1(v305_0),
    .A2(v306_0),
    .ZN(v307_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0309_ (
    .A1(v304_0),
    .A2(v307_0),
    .Z(v308_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0310_ (
    .A1(v297_0),
    .A2(v264_0),
    .ZN(v309_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0311_ (
    .A1(v296_0),
    .A2(v266_0),
    .ZN(v310_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0312_ (
    .A1(v309_0),
    .A2(v310_0),
    .ZN(v311_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0313_ (
    .A1(v272_0),
    .A2(v270_0),
    .ZN(v312_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0314_ (
    .A1(v276_0),
    .A2(v312_0),
    .ZN(v313_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0315_ (
    .A1(v295_0),
    .A2(v278_0),
    .ZN(v314_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0316_ (
    .A1(v314_0),
    .A2(v294_0),
    .ZN(v315_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0317_ (
    .A1(n6),
    .A2(n14),
    .ZN(v316_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0318_ (
    .I(n5),
    .ZN(v317_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0319_ (
    .A1(v317_0),
    .A2(n15),
    .ZN(v318_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0320_ (
    .A1(v316_0),
    .A2(v318_0),
    .Z(v319_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0321_ (
    .A1(v288_0),
    .A2(v283_0),
    .ZN(v320_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0322_ (
    .A1(v319_0),
    .A2(v320_0),
    .Z(v321_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0323_ (
    .I(v321_0),
    .ZN(v322_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0324_ (
    .A1(v269_0),
    .A2(v267_0),
    .Z(v323_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0325_ (
    .A1(v322_0),
    .A2(v323_0),
    .Z(v324_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0326_ (
    .A1(v322_0),
    .A2(v323_0),
    .ZN(v325_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0327_ (
    .A1(v324_0),
    .A2(v325_0),
    .Z(v326_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0328_ (
    .A1(v279_0),
    .A2(v290_0),
    .ZN(v327_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0329_ (
    .A1(v327_0),
    .A2(v187_0),
    .ZN(v328_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0330_ (
    .A1(n13),
    .A2(n7),
    .ZN(v329_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0331_ (
    .A1(v329_0),
    .A2(v286_0),
    .Z(v330_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0332_ (
    .I(v330_0),
    .ZN(v331_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0333_ (
    .A1(v331_0),
    .A2(v239_0),
    .Z(v332_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0334_ (
    .A1(v328_0),
    .A2(v332_0),
    .Z(v333_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0335_ (
    .A1(v328_0),
    .A2(v332_0),
    .ZN(v334_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0336_ (
    .A1(v333_0),
    .A2(v334_0),
    .Z(v335_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0337_ (
    .A1(v326_0),
    .A2(v335_0),
    .Z(v336_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0338_ (
    .A1(v315_0),
    .A2(v336_0),
    .Z(v337_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0339_ (
    .A1(v313_0),
    .A2(v337_0),
    .Z(v338_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0340_ (
    .A1(v311_0),
    .A2(v338_0),
    .Z(v339_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0341_ (
    .A1(v306_0),
    .A2(v303_0),
    .Z(v340_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0342_ (
    .A1(v305_0),
    .A2(v340_0),
    .ZN(v341_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0343_ (
    .A1(v341_0),
    .A2(v302_0),
    .Z(v342_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0344_ (
    .A1(v339_0),
    .A2(v342_0),
    .Z(v343_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0345_ (
    .A1(v320_0),
    .A2(v319_0),
    .ZN(v344_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0346_ (
    .A1(v324_0),
    .A2(v344_0),
    .ZN(v345_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0347_ (
    .A1(v335_0),
    .A2(v326_0),
    .ZN(v346_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0348_ (
    .A1(v346_0),
    .A2(v334_0),
    .ZN(v347_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0349_ (
    .A1(v239_0),
    .A2(v331_0),
    .Z(v348_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0350_ (
    .A1(v348_0),
    .A2(v187_0),
    .ZN(v349_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0351_ (
    .A1(v331_0),
    .A2(v187_0),
    .Z(v350_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0352_ (
    .A1(v349_0),
    .A2(v350_0),
    .ZN(v351_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0353_ (
    .I(v351_0),
    .ZN(v352_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0354_ (
    .A1(v286_0),
    .A2(v329_0),
    .Z(v353_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0355_ (
    .A1(v353_0),
    .A2(v283_0),
    .ZN(v354_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0356_ (
    .I(v354_0),
    .ZN(v355_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0357_ (
    .A1(n14),
    .A2(n7),
    .ZN(v356_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0358_ (
    .I(v356_0),
    .ZN(v357_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0359_ (
    .A1(v73_0),
    .A2(n6),
    .Z(v358_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0360_ (
    .A1(v357_0),
    .A2(v358_0),
    .Z(v359_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0361_ (
    .A1(v355_0),
    .A2(v359_0),
    .Z(v360_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0362_ (
    .A1(v355_0),
    .A2(v359_0),
    .ZN(v361_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0363_ (
    .A1(v360_0),
    .A2(v361_0),
    .Z(v362_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0364_ (
    .I(v362_0),
    .ZN(v363_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0365_ (
    .A1(v318_0),
    .A2(v316_0),
    .Z(v364_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0366_ (
    .A1(v363_0),
    .A2(v364_0),
    .Z(v365_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0367_ (
    .A1(v363_0),
    .A2(v364_0),
    .ZN(v366_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0368_ (
    .A1(v365_0),
    .A2(v366_0),
    .Z(v367_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0369_ (
    .A1(v352_0),
    .A2(v367_0),
    .Z(v368_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0370_ (
    .A1(v347_0),
    .A2(v368_0),
    .Z(v369_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0371_ (
    .A1(v345_0),
    .A2(v369_0),
    .Z(v370_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0372_ (
    .A1(v337_0),
    .A2(v313_0),
    .ZN(v371_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0373_ (
    .A1(v336_0),
    .A2(v315_0),
    .ZN(v372_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0374_ (
    .A1(v371_0),
    .A2(v372_0),
    .ZN(v373_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0375_ (
    .A1(v370_0),
    .A2(v373_0),
    .Z(v374_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0376_ (
    .A1(v370_0),
    .A2(v373_0),
    .ZN(v375_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0377_ (
    .A1(v374_0),
    .A2(v375_0),
    .Z(v376_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0378_ (
    .A1(v342_0),
    .A2(v339_0),
    .ZN(v377_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0379_ (
    .A1(v338_0),
    .A2(v311_0),
    .ZN(v378_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0380_ (
    .A1(v377_0),
    .A2(v378_0),
    .ZN(v379_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0381_ (
    .A1(v376_0),
    .A2(v379_0),
    .Z(v380_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0382_ (
    .A1(v365_0),
    .A2(v360_0),
    .ZN(v381_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0383_ (
    .A1(v358_0),
    .A2(v357_0),
    .ZN(v382_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0384_ (
    .A1(v73_0),
    .A2(n7),
    .Z(v383_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0385_ (
    .A1(v382_0),
    .A2(v383_0),
    .ZN(v384_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0386_ (
    .A1(v384_0),
    .A2(v354_0),
    .Z(v385_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0387_ (
    .A1(v385_0),
    .A2(v352_0),
    .Z(v386_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0388_ (
    .A1(v367_0),
    .A2(v352_0),
    .ZN(v387_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0389_ (
    .A1(v387_0),
    .A2(v350_0),
    .ZN(v388_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0390_ (
    .A1(v386_0),
    .A2(v388_0),
    .Z(v389_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0391_ (
    .A1(v381_0),
    .A2(v389_0),
    .Z(v390_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0392_ (
    .A1(v369_0),
    .A2(v345_0),
    .ZN(v391_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0393_ (
    .A1(v368_0),
    .A2(v347_0),
    .ZN(v392_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0394_ (
    .A1(v391_0),
    .A2(v392_0),
    .ZN(v393_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0395_ (
    .A1(v390_0),
    .A2(v393_0),
    .Z(v394_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0396_ (
    .A1(v379_0),
    .A2(v374_0),
    .ZN(v395_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0397_ (
    .A1(v395_0),
    .A2(v375_0),
    .ZN(v396_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0398_ (
    .A1(v394_0),
    .A2(v396_0),
    .Z(v397_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0399_ (
    .A1(v319_0),
    .A2(v396_0),
    .ZN(v398_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0400_ (
    .A1(v397_0),
    .A2(v398_0),
    .Z(v399_0)
  );

  assign OUT[0] = v331_0;
  assign OUT[1] = v234_0;
  assign OUT[2] = v352_0;
  assign OUT[3] = v151_0;
  assign OUT[4] = v39_0;
  assign OUT[5] = v19_0;
  assign OUT[6] = v66_0;
  assign OUT[7] = v119_0;
  assign OUT[8] = v168_0;
  assign OUT[9] = v215_0;
  assign OUT[10] = v262_0;
  assign OUT[11] = v308_0;
  assign OUT[12] = v343_0;
  assign OUT[13] = v380_0;
  assign OUT[14] = v397_0;
  assign OUT[15] = v399_0;
endmodule
