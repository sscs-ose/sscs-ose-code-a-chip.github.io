# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.820000 BY  2.670000 ;
  PIN BULK
    ANTENNADIFFAREA  0.957000 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.570000 0.470000 2.100000 ;
        RECT 2.350000 0.570000 2.640000 2.100000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  0.462000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 1.460000 2.770000 2.100000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.825000 ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.100000 1.915000 0.270000 ;
        RECT 0.905000 2.400000 1.915000 2.570000 ;
      LAYER mcon ;
        RECT 0.965000 0.100000 1.135000 0.270000 ;
        RECT 0.965000 2.400000 1.135000 2.570000 ;
        RECT 1.325000 0.100000 1.495000 0.270000 ;
        RECT 1.325000 2.400000 1.495000 2.570000 ;
        RECT 1.685000 0.100000 1.855000 0.270000 ;
        RECT 1.685000 2.400000 1.855000 2.570000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.905000 0.000000 1.915000 0.330000 ;
        RECT 0.905000 2.340000 1.915000 2.670000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.570000 2.770000 1.210000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.660000 0.410000 2.010000 ;
      RECT 0.795000 0.490000 0.965000 2.180000 ;
      RECT 1.325000 0.490000 1.495000 2.180000 ;
      RECT 1.855000 0.490000 2.025000 2.180000 ;
      RECT 2.410000 0.660000 2.580000 2.010000 ;
    LAYER mcon ;
      RECT 0.240000 0.710000 0.410000 0.880000 ;
      RECT 0.240000 1.070000 0.410000 1.240000 ;
      RECT 0.240000 1.430000 0.410000 1.600000 ;
      RECT 0.240000 1.790000 0.410000 1.960000 ;
      RECT 0.795000 0.710000 0.965000 0.880000 ;
      RECT 0.795000 1.070000 0.965000 1.240000 ;
      RECT 0.795000 1.430000 0.965000 1.600000 ;
      RECT 0.795000 1.790000 0.965000 1.960000 ;
      RECT 1.325000 0.710000 1.495000 0.880000 ;
      RECT 1.325000 1.070000 1.495000 1.240000 ;
      RECT 1.325000 1.430000 1.495000 1.600000 ;
      RECT 1.325000 1.790000 1.495000 1.960000 ;
      RECT 1.855000 0.710000 2.025000 0.880000 ;
      RECT 1.855000 1.070000 2.025000 1.240000 ;
      RECT 1.855000 1.430000 2.025000 1.600000 ;
      RECT 1.855000 1.790000 2.025000 1.960000 ;
      RECT 2.410000 0.710000 2.580000 0.880000 ;
      RECT 2.410000 1.070000 2.580000 1.240000 ;
      RECT 2.410000 1.430000 2.580000 1.600000 ;
      RECT 2.410000 1.790000 2.580000 1.960000 ;
    LAYER met1 ;
      RECT 0.750000 0.570000 1.010000 2.100000 ;
      RECT 1.280000 0.570000 1.540000 2.100000 ;
      RECT 1.810000 0.570000 2.070000 2.100000 ;
    LAYER via ;
      RECT 0.750000 0.600000 1.010000 0.860000 ;
      RECT 0.750000 0.920000 1.010000 1.180000 ;
      RECT 1.280000 1.490000 1.540000 1.750000 ;
      RECT 1.280000 1.810000 1.540000 2.070000 ;
      RECT 1.810000 0.600000 2.070000 0.860000 ;
      RECT 1.810000 0.920000 2.070000 1.180000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25
END LIBRARY
