** sch_path: /foss/designs/can_ic_v3/jupyter/xschem/can_ic/can_ic.sch
**.subckt can_ic DRIVER_VCC TX CAN+ CAN- DRIVER_VSS RX RS
*.iopin DRIVER_VCC
*.iopin DRIVER_VSS
*.ipin TX
*.opin CAN+
*.opin CAN-
*.iopin RS
*.opin RX
XM4 CAN- inv_tx DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=0.15 W=12 nf=1 ad=3.48 as=3.48 pd=24.58 ps=24.58
+ nrd=0.0241666666666667 nrs=0.0241666666666667 sa=0 sb=0 sd=0 mult=20 m=20
XM5 CAN+ TX DRIVER_VCC DRIVER_VCC sky130_fd_pr__pfet_01v8 L=0.15 W=30 nf=1 ad=8.7 as=8.7 pd=60.58 ps=60.58 nrd=0.00966666666666667
+ nrs=0.00966666666666667 sa=0 sb=0 sd=0 mult=20 m=20
XM1 inv_tx TX DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=0.8 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0
+ sb=0 sd=0 mult=4 m=4
XM2 net1 net2 DRIVER_VCC DRIVER_VCC sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 net2 net2 DRIVER_VCC DRIVER_VCC sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM6 net1 net1 DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM7 net8 net1 RS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM8 net3 net2 DRIVER_VCC DRIVER_VCC sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM9 net4 net6 net3 DRIVER_VCC sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM10 net5 net7 net3 DRIVER_VCC sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM11 net4 net4 DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM12 net5 net4 DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM13 RX net5 DRIVER_VSS DRIVER_VSS sky130_fd_pr__nfet_01v8 L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XR7 inv_tx DRIVER_VCC DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=40 mult=1 m=1
XR5 net7 CAN- DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=42 mult=1 m=1
XR1 CAN+ net6 DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=42 mult=1 m=1
XR3 DRIVER_VCC RX DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=42 mult=1 m=1
XR4 RX net7 DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=64 mult=1 m=1
XR2 DRIVER_VCC TX DRIVER_VCC sky130_fd_pr__res_high_po_1p41 L=42 mult=1 m=1
**.ends
.end
