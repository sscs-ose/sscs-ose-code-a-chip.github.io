# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  3.870000 BY  3.540000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.895000 3.940000 2.535000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.215000 0.000000 2.795000 0.695000 ;
        RECT 1.215000 2.845000 2.795000 3.540000 ;
      LAYER mcon ;
        RECT 1.275000 0.095000 1.445000 0.265000 ;
        RECT 1.275000 0.455000 1.445000 0.625000 ;
        RECT 1.275000 2.915000 1.445000 3.085000 ;
        RECT 1.275000 3.275000 1.445000 3.445000 ;
        RECT 1.685000 0.095000 1.855000 0.265000 ;
        RECT 1.685000 0.455000 1.855000 0.625000 ;
        RECT 1.685000 2.915000 1.855000 3.085000 ;
        RECT 1.685000 3.275000 1.855000 3.445000 ;
        RECT 2.155000 0.095000 2.325000 0.265000 ;
        RECT 2.155000 0.455000 2.325000 0.625000 ;
        RECT 2.155000 2.915000 2.325000 3.085000 ;
        RECT 2.155000 3.275000 2.325000 3.445000 ;
        RECT 2.565000 0.095000 2.735000 0.265000 ;
        RECT 2.565000 0.455000 2.735000 0.625000 ;
        RECT 2.565000 2.915000 2.735000 3.085000 ;
        RECT 2.565000 3.275000 2.735000 3.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.215000 0.000000 2.795000 0.685000 ;
        RECT 1.215000 2.855000 2.795000 3.540000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.005000 3.940000 1.645000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.072500 ;
    ANTENNAGATEAREA  0.247500 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.005000 0.500000 2.535000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.510000 1.005000 3.805000 2.535000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 0.800000 2.615000 ;
      RECT 0.600000 0.485000 0.930000 0.815000 ;
      RECT 0.600000 0.815000 0.800000 0.925000 ;
      RECT 0.600000 2.615000 0.800000 2.725000 ;
      RECT 0.600000 2.725000 0.930000 3.055000 ;
      RECT 1.060000 0.925000 1.230000 2.615000 ;
      RECT 1.490000 0.925000 1.660000 2.615000 ;
      RECT 1.920000 0.925000 2.090000 2.615000 ;
      RECT 2.350000 0.925000 2.520000 2.615000 ;
      RECT 2.780000 0.925000 2.950000 2.615000 ;
      RECT 3.080000 0.485000 3.410000 0.815000 ;
      RECT 3.080000 2.725000 3.410000 3.055000 ;
      RECT 3.210000 0.815000 3.410000 0.925000 ;
      RECT 3.210000 0.925000 3.805000 2.615000 ;
      RECT 3.210000 2.615000 3.410000 2.725000 ;
    LAYER mcon ;
      RECT 0.300000 1.145000 0.470000 1.315000 ;
      RECT 0.300000 1.505000 0.470000 1.675000 ;
      RECT 0.300000 1.865000 0.470000 2.035000 ;
      RECT 0.300000 2.225000 0.470000 2.395000 ;
      RECT 1.060000 1.145000 1.230000 1.315000 ;
      RECT 1.060000 1.505000 1.230000 1.675000 ;
      RECT 1.060000 1.865000 1.230000 2.035000 ;
      RECT 1.060000 2.225000 1.230000 2.395000 ;
      RECT 1.490000 1.145000 1.660000 1.315000 ;
      RECT 1.490000 1.505000 1.660000 1.675000 ;
      RECT 1.490000 1.865000 1.660000 2.035000 ;
      RECT 1.490000 2.225000 1.660000 2.395000 ;
      RECT 1.920000 1.145000 2.090000 1.315000 ;
      RECT 1.920000 1.505000 2.090000 1.675000 ;
      RECT 1.920000 1.865000 2.090000 2.035000 ;
      RECT 1.920000 2.225000 2.090000 2.395000 ;
      RECT 2.350000 1.145000 2.520000 1.315000 ;
      RECT 2.350000 1.505000 2.520000 1.675000 ;
      RECT 2.350000 1.865000 2.520000 2.035000 ;
      RECT 2.350000 2.225000 2.520000 2.395000 ;
      RECT 2.780000 1.145000 2.950000 1.315000 ;
      RECT 2.780000 1.505000 2.950000 1.675000 ;
      RECT 2.780000 1.865000 2.950000 2.035000 ;
      RECT 2.780000 2.225000 2.950000 2.395000 ;
      RECT 3.540000 1.145000 3.710000 1.315000 ;
      RECT 3.540000 1.505000 3.710000 1.675000 ;
      RECT 3.540000 1.865000 3.710000 2.035000 ;
      RECT 3.540000 2.225000 3.710000 2.395000 ;
    LAYER met1 ;
      RECT 1.015000 1.005000 1.275000 2.535000 ;
      RECT 1.445000 1.005000 1.705000 2.535000 ;
      RECT 1.875000 1.005000 2.135000 2.535000 ;
      RECT 2.305000 1.005000 2.565000 2.535000 ;
      RECT 2.735000 1.005000 2.995000 2.535000 ;
    LAYER via ;
      RECT 1.015000 1.035000 1.275000 1.295000 ;
      RECT 1.015000 1.355000 1.275000 1.615000 ;
      RECT 1.445000 1.925000 1.705000 2.185000 ;
      RECT 1.445000 2.245000 1.705000 2.505000 ;
      RECT 1.875000 1.035000 2.135000 1.295000 ;
      RECT 1.875000 1.355000 2.135000 1.615000 ;
      RECT 2.305000 1.925000 2.565000 2.185000 ;
      RECT 2.305000 2.245000 2.565000 2.505000 ;
      RECT 2.735000 1.035000 2.995000 1.295000 ;
      RECT 2.735000 1.355000 2.995000 1.615000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15
END LIBRARY
