MACRO NMOS_S_12565100_X74_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_12565100_X74_Y2 0 0 ;
  SIZE 65360 BY 13440 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 32110 260 32390 6460 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 32540 4460 32820 10660 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 32970 680 33250 12760 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 13105 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 13105 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 13105 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 13105 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 13105 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 13105 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 13105 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 13105 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 13105 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 13105 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 9745 ;
    LAYER M1 ;
      RECT 9765 9995 10015 11005 ;
    LAYER M1 ;
      RECT 9765 12095 10015 13105 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 6215 10445 9745 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 9745 ;
    LAYER M1 ;
      RECT 10625 9995 10875 11005 ;
    LAYER M1 ;
      RECT 10625 12095 10875 13105 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11055 6215 11305 9745 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 9745 ;
    LAYER M1 ;
      RECT 11485 9995 11735 11005 ;
    LAYER M1 ;
      RECT 11485 12095 11735 13105 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 11915 6215 12165 9745 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 9745 ;
    LAYER M1 ;
      RECT 12345 9995 12595 11005 ;
    LAYER M1 ;
      RECT 12345 12095 12595 13105 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 12775 6215 13025 9745 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 9745 ;
    LAYER M1 ;
      RECT 13205 9995 13455 11005 ;
    LAYER M1 ;
      RECT 13205 12095 13455 13105 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 13635 6215 13885 9745 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 9745 ;
    LAYER M1 ;
      RECT 14065 9995 14315 11005 ;
    LAYER M1 ;
      RECT 14065 12095 14315 13105 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14495 6215 14745 9745 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 9745 ;
    LAYER M1 ;
      RECT 14925 9995 15175 11005 ;
    LAYER M1 ;
      RECT 14925 12095 15175 13105 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15355 6215 15605 9745 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 9745 ;
    LAYER M1 ;
      RECT 15785 9995 16035 11005 ;
    LAYER M1 ;
      RECT 15785 12095 16035 13105 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16215 6215 16465 9745 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 9745 ;
    LAYER M1 ;
      RECT 16645 9995 16895 11005 ;
    LAYER M1 ;
      RECT 16645 12095 16895 13105 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17075 6215 17325 9745 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 9745 ;
    LAYER M1 ;
      RECT 17505 9995 17755 11005 ;
    LAYER M1 ;
      RECT 17505 12095 17755 13105 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 17935 6215 18185 9745 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 9745 ;
    LAYER M1 ;
      RECT 18365 9995 18615 11005 ;
    LAYER M1 ;
      RECT 18365 12095 18615 13105 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 18795 6215 19045 9745 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 9745 ;
    LAYER M1 ;
      RECT 19225 9995 19475 11005 ;
    LAYER M1 ;
      RECT 19225 12095 19475 13105 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 19655 6215 19905 9745 ;
    LAYER M1 ;
      RECT 20085 335 20335 3865 ;
    LAYER M1 ;
      RECT 20085 4115 20335 5125 ;
    LAYER M1 ;
      RECT 20085 6215 20335 9745 ;
    LAYER M1 ;
      RECT 20085 9995 20335 11005 ;
    LAYER M1 ;
      RECT 20085 12095 20335 13105 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20515 6215 20765 9745 ;
    LAYER M1 ;
      RECT 20945 335 21195 3865 ;
    LAYER M1 ;
      RECT 20945 4115 21195 5125 ;
    LAYER M1 ;
      RECT 20945 6215 21195 9745 ;
    LAYER M1 ;
      RECT 20945 9995 21195 11005 ;
    LAYER M1 ;
      RECT 20945 12095 21195 13105 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 21375 6215 21625 9745 ;
    LAYER M1 ;
      RECT 21805 335 22055 3865 ;
    LAYER M1 ;
      RECT 21805 4115 22055 5125 ;
    LAYER M1 ;
      RECT 21805 6215 22055 9745 ;
    LAYER M1 ;
      RECT 21805 9995 22055 11005 ;
    LAYER M1 ;
      RECT 21805 12095 22055 13105 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22235 6215 22485 9745 ;
    LAYER M1 ;
      RECT 22665 335 22915 3865 ;
    LAYER M1 ;
      RECT 22665 4115 22915 5125 ;
    LAYER M1 ;
      RECT 22665 6215 22915 9745 ;
    LAYER M1 ;
      RECT 22665 9995 22915 11005 ;
    LAYER M1 ;
      RECT 22665 12095 22915 13105 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23095 6215 23345 9745 ;
    LAYER M1 ;
      RECT 23525 335 23775 3865 ;
    LAYER M1 ;
      RECT 23525 4115 23775 5125 ;
    LAYER M1 ;
      RECT 23525 6215 23775 9745 ;
    LAYER M1 ;
      RECT 23525 9995 23775 11005 ;
    LAYER M1 ;
      RECT 23525 12095 23775 13105 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 23955 6215 24205 9745 ;
    LAYER M1 ;
      RECT 24385 335 24635 3865 ;
    LAYER M1 ;
      RECT 24385 4115 24635 5125 ;
    LAYER M1 ;
      RECT 24385 6215 24635 9745 ;
    LAYER M1 ;
      RECT 24385 9995 24635 11005 ;
    LAYER M1 ;
      RECT 24385 12095 24635 13105 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M1 ;
      RECT 24815 6215 25065 9745 ;
    LAYER M1 ;
      RECT 25245 335 25495 3865 ;
    LAYER M1 ;
      RECT 25245 4115 25495 5125 ;
    LAYER M1 ;
      RECT 25245 6215 25495 9745 ;
    LAYER M1 ;
      RECT 25245 9995 25495 11005 ;
    LAYER M1 ;
      RECT 25245 12095 25495 13105 ;
    LAYER M1 ;
      RECT 25675 335 25925 3865 ;
    LAYER M1 ;
      RECT 25675 6215 25925 9745 ;
    LAYER M1 ;
      RECT 26105 335 26355 3865 ;
    LAYER M1 ;
      RECT 26105 4115 26355 5125 ;
    LAYER M1 ;
      RECT 26105 6215 26355 9745 ;
    LAYER M1 ;
      RECT 26105 9995 26355 11005 ;
    LAYER M1 ;
      RECT 26105 12095 26355 13105 ;
    LAYER M1 ;
      RECT 26535 335 26785 3865 ;
    LAYER M1 ;
      RECT 26535 6215 26785 9745 ;
    LAYER M1 ;
      RECT 26965 335 27215 3865 ;
    LAYER M1 ;
      RECT 26965 4115 27215 5125 ;
    LAYER M1 ;
      RECT 26965 6215 27215 9745 ;
    LAYER M1 ;
      RECT 26965 9995 27215 11005 ;
    LAYER M1 ;
      RECT 26965 12095 27215 13105 ;
    LAYER M1 ;
      RECT 27395 335 27645 3865 ;
    LAYER M1 ;
      RECT 27395 6215 27645 9745 ;
    LAYER M1 ;
      RECT 27825 335 28075 3865 ;
    LAYER M1 ;
      RECT 27825 4115 28075 5125 ;
    LAYER M1 ;
      RECT 27825 6215 28075 9745 ;
    LAYER M1 ;
      RECT 27825 9995 28075 11005 ;
    LAYER M1 ;
      RECT 27825 12095 28075 13105 ;
    LAYER M1 ;
      RECT 28255 335 28505 3865 ;
    LAYER M1 ;
      RECT 28255 6215 28505 9745 ;
    LAYER M1 ;
      RECT 28685 335 28935 3865 ;
    LAYER M1 ;
      RECT 28685 4115 28935 5125 ;
    LAYER M1 ;
      RECT 28685 6215 28935 9745 ;
    LAYER M1 ;
      RECT 28685 9995 28935 11005 ;
    LAYER M1 ;
      RECT 28685 12095 28935 13105 ;
    LAYER M1 ;
      RECT 29115 335 29365 3865 ;
    LAYER M1 ;
      RECT 29115 6215 29365 9745 ;
    LAYER M1 ;
      RECT 29545 335 29795 3865 ;
    LAYER M1 ;
      RECT 29545 4115 29795 5125 ;
    LAYER M1 ;
      RECT 29545 6215 29795 9745 ;
    LAYER M1 ;
      RECT 29545 9995 29795 11005 ;
    LAYER M1 ;
      RECT 29545 12095 29795 13105 ;
    LAYER M1 ;
      RECT 29975 335 30225 3865 ;
    LAYER M1 ;
      RECT 29975 6215 30225 9745 ;
    LAYER M1 ;
      RECT 30405 335 30655 3865 ;
    LAYER M1 ;
      RECT 30405 4115 30655 5125 ;
    LAYER M1 ;
      RECT 30405 6215 30655 9745 ;
    LAYER M1 ;
      RECT 30405 9995 30655 11005 ;
    LAYER M1 ;
      RECT 30405 12095 30655 13105 ;
    LAYER M1 ;
      RECT 30835 335 31085 3865 ;
    LAYER M1 ;
      RECT 30835 6215 31085 9745 ;
    LAYER M1 ;
      RECT 31265 335 31515 3865 ;
    LAYER M1 ;
      RECT 31265 4115 31515 5125 ;
    LAYER M1 ;
      RECT 31265 6215 31515 9745 ;
    LAYER M1 ;
      RECT 31265 9995 31515 11005 ;
    LAYER M1 ;
      RECT 31265 12095 31515 13105 ;
    LAYER M1 ;
      RECT 31695 335 31945 3865 ;
    LAYER M1 ;
      RECT 31695 6215 31945 9745 ;
    LAYER M1 ;
      RECT 32125 335 32375 3865 ;
    LAYER M1 ;
      RECT 32125 4115 32375 5125 ;
    LAYER M1 ;
      RECT 32125 6215 32375 9745 ;
    LAYER M1 ;
      RECT 32125 9995 32375 11005 ;
    LAYER M1 ;
      RECT 32125 12095 32375 13105 ;
    LAYER M1 ;
      RECT 32555 335 32805 3865 ;
    LAYER M1 ;
      RECT 32555 6215 32805 9745 ;
    LAYER M1 ;
      RECT 32985 335 33235 3865 ;
    LAYER M1 ;
      RECT 32985 4115 33235 5125 ;
    LAYER M1 ;
      RECT 32985 6215 33235 9745 ;
    LAYER M1 ;
      RECT 32985 9995 33235 11005 ;
    LAYER M1 ;
      RECT 32985 12095 33235 13105 ;
    LAYER M1 ;
      RECT 33415 335 33665 3865 ;
    LAYER M1 ;
      RECT 33415 6215 33665 9745 ;
    LAYER M1 ;
      RECT 33845 335 34095 3865 ;
    LAYER M1 ;
      RECT 33845 4115 34095 5125 ;
    LAYER M1 ;
      RECT 33845 6215 34095 9745 ;
    LAYER M1 ;
      RECT 33845 9995 34095 11005 ;
    LAYER M1 ;
      RECT 33845 12095 34095 13105 ;
    LAYER M1 ;
      RECT 34275 335 34525 3865 ;
    LAYER M1 ;
      RECT 34275 6215 34525 9745 ;
    LAYER M1 ;
      RECT 34705 335 34955 3865 ;
    LAYER M1 ;
      RECT 34705 4115 34955 5125 ;
    LAYER M1 ;
      RECT 34705 6215 34955 9745 ;
    LAYER M1 ;
      RECT 34705 9995 34955 11005 ;
    LAYER M1 ;
      RECT 34705 12095 34955 13105 ;
    LAYER M1 ;
      RECT 35135 335 35385 3865 ;
    LAYER M1 ;
      RECT 35135 6215 35385 9745 ;
    LAYER M1 ;
      RECT 35565 335 35815 3865 ;
    LAYER M1 ;
      RECT 35565 4115 35815 5125 ;
    LAYER M1 ;
      RECT 35565 6215 35815 9745 ;
    LAYER M1 ;
      RECT 35565 9995 35815 11005 ;
    LAYER M1 ;
      RECT 35565 12095 35815 13105 ;
    LAYER M1 ;
      RECT 35995 335 36245 3865 ;
    LAYER M1 ;
      RECT 35995 6215 36245 9745 ;
    LAYER M1 ;
      RECT 36425 335 36675 3865 ;
    LAYER M1 ;
      RECT 36425 4115 36675 5125 ;
    LAYER M1 ;
      RECT 36425 6215 36675 9745 ;
    LAYER M1 ;
      RECT 36425 9995 36675 11005 ;
    LAYER M1 ;
      RECT 36425 12095 36675 13105 ;
    LAYER M1 ;
      RECT 36855 335 37105 3865 ;
    LAYER M1 ;
      RECT 36855 6215 37105 9745 ;
    LAYER M1 ;
      RECT 37285 335 37535 3865 ;
    LAYER M1 ;
      RECT 37285 4115 37535 5125 ;
    LAYER M1 ;
      RECT 37285 6215 37535 9745 ;
    LAYER M1 ;
      RECT 37285 9995 37535 11005 ;
    LAYER M1 ;
      RECT 37285 12095 37535 13105 ;
    LAYER M1 ;
      RECT 37715 335 37965 3865 ;
    LAYER M1 ;
      RECT 37715 6215 37965 9745 ;
    LAYER M1 ;
      RECT 38145 335 38395 3865 ;
    LAYER M1 ;
      RECT 38145 4115 38395 5125 ;
    LAYER M1 ;
      RECT 38145 6215 38395 9745 ;
    LAYER M1 ;
      RECT 38145 9995 38395 11005 ;
    LAYER M1 ;
      RECT 38145 12095 38395 13105 ;
    LAYER M1 ;
      RECT 38575 335 38825 3865 ;
    LAYER M1 ;
      RECT 38575 6215 38825 9745 ;
    LAYER M1 ;
      RECT 39005 335 39255 3865 ;
    LAYER M1 ;
      RECT 39005 4115 39255 5125 ;
    LAYER M1 ;
      RECT 39005 6215 39255 9745 ;
    LAYER M1 ;
      RECT 39005 9995 39255 11005 ;
    LAYER M1 ;
      RECT 39005 12095 39255 13105 ;
    LAYER M1 ;
      RECT 39435 335 39685 3865 ;
    LAYER M1 ;
      RECT 39435 6215 39685 9745 ;
    LAYER M1 ;
      RECT 39865 335 40115 3865 ;
    LAYER M1 ;
      RECT 39865 4115 40115 5125 ;
    LAYER M1 ;
      RECT 39865 6215 40115 9745 ;
    LAYER M1 ;
      RECT 39865 9995 40115 11005 ;
    LAYER M1 ;
      RECT 39865 12095 40115 13105 ;
    LAYER M1 ;
      RECT 40295 335 40545 3865 ;
    LAYER M1 ;
      RECT 40295 6215 40545 9745 ;
    LAYER M1 ;
      RECT 40725 335 40975 3865 ;
    LAYER M1 ;
      RECT 40725 4115 40975 5125 ;
    LAYER M1 ;
      RECT 40725 6215 40975 9745 ;
    LAYER M1 ;
      RECT 40725 9995 40975 11005 ;
    LAYER M1 ;
      RECT 40725 12095 40975 13105 ;
    LAYER M1 ;
      RECT 41155 335 41405 3865 ;
    LAYER M1 ;
      RECT 41155 6215 41405 9745 ;
    LAYER M1 ;
      RECT 41585 335 41835 3865 ;
    LAYER M1 ;
      RECT 41585 4115 41835 5125 ;
    LAYER M1 ;
      RECT 41585 6215 41835 9745 ;
    LAYER M1 ;
      RECT 41585 9995 41835 11005 ;
    LAYER M1 ;
      RECT 41585 12095 41835 13105 ;
    LAYER M1 ;
      RECT 42015 335 42265 3865 ;
    LAYER M1 ;
      RECT 42015 6215 42265 9745 ;
    LAYER M1 ;
      RECT 42445 335 42695 3865 ;
    LAYER M1 ;
      RECT 42445 4115 42695 5125 ;
    LAYER M1 ;
      RECT 42445 6215 42695 9745 ;
    LAYER M1 ;
      RECT 42445 9995 42695 11005 ;
    LAYER M1 ;
      RECT 42445 12095 42695 13105 ;
    LAYER M1 ;
      RECT 42875 335 43125 3865 ;
    LAYER M1 ;
      RECT 42875 6215 43125 9745 ;
    LAYER M1 ;
      RECT 43305 335 43555 3865 ;
    LAYER M1 ;
      RECT 43305 4115 43555 5125 ;
    LAYER M1 ;
      RECT 43305 6215 43555 9745 ;
    LAYER M1 ;
      RECT 43305 9995 43555 11005 ;
    LAYER M1 ;
      RECT 43305 12095 43555 13105 ;
    LAYER M1 ;
      RECT 43735 335 43985 3865 ;
    LAYER M1 ;
      RECT 43735 6215 43985 9745 ;
    LAYER M1 ;
      RECT 44165 335 44415 3865 ;
    LAYER M1 ;
      RECT 44165 4115 44415 5125 ;
    LAYER M1 ;
      RECT 44165 6215 44415 9745 ;
    LAYER M1 ;
      RECT 44165 9995 44415 11005 ;
    LAYER M1 ;
      RECT 44165 12095 44415 13105 ;
    LAYER M1 ;
      RECT 44595 335 44845 3865 ;
    LAYER M1 ;
      RECT 44595 6215 44845 9745 ;
    LAYER M1 ;
      RECT 45025 335 45275 3865 ;
    LAYER M1 ;
      RECT 45025 4115 45275 5125 ;
    LAYER M1 ;
      RECT 45025 6215 45275 9745 ;
    LAYER M1 ;
      RECT 45025 9995 45275 11005 ;
    LAYER M1 ;
      RECT 45025 12095 45275 13105 ;
    LAYER M1 ;
      RECT 45455 335 45705 3865 ;
    LAYER M1 ;
      RECT 45455 6215 45705 9745 ;
    LAYER M1 ;
      RECT 45885 335 46135 3865 ;
    LAYER M1 ;
      RECT 45885 4115 46135 5125 ;
    LAYER M1 ;
      RECT 45885 6215 46135 9745 ;
    LAYER M1 ;
      RECT 45885 9995 46135 11005 ;
    LAYER M1 ;
      RECT 45885 12095 46135 13105 ;
    LAYER M1 ;
      RECT 46315 335 46565 3865 ;
    LAYER M1 ;
      RECT 46315 6215 46565 9745 ;
    LAYER M1 ;
      RECT 46745 335 46995 3865 ;
    LAYER M1 ;
      RECT 46745 4115 46995 5125 ;
    LAYER M1 ;
      RECT 46745 6215 46995 9745 ;
    LAYER M1 ;
      RECT 46745 9995 46995 11005 ;
    LAYER M1 ;
      RECT 46745 12095 46995 13105 ;
    LAYER M1 ;
      RECT 47175 335 47425 3865 ;
    LAYER M1 ;
      RECT 47175 6215 47425 9745 ;
    LAYER M1 ;
      RECT 47605 335 47855 3865 ;
    LAYER M1 ;
      RECT 47605 4115 47855 5125 ;
    LAYER M1 ;
      RECT 47605 6215 47855 9745 ;
    LAYER M1 ;
      RECT 47605 9995 47855 11005 ;
    LAYER M1 ;
      RECT 47605 12095 47855 13105 ;
    LAYER M1 ;
      RECT 48035 335 48285 3865 ;
    LAYER M1 ;
      RECT 48035 6215 48285 9745 ;
    LAYER M1 ;
      RECT 48465 335 48715 3865 ;
    LAYER M1 ;
      RECT 48465 4115 48715 5125 ;
    LAYER M1 ;
      RECT 48465 6215 48715 9745 ;
    LAYER M1 ;
      RECT 48465 9995 48715 11005 ;
    LAYER M1 ;
      RECT 48465 12095 48715 13105 ;
    LAYER M1 ;
      RECT 48895 335 49145 3865 ;
    LAYER M1 ;
      RECT 48895 6215 49145 9745 ;
    LAYER M1 ;
      RECT 49325 335 49575 3865 ;
    LAYER M1 ;
      RECT 49325 4115 49575 5125 ;
    LAYER M1 ;
      RECT 49325 6215 49575 9745 ;
    LAYER M1 ;
      RECT 49325 9995 49575 11005 ;
    LAYER M1 ;
      RECT 49325 12095 49575 13105 ;
    LAYER M1 ;
      RECT 49755 335 50005 3865 ;
    LAYER M1 ;
      RECT 49755 6215 50005 9745 ;
    LAYER M1 ;
      RECT 50185 335 50435 3865 ;
    LAYER M1 ;
      RECT 50185 4115 50435 5125 ;
    LAYER M1 ;
      RECT 50185 6215 50435 9745 ;
    LAYER M1 ;
      RECT 50185 9995 50435 11005 ;
    LAYER M1 ;
      RECT 50185 12095 50435 13105 ;
    LAYER M1 ;
      RECT 50615 335 50865 3865 ;
    LAYER M1 ;
      RECT 50615 6215 50865 9745 ;
    LAYER M1 ;
      RECT 51045 335 51295 3865 ;
    LAYER M1 ;
      RECT 51045 4115 51295 5125 ;
    LAYER M1 ;
      RECT 51045 6215 51295 9745 ;
    LAYER M1 ;
      RECT 51045 9995 51295 11005 ;
    LAYER M1 ;
      RECT 51045 12095 51295 13105 ;
    LAYER M1 ;
      RECT 51475 335 51725 3865 ;
    LAYER M1 ;
      RECT 51475 6215 51725 9745 ;
    LAYER M1 ;
      RECT 51905 335 52155 3865 ;
    LAYER M1 ;
      RECT 51905 4115 52155 5125 ;
    LAYER M1 ;
      RECT 51905 6215 52155 9745 ;
    LAYER M1 ;
      RECT 51905 9995 52155 11005 ;
    LAYER M1 ;
      RECT 51905 12095 52155 13105 ;
    LAYER M1 ;
      RECT 52335 335 52585 3865 ;
    LAYER M1 ;
      RECT 52335 6215 52585 9745 ;
    LAYER M1 ;
      RECT 52765 335 53015 3865 ;
    LAYER M1 ;
      RECT 52765 4115 53015 5125 ;
    LAYER M1 ;
      RECT 52765 6215 53015 9745 ;
    LAYER M1 ;
      RECT 52765 9995 53015 11005 ;
    LAYER M1 ;
      RECT 52765 12095 53015 13105 ;
    LAYER M1 ;
      RECT 53195 335 53445 3865 ;
    LAYER M1 ;
      RECT 53195 6215 53445 9745 ;
    LAYER M1 ;
      RECT 53625 335 53875 3865 ;
    LAYER M1 ;
      RECT 53625 4115 53875 5125 ;
    LAYER M1 ;
      RECT 53625 6215 53875 9745 ;
    LAYER M1 ;
      RECT 53625 9995 53875 11005 ;
    LAYER M1 ;
      RECT 53625 12095 53875 13105 ;
    LAYER M1 ;
      RECT 54055 335 54305 3865 ;
    LAYER M1 ;
      RECT 54055 6215 54305 9745 ;
    LAYER M1 ;
      RECT 54485 335 54735 3865 ;
    LAYER M1 ;
      RECT 54485 4115 54735 5125 ;
    LAYER M1 ;
      RECT 54485 6215 54735 9745 ;
    LAYER M1 ;
      RECT 54485 9995 54735 11005 ;
    LAYER M1 ;
      RECT 54485 12095 54735 13105 ;
    LAYER M1 ;
      RECT 54915 335 55165 3865 ;
    LAYER M1 ;
      RECT 54915 6215 55165 9745 ;
    LAYER M1 ;
      RECT 55345 335 55595 3865 ;
    LAYER M1 ;
      RECT 55345 4115 55595 5125 ;
    LAYER M1 ;
      RECT 55345 6215 55595 9745 ;
    LAYER M1 ;
      RECT 55345 9995 55595 11005 ;
    LAYER M1 ;
      RECT 55345 12095 55595 13105 ;
    LAYER M1 ;
      RECT 55775 335 56025 3865 ;
    LAYER M1 ;
      RECT 55775 6215 56025 9745 ;
    LAYER M1 ;
      RECT 56205 335 56455 3865 ;
    LAYER M1 ;
      RECT 56205 4115 56455 5125 ;
    LAYER M1 ;
      RECT 56205 6215 56455 9745 ;
    LAYER M1 ;
      RECT 56205 9995 56455 11005 ;
    LAYER M1 ;
      RECT 56205 12095 56455 13105 ;
    LAYER M1 ;
      RECT 56635 335 56885 3865 ;
    LAYER M1 ;
      RECT 56635 6215 56885 9745 ;
    LAYER M1 ;
      RECT 57065 335 57315 3865 ;
    LAYER M1 ;
      RECT 57065 4115 57315 5125 ;
    LAYER M1 ;
      RECT 57065 6215 57315 9745 ;
    LAYER M1 ;
      RECT 57065 9995 57315 11005 ;
    LAYER M1 ;
      RECT 57065 12095 57315 13105 ;
    LAYER M1 ;
      RECT 57495 335 57745 3865 ;
    LAYER M1 ;
      RECT 57495 6215 57745 9745 ;
    LAYER M1 ;
      RECT 57925 335 58175 3865 ;
    LAYER M1 ;
      RECT 57925 4115 58175 5125 ;
    LAYER M1 ;
      RECT 57925 6215 58175 9745 ;
    LAYER M1 ;
      RECT 57925 9995 58175 11005 ;
    LAYER M1 ;
      RECT 57925 12095 58175 13105 ;
    LAYER M1 ;
      RECT 58355 335 58605 3865 ;
    LAYER M1 ;
      RECT 58355 6215 58605 9745 ;
    LAYER M1 ;
      RECT 58785 335 59035 3865 ;
    LAYER M1 ;
      RECT 58785 4115 59035 5125 ;
    LAYER M1 ;
      RECT 58785 6215 59035 9745 ;
    LAYER M1 ;
      RECT 58785 9995 59035 11005 ;
    LAYER M1 ;
      RECT 58785 12095 59035 13105 ;
    LAYER M1 ;
      RECT 59215 335 59465 3865 ;
    LAYER M1 ;
      RECT 59215 6215 59465 9745 ;
    LAYER M1 ;
      RECT 59645 335 59895 3865 ;
    LAYER M1 ;
      RECT 59645 4115 59895 5125 ;
    LAYER M1 ;
      RECT 59645 6215 59895 9745 ;
    LAYER M1 ;
      RECT 59645 9995 59895 11005 ;
    LAYER M1 ;
      RECT 59645 12095 59895 13105 ;
    LAYER M1 ;
      RECT 60075 335 60325 3865 ;
    LAYER M1 ;
      RECT 60075 6215 60325 9745 ;
    LAYER M1 ;
      RECT 60505 335 60755 3865 ;
    LAYER M1 ;
      RECT 60505 4115 60755 5125 ;
    LAYER M1 ;
      RECT 60505 6215 60755 9745 ;
    LAYER M1 ;
      RECT 60505 9995 60755 11005 ;
    LAYER M1 ;
      RECT 60505 12095 60755 13105 ;
    LAYER M1 ;
      RECT 60935 335 61185 3865 ;
    LAYER M1 ;
      RECT 60935 6215 61185 9745 ;
    LAYER M1 ;
      RECT 61365 335 61615 3865 ;
    LAYER M1 ;
      RECT 61365 4115 61615 5125 ;
    LAYER M1 ;
      RECT 61365 6215 61615 9745 ;
    LAYER M1 ;
      RECT 61365 9995 61615 11005 ;
    LAYER M1 ;
      RECT 61365 12095 61615 13105 ;
    LAYER M1 ;
      RECT 61795 335 62045 3865 ;
    LAYER M1 ;
      RECT 61795 6215 62045 9745 ;
    LAYER M1 ;
      RECT 62225 335 62475 3865 ;
    LAYER M1 ;
      RECT 62225 4115 62475 5125 ;
    LAYER M1 ;
      RECT 62225 6215 62475 9745 ;
    LAYER M1 ;
      RECT 62225 9995 62475 11005 ;
    LAYER M1 ;
      RECT 62225 12095 62475 13105 ;
    LAYER M1 ;
      RECT 62655 335 62905 3865 ;
    LAYER M1 ;
      RECT 62655 6215 62905 9745 ;
    LAYER M1 ;
      RECT 63085 335 63335 3865 ;
    LAYER M1 ;
      RECT 63085 4115 63335 5125 ;
    LAYER M1 ;
      RECT 63085 6215 63335 9745 ;
    LAYER M1 ;
      RECT 63085 9995 63335 11005 ;
    LAYER M1 ;
      RECT 63085 12095 63335 13105 ;
    LAYER M1 ;
      RECT 63515 335 63765 3865 ;
    LAYER M1 ;
      RECT 63515 6215 63765 9745 ;
    LAYER M1 ;
      RECT 63945 335 64195 3865 ;
    LAYER M1 ;
      RECT 63945 4115 64195 5125 ;
    LAYER M1 ;
      RECT 63945 6215 64195 9745 ;
    LAYER M1 ;
      RECT 63945 9995 64195 11005 ;
    LAYER M1 ;
      RECT 63945 12095 64195 13105 ;
    LAYER M1 ;
      RECT 64375 335 64625 3865 ;
    LAYER M1 ;
      RECT 64375 6215 64625 9745 ;
    LAYER M2 ;
      RECT 1120 280 64240 560 ;
    LAYER M2 ;
      RECT 1120 4480 64240 4760 ;
    LAYER M2 ;
      RECT 690 700 64670 980 ;
    LAYER M2 ;
      RECT 1120 6160 64240 6440 ;
    LAYER M2 ;
      RECT 1120 10360 64240 10640 ;
    LAYER M2 ;
      RECT 1120 12460 64240 12740 ;
    LAYER M2 ;
      RECT 690 6580 64670 6860 ;
    LAYER V1 ;
      RECT 54525 335 54695 505 ;
    LAYER V1 ;
      RECT 54525 4535 54695 4705 ;
    LAYER V1 ;
      RECT 54525 6215 54695 6385 ;
    LAYER V1 ;
      RECT 54525 10415 54695 10585 ;
    LAYER V1 ;
      RECT 54525 12515 54695 12685 ;
    LAYER V1 ;
      RECT 55385 335 55555 505 ;
    LAYER V1 ;
      RECT 55385 4535 55555 4705 ;
    LAYER V1 ;
      RECT 55385 6215 55555 6385 ;
    LAYER V1 ;
      RECT 55385 10415 55555 10585 ;
    LAYER V1 ;
      RECT 55385 12515 55555 12685 ;
    LAYER V1 ;
      RECT 56245 335 56415 505 ;
    LAYER V1 ;
      RECT 56245 4535 56415 4705 ;
    LAYER V1 ;
      RECT 56245 6215 56415 6385 ;
    LAYER V1 ;
      RECT 56245 10415 56415 10585 ;
    LAYER V1 ;
      RECT 56245 12515 56415 12685 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12515 1375 12685 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12515 2235 12685 ;
    LAYER V1 ;
      RECT 57105 335 57275 505 ;
    LAYER V1 ;
      RECT 57105 4535 57275 4705 ;
    LAYER V1 ;
      RECT 57105 6215 57275 6385 ;
    LAYER V1 ;
      RECT 57105 10415 57275 10585 ;
    LAYER V1 ;
      RECT 57105 12515 57275 12685 ;
    LAYER V1 ;
      RECT 57965 335 58135 505 ;
    LAYER V1 ;
      RECT 57965 4535 58135 4705 ;
    LAYER V1 ;
      RECT 57965 6215 58135 6385 ;
    LAYER V1 ;
      RECT 57965 10415 58135 10585 ;
    LAYER V1 ;
      RECT 57965 12515 58135 12685 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12515 3095 12685 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12515 3955 12685 ;
    LAYER V1 ;
      RECT 58825 335 58995 505 ;
    LAYER V1 ;
      RECT 58825 4535 58995 4705 ;
    LAYER V1 ;
      RECT 58825 6215 58995 6385 ;
    LAYER V1 ;
      RECT 58825 10415 58995 10585 ;
    LAYER V1 ;
      RECT 58825 12515 58995 12685 ;
    LAYER V1 ;
      RECT 59685 335 59855 505 ;
    LAYER V1 ;
      RECT 59685 4535 59855 4705 ;
    LAYER V1 ;
      RECT 59685 6215 59855 6385 ;
    LAYER V1 ;
      RECT 59685 10415 59855 10585 ;
    LAYER V1 ;
      RECT 59685 12515 59855 12685 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12515 4815 12685 ;
    LAYER V1 ;
      RECT 60545 335 60715 505 ;
    LAYER V1 ;
      RECT 60545 4535 60715 4705 ;
    LAYER V1 ;
      RECT 60545 6215 60715 6385 ;
    LAYER V1 ;
      RECT 60545 10415 60715 10585 ;
    LAYER V1 ;
      RECT 60545 12515 60715 12685 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12515 5675 12685 ;
    LAYER V1 ;
      RECT 61405 335 61575 505 ;
    LAYER V1 ;
      RECT 61405 4535 61575 4705 ;
    LAYER V1 ;
      RECT 61405 6215 61575 6385 ;
    LAYER V1 ;
      RECT 61405 10415 61575 10585 ;
    LAYER V1 ;
      RECT 61405 12515 61575 12685 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12515 6535 12685 ;
    LAYER V1 ;
      RECT 62265 335 62435 505 ;
    LAYER V1 ;
      RECT 62265 4535 62435 4705 ;
    LAYER V1 ;
      RECT 62265 6215 62435 6385 ;
    LAYER V1 ;
      RECT 62265 10415 62435 10585 ;
    LAYER V1 ;
      RECT 62265 12515 62435 12685 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12515 7395 12685 ;
    LAYER V1 ;
      RECT 63125 335 63295 505 ;
    LAYER V1 ;
      RECT 63125 4535 63295 4705 ;
    LAYER V1 ;
      RECT 63125 6215 63295 6385 ;
    LAYER V1 ;
      RECT 63125 10415 63295 10585 ;
    LAYER V1 ;
      RECT 63125 12515 63295 12685 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12515 8255 12685 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12515 9115 12685 ;
    LAYER V1 ;
      RECT 63985 335 64155 505 ;
    LAYER V1 ;
      RECT 63985 4535 64155 4705 ;
    LAYER V1 ;
      RECT 63985 6215 64155 6385 ;
    LAYER V1 ;
      RECT 63985 10415 64155 10585 ;
    LAYER V1 ;
      RECT 63985 12515 64155 12685 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6215 9975 6385 ;
    LAYER V1 ;
      RECT 9805 10415 9975 10585 ;
    LAYER V1 ;
      RECT 9805 12515 9975 12685 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6215 10835 6385 ;
    LAYER V1 ;
      RECT 10665 10415 10835 10585 ;
    LAYER V1 ;
      RECT 10665 12515 10835 12685 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6215 11695 6385 ;
    LAYER V1 ;
      RECT 11525 10415 11695 10585 ;
    LAYER V1 ;
      RECT 11525 12515 11695 12685 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6215 12555 6385 ;
    LAYER V1 ;
      RECT 12385 10415 12555 10585 ;
    LAYER V1 ;
      RECT 12385 12515 12555 12685 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6215 13415 6385 ;
    LAYER V1 ;
      RECT 13245 10415 13415 10585 ;
    LAYER V1 ;
      RECT 13245 12515 13415 12685 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6215 14275 6385 ;
    LAYER V1 ;
      RECT 14105 10415 14275 10585 ;
    LAYER V1 ;
      RECT 14105 12515 14275 12685 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6215 15135 6385 ;
    LAYER V1 ;
      RECT 14965 10415 15135 10585 ;
    LAYER V1 ;
      RECT 14965 12515 15135 12685 ;
    LAYER V1 ;
      RECT 15825 335 15995 505 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6215 15995 6385 ;
    LAYER V1 ;
      RECT 15825 10415 15995 10585 ;
    LAYER V1 ;
      RECT 15825 12515 15995 12685 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6215 16855 6385 ;
    LAYER V1 ;
      RECT 16685 10415 16855 10585 ;
    LAYER V1 ;
      RECT 16685 12515 16855 12685 ;
    LAYER V1 ;
      RECT 17545 335 17715 505 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6215 17715 6385 ;
    LAYER V1 ;
      RECT 17545 10415 17715 10585 ;
    LAYER V1 ;
      RECT 17545 12515 17715 12685 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6215 18575 6385 ;
    LAYER V1 ;
      RECT 18405 10415 18575 10585 ;
    LAYER V1 ;
      RECT 18405 12515 18575 12685 ;
    LAYER V1 ;
      RECT 19265 335 19435 505 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6215 19435 6385 ;
    LAYER V1 ;
      RECT 19265 10415 19435 10585 ;
    LAYER V1 ;
      RECT 19265 12515 19435 12685 ;
    LAYER V1 ;
      RECT 20125 335 20295 505 ;
    LAYER V1 ;
      RECT 20125 4535 20295 4705 ;
    LAYER V1 ;
      RECT 20125 6215 20295 6385 ;
    LAYER V1 ;
      RECT 20125 10415 20295 10585 ;
    LAYER V1 ;
      RECT 20125 12515 20295 12685 ;
    LAYER V1 ;
      RECT 20985 335 21155 505 ;
    LAYER V1 ;
      RECT 20985 4535 21155 4705 ;
    LAYER V1 ;
      RECT 20985 6215 21155 6385 ;
    LAYER V1 ;
      RECT 20985 10415 21155 10585 ;
    LAYER V1 ;
      RECT 20985 12515 21155 12685 ;
    LAYER V1 ;
      RECT 21845 335 22015 505 ;
    LAYER V1 ;
      RECT 21845 4535 22015 4705 ;
    LAYER V1 ;
      RECT 21845 6215 22015 6385 ;
    LAYER V1 ;
      RECT 21845 10415 22015 10585 ;
    LAYER V1 ;
      RECT 21845 12515 22015 12685 ;
    LAYER V1 ;
      RECT 22705 335 22875 505 ;
    LAYER V1 ;
      RECT 22705 4535 22875 4705 ;
    LAYER V1 ;
      RECT 22705 6215 22875 6385 ;
    LAYER V1 ;
      RECT 22705 10415 22875 10585 ;
    LAYER V1 ;
      RECT 22705 12515 22875 12685 ;
    LAYER V1 ;
      RECT 23565 335 23735 505 ;
    LAYER V1 ;
      RECT 23565 4535 23735 4705 ;
    LAYER V1 ;
      RECT 23565 6215 23735 6385 ;
    LAYER V1 ;
      RECT 23565 10415 23735 10585 ;
    LAYER V1 ;
      RECT 23565 12515 23735 12685 ;
    LAYER V1 ;
      RECT 24425 335 24595 505 ;
    LAYER V1 ;
      RECT 24425 4535 24595 4705 ;
    LAYER V1 ;
      RECT 24425 6215 24595 6385 ;
    LAYER V1 ;
      RECT 24425 10415 24595 10585 ;
    LAYER V1 ;
      RECT 24425 12515 24595 12685 ;
    LAYER V1 ;
      RECT 25285 335 25455 505 ;
    LAYER V1 ;
      RECT 25285 4535 25455 4705 ;
    LAYER V1 ;
      RECT 25285 6215 25455 6385 ;
    LAYER V1 ;
      RECT 25285 10415 25455 10585 ;
    LAYER V1 ;
      RECT 25285 12515 25455 12685 ;
    LAYER V1 ;
      RECT 26145 335 26315 505 ;
    LAYER V1 ;
      RECT 26145 4535 26315 4705 ;
    LAYER V1 ;
      RECT 26145 6215 26315 6385 ;
    LAYER V1 ;
      RECT 26145 10415 26315 10585 ;
    LAYER V1 ;
      RECT 26145 12515 26315 12685 ;
    LAYER V1 ;
      RECT 27005 335 27175 505 ;
    LAYER V1 ;
      RECT 27005 4535 27175 4705 ;
    LAYER V1 ;
      RECT 27005 6215 27175 6385 ;
    LAYER V1 ;
      RECT 27005 10415 27175 10585 ;
    LAYER V1 ;
      RECT 27005 12515 27175 12685 ;
    LAYER V1 ;
      RECT 27865 335 28035 505 ;
    LAYER V1 ;
      RECT 27865 4535 28035 4705 ;
    LAYER V1 ;
      RECT 27865 6215 28035 6385 ;
    LAYER V1 ;
      RECT 27865 10415 28035 10585 ;
    LAYER V1 ;
      RECT 27865 12515 28035 12685 ;
    LAYER V1 ;
      RECT 28725 335 28895 505 ;
    LAYER V1 ;
      RECT 28725 4535 28895 4705 ;
    LAYER V1 ;
      RECT 28725 6215 28895 6385 ;
    LAYER V1 ;
      RECT 28725 10415 28895 10585 ;
    LAYER V1 ;
      RECT 28725 12515 28895 12685 ;
    LAYER V1 ;
      RECT 29585 335 29755 505 ;
    LAYER V1 ;
      RECT 29585 4535 29755 4705 ;
    LAYER V1 ;
      RECT 29585 6215 29755 6385 ;
    LAYER V1 ;
      RECT 29585 10415 29755 10585 ;
    LAYER V1 ;
      RECT 29585 12515 29755 12685 ;
    LAYER V1 ;
      RECT 30445 335 30615 505 ;
    LAYER V1 ;
      RECT 30445 4535 30615 4705 ;
    LAYER V1 ;
      RECT 30445 6215 30615 6385 ;
    LAYER V1 ;
      RECT 30445 10415 30615 10585 ;
    LAYER V1 ;
      RECT 30445 12515 30615 12685 ;
    LAYER V1 ;
      RECT 31305 335 31475 505 ;
    LAYER V1 ;
      RECT 31305 4535 31475 4705 ;
    LAYER V1 ;
      RECT 31305 6215 31475 6385 ;
    LAYER V1 ;
      RECT 31305 10415 31475 10585 ;
    LAYER V1 ;
      RECT 31305 12515 31475 12685 ;
    LAYER V1 ;
      RECT 32165 335 32335 505 ;
    LAYER V1 ;
      RECT 32165 4535 32335 4705 ;
    LAYER V1 ;
      RECT 32165 6215 32335 6385 ;
    LAYER V1 ;
      RECT 32165 10415 32335 10585 ;
    LAYER V1 ;
      RECT 32165 12515 32335 12685 ;
    LAYER V1 ;
      RECT 33025 335 33195 505 ;
    LAYER V1 ;
      RECT 33025 4535 33195 4705 ;
    LAYER V1 ;
      RECT 33025 6215 33195 6385 ;
    LAYER V1 ;
      RECT 33025 10415 33195 10585 ;
    LAYER V1 ;
      RECT 33025 12515 33195 12685 ;
    LAYER V1 ;
      RECT 33885 335 34055 505 ;
    LAYER V1 ;
      RECT 33885 4535 34055 4705 ;
    LAYER V1 ;
      RECT 33885 6215 34055 6385 ;
    LAYER V1 ;
      RECT 33885 10415 34055 10585 ;
    LAYER V1 ;
      RECT 33885 12515 34055 12685 ;
    LAYER V1 ;
      RECT 34745 335 34915 505 ;
    LAYER V1 ;
      RECT 34745 4535 34915 4705 ;
    LAYER V1 ;
      RECT 34745 6215 34915 6385 ;
    LAYER V1 ;
      RECT 34745 10415 34915 10585 ;
    LAYER V1 ;
      RECT 34745 12515 34915 12685 ;
    LAYER V1 ;
      RECT 35605 335 35775 505 ;
    LAYER V1 ;
      RECT 35605 4535 35775 4705 ;
    LAYER V1 ;
      RECT 35605 6215 35775 6385 ;
    LAYER V1 ;
      RECT 35605 10415 35775 10585 ;
    LAYER V1 ;
      RECT 35605 12515 35775 12685 ;
    LAYER V1 ;
      RECT 36465 335 36635 505 ;
    LAYER V1 ;
      RECT 36465 4535 36635 4705 ;
    LAYER V1 ;
      RECT 36465 6215 36635 6385 ;
    LAYER V1 ;
      RECT 36465 10415 36635 10585 ;
    LAYER V1 ;
      RECT 36465 12515 36635 12685 ;
    LAYER V1 ;
      RECT 37325 335 37495 505 ;
    LAYER V1 ;
      RECT 37325 4535 37495 4705 ;
    LAYER V1 ;
      RECT 37325 6215 37495 6385 ;
    LAYER V1 ;
      RECT 37325 10415 37495 10585 ;
    LAYER V1 ;
      RECT 37325 12515 37495 12685 ;
    LAYER V1 ;
      RECT 38185 335 38355 505 ;
    LAYER V1 ;
      RECT 38185 4535 38355 4705 ;
    LAYER V1 ;
      RECT 38185 6215 38355 6385 ;
    LAYER V1 ;
      RECT 38185 10415 38355 10585 ;
    LAYER V1 ;
      RECT 38185 12515 38355 12685 ;
    LAYER V1 ;
      RECT 39045 335 39215 505 ;
    LAYER V1 ;
      RECT 39045 4535 39215 4705 ;
    LAYER V1 ;
      RECT 39045 6215 39215 6385 ;
    LAYER V1 ;
      RECT 39045 10415 39215 10585 ;
    LAYER V1 ;
      RECT 39045 12515 39215 12685 ;
    LAYER V1 ;
      RECT 39905 335 40075 505 ;
    LAYER V1 ;
      RECT 39905 4535 40075 4705 ;
    LAYER V1 ;
      RECT 39905 6215 40075 6385 ;
    LAYER V1 ;
      RECT 39905 10415 40075 10585 ;
    LAYER V1 ;
      RECT 39905 12515 40075 12685 ;
    LAYER V1 ;
      RECT 40765 335 40935 505 ;
    LAYER V1 ;
      RECT 40765 4535 40935 4705 ;
    LAYER V1 ;
      RECT 40765 6215 40935 6385 ;
    LAYER V1 ;
      RECT 40765 10415 40935 10585 ;
    LAYER V1 ;
      RECT 40765 12515 40935 12685 ;
    LAYER V1 ;
      RECT 41625 335 41795 505 ;
    LAYER V1 ;
      RECT 41625 4535 41795 4705 ;
    LAYER V1 ;
      RECT 41625 6215 41795 6385 ;
    LAYER V1 ;
      RECT 41625 10415 41795 10585 ;
    LAYER V1 ;
      RECT 41625 12515 41795 12685 ;
    LAYER V1 ;
      RECT 42485 335 42655 505 ;
    LAYER V1 ;
      RECT 42485 4535 42655 4705 ;
    LAYER V1 ;
      RECT 42485 6215 42655 6385 ;
    LAYER V1 ;
      RECT 42485 10415 42655 10585 ;
    LAYER V1 ;
      RECT 42485 12515 42655 12685 ;
    LAYER V1 ;
      RECT 43345 335 43515 505 ;
    LAYER V1 ;
      RECT 43345 4535 43515 4705 ;
    LAYER V1 ;
      RECT 43345 6215 43515 6385 ;
    LAYER V1 ;
      RECT 43345 10415 43515 10585 ;
    LAYER V1 ;
      RECT 43345 12515 43515 12685 ;
    LAYER V1 ;
      RECT 44205 335 44375 505 ;
    LAYER V1 ;
      RECT 44205 4535 44375 4705 ;
    LAYER V1 ;
      RECT 44205 6215 44375 6385 ;
    LAYER V1 ;
      RECT 44205 10415 44375 10585 ;
    LAYER V1 ;
      RECT 44205 12515 44375 12685 ;
    LAYER V1 ;
      RECT 45065 335 45235 505 ;
    LAYER V1 ;
      RECT 45065 4535 45235 4705 ;
    LAYER V1 ;
      RECT 45065 6215 45235 6385 ;
    LAYER V1 ;
      RECT 45065 10415 45235 10585 ;
    LAYER V1 ;
      RECT 45065 12515 45235 12685 ;
    LAYER V1 ;
      RECT 45925 335 46095 505 ;
    LAYER V1 ;
      RECT 45925 4535 46095 4705 ;
    LAYER V1 ;
      RECT 45925 6215 46095 6385 ;
    LAYER V1 ;
      RECT 45925 10415 46095 10585 ;
    LAYER V1 ;
      RECT 45925 12515 46095 12685 ;
    LAYER V1 ;
      RECT 46785 335 46955 505 ;
    LAYER V1 ;
      RECT 46785 4535 46955 4705 ;
    LAYER V1 ;
      RECT 46785 6215 46955 6385 ;
    LAYER V1 ;
      RECT 46785 10415 46955 10585 ;
    LAYER V1 ;
      RECT 46785 12515 46955 12685 ;
    LAYER V1 ;
      RECT 47645 335 47815 505 ;
    LAYER V1 ;
      RECT 47645 4535 47815 4705 ;
    LAYER V1 ;
      RECT 47645 6215 47815 6385 ;
    LAYER V1 ;
      RECT 47645 10415 47815 10585 ;
    LAYER V1 ;
      RECT 47645 12515 47815 12685 ;
    LAYER V1 ;
      RECT 48505 335 48675 505 ;
    LAYER V1 ;
      RECT 48505 4535 48675 4705 ;
    LAYER V1 ;
      RECT 48505 6215 48675 6385 ;
    LAYER V1 ;
      RECT 48505 10415 48675 10585 ;
    LAYER V1 ;
      RECT 48505 12515 48675 12685 ;
    LAYER V1 ;
      RECT 49365 335 49535 505 ;
    LAYER V1 ;
      RECT 49365 4535 49535 4705 ;
    LAYER V1 ;
      RECT 49365 6215 49535 6385 ;
    LAYER V1 ;
      RECT 49365 10415 49535 10585 ;
    LAYER V1 ;
      RECT 49365 12515 49535 12685 ;
    LAYER V1 ;
      RECT 50225 335 50395 505 ;
    LAYER V1 ;
      RECT 50225 4535 50395 4705 ;
    LAYER V1 ;
      RECT 50225 6215 50395 6385 ;
    LAYER V1 ;
      RECT 50225 10415 50395 10585 ;
    LAYER V1 ;
      RECT 50225 12515 50395 12685 ;
    LAYER V1 ;
      RECT 51085 335 51255 505 ;
    LAYER V1 ;
      RECT 51085 4535 51255 4705 ;
    LAYER V1 ;
      RECT 51085 6215 51255 6385 ;
    LAYER V1 ;
      RECT 51085 10415 51255 10585 ;
    LAYER V1 ;
      RECT 51085 12515 51255 12685 ;
    LAYER V1 ;
      RECT 51945 335 52115 505 ;
    LAYER V1 ;
      RECT 51945 4535 52115 4705 ;
    LAYER V1 ;
      RECT 51945 6215 52115 6385 ;
    LAYER V1 ;
      RECT 51945 10415 52115 10585 ;
    LAYER V1 ;
      RECT 51945 12515 52115 12685 ;
    LAYER V1 ;
      RECT 52805 335 52975 505 ;
    LAYER V1 ;
      RECT 52805 4535 52975 4705 ;
    LAYER V1 ;
      RECT 52805 6215 52975 6385 ;
    LAYER V1 ;
      RECT 52805 10415 52975 10585 ;
    LAYER V1 ;
      RECT 52805 12515 52975 12685 ;
    LAYER V1 ;
      RECT 53665 335 53835 505 ;
    LAYER V1 ;
      RECT 53665 4535 53835 4705 ;
    LAYER V1 ;
      RECT 53665 6215 53835 6385 ;
    LAYER V1 ;
      RECT 53665 10415 53835 10585 ;
    LAYER V1 ;
      RECT 53665 12515 53835 12685 ;
    LAYER V1 ;
      RECT 54955 755 55125 925 ;
    LAYER V1 ;
      RECT 54955 6635 55125 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 55815 755 55985 925 ;
    LAYER V1 ;
      RECT 55815 6635 55985 6805 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 56675 755 56845 925 ;
    LAYER V1 ;
      RECT 56675 6635 56845 6805 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 57535 755 57705 925 ;
    LAYER V1 ;
      RECT 57535 6635 57705 6805 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 58395 755 58565 925 ;
    LAYER V1 ;
      RECT 58395 6635 58565 6805 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 59255 755 59425 925 ;
    LAYER V1 ;
      RECT 59255 6635 59425 6805 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 60115 755 60285 925 ;
    LAYER V1 ;
      RECT 60115 6635 60285 6805 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 60975 755 61145 925 ;
    LAYER V1 ;
      RECT 60975 6635 61145 6805 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 61835 755 62005 925 ;
    LAYER V1 ;
      RECT 61835 6635 62005 6805 ;
    LAYER V1 ;
      RECT 62695 755 62865 925 ;
    LAYER V1 ;
      RECT 62695 6635 62865 6805 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 63555 755 63725 925 ;
    LAYER V1 ;
      RECT 63555 6635 63725 6805 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 9375 6635 9545 6805 ;
    LAYER V1 ;
      RECT 64415 755 64585 925 ;
    LAYER V1 ;
      RECT 64415 6635 64585 6805 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 10235 6635 10405 6805 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11095 6635 11265 6805 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 11955 6635 12125 6805 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 12815 6635 12985 6805 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 13675 6635 13845 6805 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 14535 6635 14705 6805 ;
    LAYER V1 ;
      RECT 15395 755 15565 925 ;
    LAYER V1 ;
      RECT 15395 6635 15565 6805 ;
    LAYER V1 ;
      RECT 16255 755 16425 925 ;
    LAYER V1 ;
      RECT 16255 6635 16425 6805 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17115 6635 17285 6805 ;
    LAYER V1 ;
      RECT 17975 755 18145 925 ;
    LAYER V1 ;
      RECT 17975 6635 18145 6805 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 18835 6635 19005 6805 ;
    LAYER V1 ;
      RECT 19695 755 19865 925 ;
    LAYER V1 ;
      RECT 19695 6635 19865 6805 ;
    LAYER V1 ;
      RECT 20555 755 20725 925 ;
    LAYER V1 ;
      RECT 20555 6635 20725 6805 ;
    LAYER V1 ;
      RECT 21415 755 21585 925 ;
    LAYER V1 ;
      RECT 21415 6635 21585 6805 ;
    LAYER V1 ;
      RECT 22275 755 22445 925 ;
    LAYER V1 ;
      RECT 22275 6635 22445 6805 ;
    LAYER V1 ;
      RECT 23135 755 23305 925 ;
    LAYER V1 ;
      RECT 23135 6635 23305 6805 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 23995 6635 24165 6805 ;
    LAYER V1 ;
      RECT 24855 755 25025 925 ;
    LAYER V1 ;
      RECT 24855 6635 25025 6805 ;
    LAYER V1 ;
      RECT 25715 755 25885 925 ;
    LAYER V1 ;
      RECT 25715 6635 25885 6805 ;
    LAYER V1 ;
      RECT 26575 755 26745 925 ;
    LAYER V1 ;
      RECT 26575 6635 26745 6805 ;
    LAYER V1 ;
      RECT 27435 755 27605 925 ;
    LAYER V1 ;
      RECT 27435 6635 27605 6805 ;
    LAYER V1 ;
      RECT 28295 755 28465 925 ;
    LAYER V1 ;
      RECT 28295 6635 28465 6805 ;
    LAYER V1 ;
      RECT 29155 755 29325 925 ;
    LAYER V1 ;
      RECT 29155 6635 29325 6805 ;
    LAYER V1 ;
      RECT 30015 755 30185 925 ;
    LAYER V1 ;
      RECT 30015 6635 30185 6805 ;
    LAYER V1 ;
      RECT 30875 755 31045 925 ;
    LAYER V1 ;
      RECT 30875 6635 31045 6805 ;
    LAYER V1 ;
      RECT 31735 755 31905 925 ;
    LAYER V1 ;
      RECT 31735 6635 31905 6805 ;
    LAYER V1 ;
      RECT 32595 755 32765 925 ;
    LAYER V1 ;
      RECT 32595 6635 32765 6805 ;
    LAYER V1 ;
      RECT 33455 755 33625 925 ;
    LAYER V1 ;
      RECT 33455 6635 33625 6805 ;
    LAYER V1 ;
      RECT 34315 755 34485 925 ;
    LAYER V1 ;
      RECT 34315 6635 34485 6805 ;
    LAYER V1 ;
      RECT 35175 755 35345 925 ;
    LAYER V1 ;
      RECT 35175 6635 35345 6805 ;
    LAYER V1 ;
      RECT 36035 755 36205 925 ;
    LAYER V1 ;
      RECT 36035 6635 36205 6805 ;
    LAYER V1 ;
      RECT 36895 755 37065 925 ;
    LAYER V1 ;
      RECT 36895 6635 37065 6805 ;
    LAYER V1 ;
      RECT 37755 755 37925 925 ;
    LAYER V1 ;
      RECT 37755 6635 37925 6805 ;
    LAYER V1 ;
      RECT 38615 755 38785 925 ;
    LAYER V1 ;
      RECT 38615 6635 38785 6805 ;
    LAYER V1 ;
      RECT 39475 755 39645 925 ;
    LAYER V1 ;
      RECT 39475 6635 39645 6805 ;
    LAYER V1 ;
      RECT 40335 755 40505 925 ;
    LAYER V1 ;
      RECT 40335 6635 40505 6805 ;
    LAYER V1 ;
      RECT 41195 755 41365 925 ;
    LAYER V1 ;
      RECT 41195 6635 41365 6805 ;
    LAYER V1 ;
      RECT 42055 755 42225 925 ;
    LAYER V1 ;
      RECT 42055 6635 42225 6805 ;
    LAYER V1 ;
      RECT 42915 755 43085 925 ;
    LAYER V1 ;
      RECT 42915 6635 43085 6805 ;
    LAYER V1 ;
      RECT 43775 755 43945 925 ;
    LAYER V1 ;
      RECT 43775 6635 43945 6805 ;
    LAYER V1 ;
      RECT 44635 755 44805 925 ;
    LAYER V1 ;
      RECT 44635 6635 44805 6805 ;
    LAYER V1 ;
      RECT 45495 755 45665 925 ;
    LAYER V1 ;
      RECT 45495 6635 45665 6805 ;
    LAYER V1 ;
      RECT 46355 755 46525 925 ;
    LAYER V1 ;
      RECT 46355 6635 46525 6805 ;
    LAYER V1 ;
      RECT 47215 755 47385 925 ;
    LAYER V1 ;
      RECT 47215 6635 47385 6805 ;
    LAYER V1 ;
      RECT 48075 755 48245 925 ;
    LAYER V1 ;
      RECT 48075 6635 48245 6805 ;
    LAYER V1 ;
      RECT 48935 755 49105 925 ;
    LAYER V1 ;
      RECT 48935 6635 49105 6805 ;
    LAYER V1 ;
      RECT 49795 755 49965 925 ;
    LAYER V1 ;
      RECT 49795 6635 49965 6805 ;
    LAYER V1 ;
      RECT 50655 755 50825 925 ;
    LAYER V1 ;
      RECT 50655 6635 50825 6805 ;
    LAYER V1 ;
      RECT 51515 755 51685 925 ;
    LAYER V1 ;
      RECT 51515 6635 51685 6805 ;
    LAYER V1 ;
      RECT 52375 755 52545 925 ;
    LAYER V1 ;
      RECT 52375 6635 52545 6805 ;
    LAYER V1 ;
      RECT 53235 755 53405 925 ;
    LAYER V1 ;
      RECT 53235 6635 53405 6805 ;
    LAYER V1 ;
      RECT 54095 755 54265 925 ;
    LAYER V1 ;
      RECT 54095 6635 54265 6805 ;
    LAYER V2 ;
      RECT 32175 345 32325 495 ;
    LAYER V2 ;
      RECT 32175 6225 32325 6375 ;
    LAYER V2 ;
      RECT 32605 4545 32755 4695 ;
    LAYER V2 ;
      RECT 32605 10425 32755 10575 ;
    LAYER V2 ;
      RECT 33035 765 33185 915 ;
    LAYER V2 ;
      RECT 33035 6645 33185 6795 ;
    LAYER V2 ;
      RECT 33035 12525 33185 12675 ;
  END
END NMOS_S_12565100_X74_Y2
