# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.41000 BY  11.69000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT  0.000000  0.000000  5.430000  0.330000 ;
        RECT  0.000000  0.330000  0.330000  0.750000 ;
        RECT  0.000000  0.750000  5.430000  0.890000 ;
        RECT  0.000000  0.890000  0.330000  1.310000 ;
        RECT  0.000000  1.310000  5.430000  1.450000 ;
        RECT  0.000000  1.450000  0.330000  1.870000 ;
        RECT  0.000000  1.870000  5.430000  2.010000 ;
        RECT  0.000000  2.010000  0.330000  2.430000 ;
        RECT  0.000000  2.430000  5.430000  2.570000 ;
        RECT  0.000000  2.570000  0.330000  2.990000 ;
        RECT  0.000000  2.990000  5.430000  3.130000 ;
        RECT  0.000000  3.130000  0.330000  3.550000 ;
        RECT  0.000000  3.550000  5.430000  3.690000 ;
        RECT  0.000000  3.690000  0.330000  4.110000 ;
        RECT  0.000000  4.110000  5.430000  4.250000 ;
        RECT  0.000000  4.250000  0.330000  4.670000 ;
        RECT  0.000000  4.670000  5.430000  4.810000 ;
        RECT  0.000000  4.810000  0.330000  5.230000 ;
        RECT  0.000000  5.230000  5.430000  5.370000 ;
        RECT  0.000000  5.370000  0.330000  5.570000 ;
        RECT  0.000000  6.120000  0.330000  6.320000 ;
        RECT  0.000000  6.320000  5.430000  6.460000 ;
        RECT  0.000000  6.460000  0.330000  6.880000 ;
        RECT  0.000000  6.880000  5.430000  7.020000 ;
        RECT  0.000000  7.020000  0.330000  7.440000 ;
        RECT  0.000000  7.440000  5.430000  7.580000 ;
        RECT  0.000000  7.580000  0.330000  8.000000 ;
        RECT  0.000000  8.000000  5.430000  8.140000 ;
        RECT  0.000000  8.140000  0.330000  8.560000 ;
        RECT  0.000000  8.560000  5.430000  8.700000 ;
        RECT  0.000000  8.700000  0.330000  9.120000 ;
        RECT  0.000000  9.120000  5.430000  9.260000 ;
        RECT  0.000000  9.260000  0.330000  9.680000 ;
        RECT  0.000000  9.680000  5.430000  9.820000 ;
        RECT  0.000000  9.820000  0.330000 10.240000 ;
        RECT  0.000000 10.240000  5.430000 10.380000 ;
        RECT  0.000000 10.380000  0.330000 10.800000 ;
        RECT  0.000000 10.800000  5.430000 10.940000 ;
        RECT  0.000000 10.940000  0.330000 11.360000 ;
        RECT  0.000000 11.360000  5.430000 11.690000 ;
        RECT  5.980000  0.000000 11.410000  0.330000 ;
        RECT  5.980000  0.750000 11.410000  0.890000 ;
        RECT  5.980000  1.310000 11.410000  1.450000 ;
        RECT  5.980000  1.870000 11.410000  2.010000 ;
        RECT  5.980000  2.430000 11.410000  2.570000 ;
        RECT  5.980000  2.990000 11.410000  3.130000 ;
        RECT  5.980000  3.550000 11.410000  3.690000 ;
        RECT  5.980000  4.110000 11.410000  4.250000 ;
        RECT  5.980000  4.670000 11.410000  4.810000 ;
        RECT  5.980000  5.230000 11.410000  5.370000 ;
        RECT  5.980000  6.320000 11.410000  6.460000 ;
        RECT  5.980000  6.880000 11.410000  7.020000 ;
        RECT  5.980000  7.440000 11.410000  7.580000 ;
        RECT  5.980000  8.000000 11.410000  8.140000 ;
        RECT  5.980000  8.560000 11.410000  8.700000 ;
        RECT  5.980000  9.120000 11.410000  9.260000 ;
        RECT  5.980000  9.680000 11.410000  9.820000 ;
        RECT  5.980000 10.240000 11.410000 10.380000 ;
        RECT  5.980000 10.800000 11.410000 10.940000 ;
        RECT  5.980000 11.360000 11.410000 11.690000 ;
        RECT 11.080000  0.330000 11.410000  0.750000 ;
        RECT 11.080000  0.890000 11.410000  1.310000 ;
        RECT 11.080000  1.450000 11.410000  1.870000 ;
        RECT 11.080000  2.010000 11.410000  2.430000 ;
        RECT 11.080000  2.570000 11.410000  2.990000 ;
        RECT 11.080000  3.130000 11.410000  3.550000 ;
        RECT 11.080000  3.690000 11.410000  4.110000 ;
        RECT 11.080000  4.250000 11.410000  4.670000 ;
        RECT 11.080000  4.810000 11.410000  5.230000 ;
        RECT 11.080000  5.370000 11.410000  5.570000 ;
        RECT 11.080000  6.120000 11.410000  6.320000 ;
        RECT 11.080000  6.460000 11.410000  6.880000 ;
        RECT 11.080000  7.020000 11.410000  7.440000 ;
        RECT 11.080000  7.580000 11.410000  8.000000 ;
        RECT 11.080000  8.140000 11.410000  8.560000 ;
        RECT 11.080000  8.700000 11.410000  9.120000 ;
        RECT 11.080000  9.260000 11.410000  9.680000 ;
        RECT 11.080000  9.820000 11.410000 10.240000 ;
        RECT 11.080000 10.380000 11.410000 10.800000 ;
        RECT 11.080000 10.940000 11.410000 11.360000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT 0.000000  5.710000 11.410000  5.980000 ;
        RECT 0.470000  0.470000 10.940000  0.610000 ;
        RECT 0.470000  1.030000 10.940000  1.170000 ;
        RECT 0.470000  1.590000 10.940000  1.730000 ;
        RECT 0.470000  2.150000 10.940000  2.290000 ;
        RECT 0.470000  2.710000 10.940000  2.850000 ;
        RECT 0.470000  3.270000 10.940000  3.410000 ;
        RECT 0.470000  3.830000 10.940000  3.970000 ;
        RECT 0.470000  4.390000 10.940000  4.530000 ;
        RECT 0.470000  4.950000 10.940000  5.090000 ;
        RECT 0.470000  6.600000 10.940000  6.740000 ;
        RECT 0.470000  7.160000 10.940000  7.300000 ;
        RECT 0.470000  7.720000 10.940000  7.860000 ;
        RECT 0.470000  8.280000 10.940000  8.420000 ;
        RECT 0.470000  8.840000 10.940000  8.980000 ;
        RECT 0.470000  9.400000 10.940000  9.540000 ;
        RECT 0.470000  9.960000 10.940000 10.100000 ;
        RECT 0.470000 10.520000 10.940000 10.660000 ;
        RECT 0.470000 11.080000 10.940000 11.220000 ;
        RECT 5.570000  0.000000  5.840000  0.470000 ;
        RECT 5.570000  0.610000  5.840000  1.030000 ;
        RECT 5.570000  1.170000  5.840000  1.590000 ;
        RECT 5.570000  1.730000  5.840000  2.150000 ;
        RECT 5.570000  2.290000  5.840000  2.710000 ;
        RECT 5.570000  2.850000  5.840000  3.270000 ;
        RECT 5.570000  3.410000  5.840000  3.830000 ;
        RECT 5.570000  3.970000  5.840000  4.390000 ;
        RECT 5.570000  4.530000  5.840000  4.950000 ;
        RECT 5.570000  5.090000  5.840000  5.710000 ;
        RECT 5.570000  5.980000  5.840000  6.600000 ;
        RECT 5.570000  6.740000  5.840000  7.160000 ;
        RECT 5.570000  7.300000  5.840000  7.720000 ;
        RECT 5.570000  7.860000  5.840000  8.280000 ;
        RECT 5.570000  8.420000  5.840000  8.840000 ;
        RECT 5.570000  8.980000  5.840000  9.400000 ;
        RECT 5.570000  9.540000  5.840000  9.960000 ;
        RECT 5.570000 10.100000  5.840000 10.520000 ;
        RECT 5.570000 10.660000  5.840000 11.080000 ;
        RECT 5.570000 11.220000  5.840000 11.690000 ;
    END
  END C1
  PIN MET3
    PORT
      LAYER met3 ;
        RECT 0.000000 0.000000 11.410000 11.690000 ;
    END
  END MET3
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 5.880000 6.445000 5.985000 6.690000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.860000 ;
      RECT  0.000000  0.860000  5.400000  1.030000 ;
      RECT  0.000000  1.030000  0.330000  1.560000 ;
      RECT  0.000000  1.560000  5.400000  1.730000 ;
      RECT  0.000000  1.730000  0.330000  2.260000 ;
      RECT  0.000000  2.260000  5.400000  2.430000 ;
      RECT  0.000000  2.430000  0.330000  2.960000 ;
      RECT  0.000000  2.960000  5.400000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.660000 ;
      RECT  0.000000  3.660000  5.400000  3.830000 ;
      RECT  0.000000  3.830000  0.330000  4.360000 ;
      RECT  0.000000  4.360000  5.400000  4.530000 ;
      RECT  0.000000  4.530000  0.330000  5.060000 ;
      RECT  0.000000  5.060000  5.400000  5.230000 ;
      RECT  0.000000  5.230000  0.330000  5.760000 ;
      RECT  0.000000  5.760000  5.400000  5.930000 ;
      RECT  0.000000  5.930000  0.330000  6.460000 ;
      RECT  0.000000  6.460000  5.400000  6.630000 ;
      RECT  0.000000  6.630000  0.330000  7.160000 ;
      RECT  0.000000  7.160000  5.400000  7.330000 ;
      RECT  0.000000  7.330000  0.330000  7.860000 ;
      RECT  0.000000  7.860000  5.400000  8.030000 ;
      RECT  0.000000  8.030000  0.330000  8.560000 ;
      RECT  0.000000  8.560000  5.400000  8.730000 ;
      RECT  0.000000  8.730000  0.330000  9.260000 ;
      RECT  0.000000  9.260000  5.400000  9.430000 ;
      RECT  0.000000  9.430000  0.330000  9.960000 ;
      RECT  0.000000  9.960000  5.400000 10.130000 ;
      RECT  0.000000 10.130000  0.330000 10.660000 ;
      RECT  0.000000 10.660000  5.400000 10.830000 ;
      RECT  0.000000 10.830000  0.330000 11.360000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.500000  0.510000 10.905000  0.680000 ;
      RECT  0.500000  1.210000 10.905000  1.380000 ;
      RECT  0.500000  1.910000 10.905000  2.080000 ;
      RECT  0.500000  2.610000 10.905000  2.780000 ;
      RECT  0.500000  3.310000 10.905000  3.480000 ;
      RECT  0.500000  4.010000 10.905000  4.180000 ;
      RECT  0.500000  4.710000 10.905000  4.880000 ;
      RECT  0.500000  5.410000 10.905000  5.580000 ;
      RECT  0.500000  6.110000 10.905000  6.280000 ;
      RECT  0.500000  6.810000 10.905000  6.980000 ;
      RECT  0.500000  7.510000 10.905000  7.680000 ;
      RECT  0.500000  8.210000 10.905000  8.380000 ;
      RECT  0.500000  8.910000 10.905000  9.080000 ;
      RECT  0.500000  9.610000 10.905000  9.780000 ;
      RECT  0.500000 10.310000 10.905000 10.480000 ;
      RECT  0.500000 11.010000 10.905000 11.180000 ;
      RECT  5.570000  0.680000  5.840000  1.210000 ;
      RECT  5.570000  1.380000  5.840000  1.910000 ;
      RECT  5.570000  2.080000  5.840000  2.610000 ;
      RECT  5.570000  2.780000  5.840000  3.310000 ;
      RECT  5.570000  3.480000  5.840000  4.010000 ;
      RECT  5.570000  4.180000  5.840000  4.710000 ;
      RECT  5.570000  4.880000  5.840000  5.410000 ;
      RECT  5.570000  5.580000  5.840000  6.110000 ;
      RECT  5.570000  6.280000  5.840000  6.810000 ;
      RECT  5.570000  6.980000  5.840000  7.510000 ;
      RECT  5.570000  7.680000  5.840000  8.210000 ;
      RECT  5.570000  8.380000  5.840000  8.910000 ;
      RECT  5.570000  9.080000  5.840000  9.610000 ;
      RECT  5.570000  9.780000  5.840000 10.310000 ;
      RECT  5.570000 10.480000  5.840000 11.010000 ;
      RECT  6.010000  0.860000 11.410000  1.030000 ;
      RECT  6.010000  1.560000 11.410000  1.730000 ;
      RECT  6.010000  2.260000 11.410000  2.430000 ;
      RECT  6.010000  2.960000 11.410000  3.130000 ;
      RECT  6.010000  3.660000 11.410000  3.830000 ;
      RECT  6.010000  4.360000 11.410000  4.530000 ;
      RECT  6.010000  5.060000 11.410000  5.230000 ;
      RECT  6.010000  5.760000 11.410000  5.930000 ;
      RECT  6.010000  6.460000 11.410000  6.630000 ;
      RECT  6.010000  7.160000 11.410000  7.330000 ;
      RECT  6.010000  7.860000 11.410000  8.030000 ;
      RECT  6.010000  8.560000 11.410000  8.730000 ;
      RECT  6.010000  9.260000 11.410000  9.430000 ;
      RECT  6.010000  9.960000 11.410000 10.130000 ;
      RECT  6.010000 10.660000 11.410000 10.830000 ;
      RECT 11.080000  0.330000 11.410000  0.860000 ;
      RECT 11.080000  1.030000 11.410000  1.560000 ;
      RECT 11.080000  1.730000 11.410000  2.260000 ;
      RECT 11.080000  2.430000 11.410000  2.960000 ;
      RECT 11.080000  3.130000 11.410000  3.660000 ;
      RECT 11.080000  3.830000 11.410000  4.360000 ;
      RECT 11.080000  4.530000 11.410000  5.060000 ;
      RECT 11.080000  5.230000 11.410000  5.760000 ;
      RECT 11.080000  5.930000 11.410000  6.460000 ;
      RECT 11.080000  6.630000 11.410000  7.160000 ;
      RECT 11.080000  7.330000 11.410000  7.860000 ;
      RECT 11.080000  8.030000 11.410000  8.560000 ;
      RECT 11.080000  8.730000 11.410000  9.260000 ;
      RECT 11.080000  9.430000 11.410000  9.960000 ;
      RECT 11.080000 10.130000 11.410000 10.660000 ;
      RECT 11.080000 10.830000 11.410000 11.360000 ;
    LAYER mcon ;
      RECT  0.080000  0.580000  0.250000  0.750000 ;
      RECT  0.080000  0.940000  0.250000  1.110000 ;
      RECT  0.080000  1.300000  0.250000  1.470000 ;
      RECT  0.080000  1.660000  0.250000  1.830000 ;
      RECT  0.080000  2.020000  0.250000  2.190000 ;
      RECT  0.080000  2.380000  0.250000  2.550000 ;
      RECT  0.080000  2.740000  0.250000  2.910000 ;
      RECT  0.080000  3.100000  0.250000  3.270000 ;
      RECT  0.080000  3.460000  0.250000  3.630000 ;
      RECT  0.080000  3.820000  0.250000  3.990000 ;
      RECT  0.080000  4.180000  0.250000  4.350000 ;
      RECT  0.080000  4.540000  0.250000  4.710000 ;
      RECT  0.080000  4.900000  0.250000  5.070000 ;
      RECT  0.080000  5.260000  0.250000  5.430000 ;
      RECT  0.080000  6.260000  0.250000  6.430000 ;
      RECT  0.080000  6.620000  0.250000  6.790000 ;
      RECT  0.080000  6.980000  0.250000  7.150000 ;
      RECT  0.080000  7.340000  0.250000  7.510000 ;
      RECT  0.080000  7.700000  0.250000  7.870000 ;
      RECT  0.080000  8.060000  0.250000  8.230000 ;
      RECT  0.080000  8.420000  0.250000  8.590000 ;
      RECT  0.080000  8.780000  0.250000  8.950000 ;
      RECT  0.080000  9.140000  0.250000  9.310000 ;
      RECT  0.080000  9.500000  0.250000  9.670000 ;
      RECT  0.080000  9.860000  0.250000 10.030000 ;
      RECT  0.080000 10.220000  0.250000 10.390000 ;
      RECT  0.080000 10.580000  0.250000 10.750000 ;
      RECT  0.080000 10.940000  0.250000 11.110000 ;
      RECT  0.400000  0.080000  0.570000  0.250000 ;
      RECT  0.400000 11.440000  0.570000 11.610000 ;
      RECT  0.760000  0.080000  0.930000  0.250000 ;
      RECT  0.760000 11.440000  0.930000 11.610000 ;
      RECT  1.120000  0.080000  1.290000  0.250000 ;
      RECT  1.120000 11.440000  1.290000 11.610000 ;
      RECT  1.480000  0.080000  1.650000  0.250000 ;
      RECT  1.480000 11.440000  1.650000 11.610000 ;
      RECT  1.840000  0.080000  2.010000  0.250000 ;
      RECT  1.840000 11.440000  2.010000 11.610000 ;
      RECT  2.200000  0.080000  2.370000  0.250000 ;
      RECT  2.200000 11.440000  2.370000 11.610000 ;
      RECT  2.560000  0.080000  2.730000  0.250000 ;
      RECT  2.560000 11.440000  2.730000 11.610000 ;
      RECT  2.920000  0.080000  3.090000  0.250000 ;
      RECT  2.920000 11.440000  3.090000 11.610000 ;
      RECT  3.280000  0.080000  3.450000  0.250000 ;
      RECT  3.280000 11.440000  3.450000 11.610000 ;
      RECT  3.640000  0.080000  3.810000  0.250000 ;
      RECT  3.640000 11.440000  3.810000 11.610000 ;
      RECT  4.000000  0.080000  4.170000  0.250000 ;
      RECT  4.000000 11.440000  4.170000 11.610000 ;
      RECT  4.360000  0.080000  4.530000  0.250000 ;
      RECT  4.360000 11.440000  4.530000 11.610000 ;
      RECT  4.720000  0.080000  4.890000  0.250000 ;
      RECT  4.720000 11.440000  4.890000 11.610000 ;
      RECT  5.080000  0.080000  5.250000  0.250000 ;
      RECT  5.080000 11.440000  5.250000 11.610000 ;
      RECT  5.440000  0.080000  5.610000  0.250000 ;
      RECT  5.440000 11.440000  5.610000 11.610000 ;
      RECT  5.620000  0.590000  5.790000  0.760000 ;
      RECT  5.620000  0.950000  5.790000  1.120000 ;
      RECT  5.620000  1.310000  5.790000  1.480000 ;
      RECT  5.620000  1.670000  5.790000  1.840000 ;
      RECT  5.620000  2.030000  5.790000  2.200000 ;
      RECT  5.620000  2.390000  5.790000  2.560000 ;
      RECT  5.620000  2.750000  5.790000  2.920000 ;
      RECT  5.620000  3.110000  5.790000  3.280000 ;
      RECT  5.620000  3.470000  5.790000  3.640000 ;
      RECT  5.620000  3.830000  5.790000  4.000000 ;
      RECT  5.620000  4.190000  5.790000  4.360000 ;
      RECT  5.620000  4.550000  5.790000  4.720000 ;
      RECT  5.620000  4.910000  5.790000  5.080000 ;
      RECT  5.620000  5.270000  5.790000  5.440000 ;
      RECT  5.620000  6.250000  5.790000  6.420000 ;
      RECT  5.620000  6.610000  5.790000  6.780000 ;
      RECT  5.620000  6.970000  5.790000  7.140000 ;
      RECT  5.620000  7.330000  5.790000  7.500000 ;
      RECT  5.620000  7.690000  5.790000  7.860000 ;
      RECT  5.620000  8.050000  5.790000  8.220000 ;
      RECT  5.620000  8.410000  5.790000  8.580000 ;
      RECT  5.620000  8.770000  5.790000  8.940000 ;
      RECT  5.620000  9.130000  5.790000  9.300000 ;
      RECT  5.620000  9.490000  5.790000  9.660000 ;
      RECT  5.620000  9.850000  5.790000 10.020000 ;
      RECT  5.620000 10.210000  5.790000 10.380000 ;
      RECT  5.620000 10.570000  5.790000 10.740000 ;
      RECT  5.620000 10.930000  5.790000 11.100000 ;
      RECT  5.800000  0.080000  5.970000  0.250000 ;
      RECT  5.800000 11.440000  5.970000 11.610000 ;
      RECT  6.160000  0.080000  6.330000  0.250000 ;
      RECT  6.160000 11.440000  6.330000 11.610000 ;
      RECT  6.520000  0.080000  6.690000  0.250000 ;
      RECT  6.520000 11.440000  6.690000 11.610000 ;
      RECT  6.880000  0.080000  7.050000  0.250000 ;
      RECT  6.880000 11.440000  7.050000 11.610000 ;
      RECT  7.240000  0.080000  7.410000  0.250000 ;
      RECT  7.240000 11.440000  7.410000 11.610000 ;
      RECT  7.600000  0.080000  7.770000  0.250000 ;
      RECT  7.600000 11.440000  7.770000 11.610000 ;
      RECT  7.960000  0.080000  8.130000  0.250000 ;
      RECT  7.960000 11.440000  8.130000 11.610000 ;
      RECT  8.320000  0.080000  8.490000  0.250000 ;
      RECT  8.320000 11.440000  8.490000 11.610000 ;
      RECT  8.680000  0.080000  8.850000  0.250000 ;
      RECT  8.680000 11.440000  8.850000 11.610000 ;
      RECT  9.040000  0.080000  9.210000  0.250000 ;
      RECT  9.040000 11.440000  9.210000 11.610000 ;
      RECT  9.400000  0.080000  9.570000  0.250000 ;
      RECT  9.400000 11.440000  9.570000 11.610000 ;
      RECT  9.760000  0.080000  9.930000  0.250000 ;
      RECT  9.760000 11.440000  9.930000 11.610000 ;
      RECT 10.120000  0.080000 10.290000  0.250000 ;
      RECT 10.120000 11.440000 10.290000 11.610000 ;
      RECT 10.480000  0.080000 10.650000  0.250000 ;
      RECT 10.480000 11.440000 10.650000 11.610000 ;
      RECT 10.840000  0.080000 11.010000  0.250000 ;
      RECT 10.840000 11.440000 11.010000 11.610000 ;
      RECT 11.160000  0.580000 11.330000  0.750000 ;
      RECT 11.160000  0.940000 11.330000  1.110000 ;
      RECT 11.160000  1.300000 11.330000  1.470000 ;
      RECT 11.160000  1.660000 11.330000  1.830000 ;
      RECT 11.160000  2.020000 11.330000  2.190000 ;
      RECT 11.160000  2.380000 11.330000  2.550000 ;
      RECT 11.160000  2.740000 11.330000  2.910000 ;
      RECT 11.160000  3.100000 11.330000  3.270000 ;
      RECT 11.160000  3.460000 11.330000  3.630000 ;
      RECT 11.160000  3.820000 11.330000  3.990000 ;
      RECT 11.160000  4.180000 11.330000  4.350000 ;
      RECT 11.160000  4.540000 11.330000  4.710000 ;
      RECT 11.160000  4.900000 11.330000  5.070000 ;
      RECT 11.160000  5.260000 11.330000  5.430000 ;
      RECT 11.160000  6.260000 11.330000  6.430000 ;
      RECT 11.160000  6.620000 11.330000  6.790000 ;
      RECT 11.160000  6.980000 11.330000  7.150000 ;
      RECT 11.160000  7.340000 11.330000  7.510000 ;
      RECT 11.160000  7.700000 11.330000  7.870000 ;
      RECT 11.160000  8.060000 11.330000  8.230000 ;
      RECT 11.160000  8.420000 11.330000  8.590000 ;
      RECT 11.160000  8.780000 11.330000  8.950000 ;
      RECT 11.160000  9.140000 11.330000  9.310000 ;
      RECT 11.160000  9.500000 11.330000  9.670000 ;
      RECT 11.160000  9.860000 11.330000 10.030000 ;
      RECT 11.160000 10.220000 11.330000 10.390000 ;
      RECT 11.160000 10.580000 11.330000 10.750000 ;
      RECT 11.160000 10.940000 11.330000 11.110000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.330000  0.330000 11.360000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.500000  0.470000  0.640000  5.685000 ;
      RECT  0.500000  5.685000 10.910000  6.005000 ;
      RECT  0.500000  6.005000  0.640000 11.220000 ;
      RECT  0.780000  0.330000  0.920000  5.545000 ;
      RECT  0.780000  6.145000  0.920000 11.360000 ;
      RECT  1.060000  0.470000  1.200000  5.685000 ;
      RECT  1.060000  6.005000  1.200000 11.220000 ;
      RECT  1.340000  0.330000  1.480000  5.545000 ;
      RECT  1.340000  6.145000  1.480000 11.360000 ;
      RECT  1.620000  0.470000  1.760000  5.685000 ;
      RECT  1.620000  6.005000  1.760000 11.220000 ;
      RECT  1.900000  0.330000  2.040000  5.545000 ;
      RECT  1.900000  6.145000  2.040000 11.360000 ;
      RECT  2.180000  0.470000  2.320000  5.685000 ;
      RECT  2.180000  6.005000  2.320000 11.220000 ;
      RECT  2.460000  0.330000  2.600000  5.545000 ;
      RECT  2.460000  6.145000  2.600000 11.360000 ;
      RECT  2.740000  0.470000  2.880000  5.685000 ;
      RECT  2.740000  6.005000  2.880000 11.220000 ;
      RECT  3.020000  0.330000  3.160000  5.545000 ;
      RECT  3.020000  6.145000  3.160000 11.360000 ;
      RECT  3.300000  0.470000  3.440000  5.685000 ;
      RECT  3.300000  6.005000  3.440000 11.220000 ;
      RECT  3.580000  0.330000  3.720000  5.545000 ;
      RECT  3.580000  6.145000  3.720000 11.360000 ;
      RECT  3.860000  0.470000  4.000000  5.685000 ;
      RECT  3.860000  6.005000  4.000000 11.220000 ;
      RECT  4.140000  0.330000  4.280000  5.545000 ;
      RECT  4.140000  6.145000  4.280000 11.360000 ;
      RECT  4.420000  0.470000  4.560000  5.685000 ;
      RECT  4.420000  6.005000  4.560000 11.220000 ;
      RECT  4.700000  0.330000  4.840000  5.545000 ;
      RECT  4.700000  6.145000  4.840000 11.360000 ;
      RECT  4.980000  0.470000  5.120000  5.685000 ;
      RECT  4.980000  6.005000  5.120000 11.220000 ;
      RECT  5.260000  0.330000  5.400000  5.545000 ;
      RECT  5.260000  6.145000  5.400000 11.360000 ;
      RECT  5.570000  0.470000  5.840000  5.685000 ;
      RECT  5.570000  6.005000  5.840000 11.220000 ;
      RECT  6.010000  0.330000  6.150000  5.545000 ;
      RECT  6.010000  6.145000  6.150000 11.360000 ;
      RECT  6.290000  0.470000  6.430000  5.685000 ;
      RECT  6.290000  6.005000  6.430000 11.220000 ;
      RECT  6.570000  0.330000  6.710000  5.545000 ;
      RECT  6.570000  6.145000  6.710000 11.360000 ;
      RECT  6.850000  0.470000  6.990000  5.685000 ;
      RECT  6.850000  6.005000  6.990000 11.220000 ;
      RECT  7.130000  0.330000  7.270000  5.545000 ;
      RECT  7.130000  6.145000  7.270000 11.360000 ;
      RECT  7.410000  0.470000  7.550000  5.685000 ;
      RECT  7.410000  6.005000  7.550000 11.220000 ;
      RECT  7.690000  0.330000  7.830000  5.545000 ;
      RECT  7.690000  6.145000  7.830000 11.360000 ;
      RECT  7.970000  0.470000  8.110000  5.685000 ;
      RECT  7.970000  6.005000  8.110000 11.220000 ;
      RECT  8.250000  0.330000  8.390000  5.545000 ;
      RECT  8.250000  6.145000  8.390000 11.360000 ;
      RECT  8.530000  0.470000  8.670000  5.685000 ;
      RECT  8.530000  6.005000  8.670000 11.220000 ;
      RECT  8.810000  0.330000  8.950000  5.545000 ;
      RECT  8.810000  6.145000  8.950000 11.360000 ;
      RECT  9.090000  0.470000  9.230000  5.685000 ;
      RECT  9.090000  6.005000  9.230000 11.220000 ;
      RECT  9.370000  0.330000  9.510000  5.545000 ;
      RECT  9.370000  6.145000  9.510000 11.360000 ;
      RECT  9.650000  0.470000  9.790000  5.685000 ;
      RECT  9.650000  6.005000  9.790000 11.220000 ;
      RECT  9.930000  0.330000 10.070000  5.545000 ;
      RECT  9.930000  6.145000 10.070000 11.360000 ;
      RECT 10.210000  0.470000 10.350000  5.685000 ;
      RECT 10.210000  6.005000 10.350000 11.220000 ;
      RECT 10.490000  0.330000 10.630000  5.545000 ;
      RECT 10.490000  6.145000 10.630000 11.360000 ;
      RECT 10.770000  0.470000 10.910000  5.685000 ;
      RECT 10.770000  6.005000 10.910000 11.220000 ;
      RECT 11.080000  0.330000 11.410000 11.360000 ;
    LAYER via ;
      RECT  0.035000  0.280000  0.295000  0.540000 ;
      RECT  0.035000  0.600000  0.295000  0.860000 ;
      RECT  0.035000  0.920000  0.295000  1.180000 ;
      RECT  0.035000  1.240000  0.295000  1.500000 ;
      RECT  0.035000  1.560000  0.295000  1.820000 ;
      RECT  0.035000  1.880000  0.295000  2.140000 ;
      RECT  0.035000  2.200000  0.295000  2.460000 ;
      RECT  0.035000  2.520000  0.295000  2.780000 ;
      RECT  0.035000  2.840000  0.295000  3.100000 ;
      RECT  0.035000  3.160000  0.295000  3.420000 ;
      RECT  0.035000  3.480000  0.295000  3.740000 ;
      RECT  0.035000  3.800000  0.295000  4.060000 ;
      RECT  0.035000  4.120000  0.295000  4.380000 ;
      RECT  0.035000  4.440000  0.295000  4.700000 ;
      RECT  0.035000  4.760000  0.295000  5.020000 ;
      RECT  0.035000  5.080000  0.295000  5.340000 ;
      RECT  0.035000  6.350000  0.295000  6.610000 ;
      RECT  0.035000  6.670000  0.295000  6.930000 ;
      RECT  0.035000  6.990000  0.295000  7.250000 ;
      RECT  0.035000  7.310000  0.295000  7.570000 ;
      RECT  0.035000  7.630000  0.295000  7.890000 ;
      RECT  0.035000  7.950000  0.295000  8.210000 ;
      RECT  0.035000  8.270000  0.295000  8.530000 ;
      RECT  0.035000  8.590000  0.295000  8.850000 ;
      RECT  0.035000  8.910000  0.295000  9.170000 ;
      RECT  0.035000  9.230000  0.295000  9.490000 ;
      RECT  0.035000  9.550000  0.295000  9.810000 ;
      RECT  0.035000  9.870000  0.295000 10.130000 ;
      RECT  0.035000 10.190000  0.295000 10.450000 ;
      RECT  0.035000 10.510000  0.295000 10.770000 ;
      RECT  0.035000 10.830000  0.295000 11.090000 ;
      RECT  0.035000 11.150000  0.295000 11.410000 ;
      RECT  0.440000  0.035000  0.700000  0.295000 ;
      RECT  0.440000 11.395000  0.700000 11.655000 ;
      RECT  0.760000  0.035000  1.020000  0.295000 ;
      RECT  0.760000  5.715000  1.020000  5.975000 ;
      RECT  0.760000 11.395000  1.020000 11.655000 ;
      RECT  1.080000  0.035000  1.340000  0.295000 ;
      RECT  1.080000  5.715000  1.340000  5.975000 ;
      RECT  1.080000 11.395000  1.340000 11.655000 ;
      RECT  1.400000  0.035000  1.660000  0.295000 ;
      RECT  1.400000  5.715000  1.660000  5.975000 ;
      RECT  1.400000 11.395000  1.660000 11.655000 ;
      RECT  1.720000  0.035000  1.980000  0.295000 ;
      RECT  1.720000  5.715000  1.980000  5.975000 ;
      RECT  1.720000 11.395000  1.980000 11.655000 ;
      RECT  2.040000  0.035000  2.300000  0.295000 ;
      RECT  2.040000  5.715000  2.300000  5.975000 ;
      RECT  2.040000 11.395000  2.300000 11.655000 ;
      RECT  2.360000  0.035000  2.620000  0.295000 ;
      RECT  2.360000  5.715000  2.620000  5.975000 ;
      RECT  2.360000 11.395000  2.620000 11.655000 ;
      RECT  2.680000  0.035000  2.940000  0.295000 ;
      RECT  2.680000  5.715000  2.940000  5.975000 ;
      RECT  2.680000 11.395000  2.940000 11.655000 ;
      RECT  3.000000  0.035000  3.260000  0.295000 ;
      RECT  3.000000  5.715000  3.260000  5.975000 ;
      RECT  3.000000 11.395000  3.260000 11.655000 ;
      RECT  3.320000  0.035000  3.580000  0.295000 ;
      RECT  3.320000  5.715000  3.580000  5.975000 ;
      RECT  3.320000 11.395000  3.580000 11.655000 ;
      RECT  3.640000  0.035000  3.900000  0.295000 ;
      RECT  3.640000  5.715000  3.900000  5.975000 ;
      RECT  3.640000 11.395000  3.900000 11.655000 ;
      RECT  3.960000  0.035000  4.220000  0.295000 ;
      RECT  3.960000  5.715000  4.220000  5.975000 ;
      RECT  3.960000 11.395000  4.220000 11.655000 ;
      RECT  4.280000  0.035000  4.540000  0.295000 ;
      RECT  4.280000  5.715000  4.540000  5.975000 ;
      RECT  4.280000 11.395000  4.540000 11.655000 ;
      RECT  4.600000  0.035000  4.860000  0.295000 ;
      RECT  4.600000  5.715000  4.860000  5.975000 ;
      RECT  4.600000 11.395000  4.860000 11.655000 ;
      RECT  4.920000  0.035000  5.180000  0.295000 ;
      RECT  4.920000  5.715000  5.180000  5.975000 ;
      RECT  4.920000 11.395000  5.180000 11.655000 ;
      RECT  5.240000  5.715000  5.500000  5.975000 ;
      RECT  5.575000  0.505000  5.835000  0.765000 ;
      RECT  5.575000  0.825000  5.835000  1.085000 ;
      RECT  5.575000  1.145000  5.835000  1.405000 ;
      RECT  5.575000  1.465000  5.835000  1.725000 ;
      RECT  5.575000  1.785000  5.835000  2.045000 ;
      RECT  5.575000  2.105000  5.835000  2.365000 ;
      RECT  5.575000  2.425000  5.835000  2.685000 ;
      RECT  5.575000  2.745000  5.835000  3.005000 ;
      RECT  5.575000  3.065000  5.835000  3.325000 ;
      RECT  5.575000  3.385000  5.835000  3.645000 ;
      RECT  5.575000  3.705000  5.835000  3.965000 ;
      RECT  5.575000  4.025000  5.835000  4.285000 ;
      RECT  5.575000  4.345000  5.835000  4.605000 ;
      RECT  5.575000  4.665000  5.835000  4.925000 ;
      RECT  5.575000  4.985000  5.835000  5.245000 ;
      RECT  5.575000  5.305000  5.835000  5.565000 ;
      RECT  5.575000  6.125000  5.835000  6.385000 ;
      RECT  5.575000  6.445000  5.835000  6.705000 ;
      RECT  5.575000  6.765000  5.835000  7.025000 ;
      RECT  5.575000  7.085000  5.835000  7.345000 ;
      RECT  5.575000  7.405000  5.835000  7.665000 ;
      RECT  5.575000  7.725000  5.835000  7.985000 ;
      RECT  5.575000  8.045000  5.835000  8.305000 ;
      RECT  5.575000  8.365000  5.835000  8.625000 ;
      RECT  5.575000  8.685000  5.835000  8.945000 ;
      RECT  5.575000  9.005000  5.835000  9.265000 ;
      RECT  5.575000  9.325000  5.835000  9.585000 ;
      RECT  5.575000  9.645000  5.835000  9.905000 ;
      RECT  5.575000  9.965000  5.835000 10.225000 ;
      RECT  5.575000 10.285000  5.835000 10.545000 ;
      RECT  5.575000 10.605000  5.835000 10.865000 ;
      RECT  5.575000 10.925000  5.835000 11.185000 ;
      RECT  5.910000  5.715000  6.170000  5.975000 ;
      RECT  6.230000  0.035000  6.490000  0.295000 ;
      RECT  6.230000  5.715000  6.490000  5.975000 ;
      RECT  6.230000 11.395000  6.490000 11.655000 ;
      RECT  6.550000  0.035000  6.810000  0.295000 ;
      RECT  6.550000  5.715000  6.810000  5.975000 ;
      RECT  6.550000 11.395000  6.810000 11.655000 ;
      RECT  6.870000  0.035000  7.130000  0.295000 ;
      RECT  6.870000  5.715000  7.130000  5.975000 ;
      RECT  6.870000 11.395000  7.130000 11.655000 ;
      RECT  7.190000  0.035000  7.450000  0.295000 ;
      RECT  7.190000  5.715000  7.450000  5.975000 ;
      RECT  7.190000 11.395000  7.450000 11.655000 ;
      RECT  7.510000  0.035000  7.770000  0.295000 ;
      RECT  7.510000  5.715000  7.770000  5.975000 ;
      RECT  7.510000 11.395000  7.770000 11.655000 ;
      RECT  7.830000  0.035000  8.090000  0.295000 ;
      RECT  7.830000  5.715000  8.090000  5.975000 ;
      RECT  7.830000 11.395000  8.090000 11.655000 ;
      RECT  8.150000  0.035000  8.410000  0.295000 ;
      RECT  8.150000  5.715000  8.410000  5.975000 ;
      RECT  8.150000 11.395000  8.410000 11.655000 ;
      RECT  8.470000  0.035000  8.730000  0.295000 ;
      RECT  8.470000  5.715000  8.730000  5.975000 ;
      RECT  8.470000 11.395000  8.730000 11.655000 ;
      RECT  8.790000  0.035000  9.050000  0.295000 ;
      RECT  8.790000  5.715000  9.050000  5.975000 ;
      RECT  8.790000 11.395000  9.050000 11.655000 ;
      RECT  9.110000  0.035000  9.370000  0.295000 ;
      RECT  9.110000  5.715000  9.370000  5.975000 ;
      RECT  9.110000 11.395000  9.370000 11.655000 ;
      RECT  9.430000  0.035000  9.690000  0.295000 ;
      RECT  9.430000  5.715000  9.690000  5.975000 ;
      RECT  9.430000 11.395000  9.690000 11.655000 ;
      RECT  9.750000  0.035000 10.010000  0.295000 ;
      RECT  9.750000  5.715000 10.010000  5.975000 ;
      RECT  9.750000 11.395000 10.010000 11.655000 ;
      RECT 10.070000  0.035000 10.330000  0.295000 ;
      RECT 10.070000  5.715000 10.330000  5.975000 ;
      RECT 10.070000 11.395000 10.330000 11.655000 ;
      RECT 10.390000  0.035000 10.650000  0.295000 ;
      RECT 10.390000  5.715000 10.650000  5.975000 ;
      RECT 10.390000 11.395000 10.650000 11.655000 ;
      RECT 10.710000  0.035000 10.970000  0.295000 ;
      RECT 10.710000 11.395000 10.970000 11.655000 ;
      RECT 11.115000  0.280000 11.375000  0.540000 ;
      RECT 11.115000  0.600000 11.375000  0.860000 ;
      RECT 11.115000  0.920000 11.375000  1.180000 ;
      RECT 11.115000  1.240000 11.375000  1.500000 ;
      RECT 11.115000  1.560000 11.375000  1.820000 ;
      RECT 11.115000  1.880000 11.375000  2.140000 ;
      RECT 11.115000  2.200000 11.375000  2.460000 ;
      RECT 11.115000  2.520000 11.375000  2.780000 ;
      RECT 11.115000  2.840000 11.375000  3.100000 ;
      RECT 11.115000  3.160000 11.375000  3.420000 ;
      RECT 11.115000  3.480000 11.375000  3.740000 ;
      RECT 11.115000  3.800000 11.375000  4.060000 ;
      RECT 11.115000  4.120000 11.375000  4.380000 ;
      RECT 11.115000  4.440000 11.375000  4.700000 ;
      RECT 11.115000  4.760000 11.375000  5.020000 ;
      RECT 11.115000  5.080000 11.375000  5.340000 ;
      RECT 11.115000  6.350000 11.375000  6.610000 ;
      RECT 11.115000  6.670000 11.375000  6.930000 ;
      RECT 11.115000  6.990000 11.375000  7.250000 ;
      RECT 11.115000  7.310000 11.375000  7.570000 ;
      RECT 11.115000  7.630000 11.375000  7.890000 ;
      RECT 11.115000  7.950000 11.375000  8.210000 ;
      RECT 11.115000  8.270000 11.375000  8.530000 ;
      RECT 11.115000  8.590000 11.375000  8.850000 ;
      RECT 11.115000  8.910000 11.375000  9.170000 ;
      RECT 11.115000  9.230000 11.375000  9.490000 ;
      RECT 11.115000  9.550000 11.375000  9.810000 ;
      RECT 11.115000  9.870000 11.375000 10.130000 ;
      RECT 11.115000 10.190000 11.375000 10.450000 ;
      RECT 11.115000 10.510000 11.375000 10.770000 ;
      RECT 11.115000 10.830000 11.375000 11.090000 ;
      RECT 11.115000 11.150000 11.375000 11.410000 ;
  END
END sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3
END LIBRARY
