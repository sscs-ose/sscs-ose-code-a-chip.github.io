MACRO SCM_NMOS_B_85279373_X2_Y4
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_85279373_X2_Y4 0 0 ;
  SIZE 8600 BY 25200 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 24220 7050 24500 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3730 260 4010 22420 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4160 680 4440 18640 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4590 1100 4870 19060 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 4115 1845 5125 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 9995 1845 11005 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 15875 1845 16885 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 21755 1845 22765 ;
    LAYER M1 ;
      RECT 1595 23855 1845 24865 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 4115 3565 5125 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 9995 3565 11005 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 15875 3565 16885 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 21755 3565 22765 ;
    LAYER M1 ;
      RECT 3315 23855 3565 24865 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 4115 5285 5125 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 9995 5285 11005 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 15875 5285 16885 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 21755 5285 22765 ;
    LAYER M1 ;
      RECT 5035 23855 5285 24865 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 4115 7005 5125 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 9995 7005 11005 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 6755 15875 7005 16885 ;
    LAYER M1 ;
      RECT 6755 17975 7005 21505 ;
    LAYER M1 ;
      RECT 6755 21755 7005 22765 ;
    LAYER M1 ;
      RECT 6755 23855 7005 24865 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 7615 17975 7865 21505 ;
    LAYER M2 ;
      RECT 1550 4480 7050 4760 ;
    LAYER M2 ;
      RECT 1550 280 7050 560 ;
    LAYER M2 ;
      RECT 3270 700 5330 980 ;
    LAYER M2 ;
      RECT 690 1120 7910 1400 ;
    LAYER M2 ;
      RECT 1550 10360 7050 10640 ;
    LAYER M2 ;
      RECT 3270 6160 5330 6440 ;
    LAYER M2 ;
      RECT 1550 6580 7050 6860 ;
    LAYER M2 ;
      RECT 690 7000 7910 7280 ;
    LAYER M2 ;
      RECT 1550 16240 7050 16520 ;
    LAYER M2 ;
      RECT 1550 12040 7050 12320 ;
    LAYER M2 ;
      RECT 3270 12460 5330 12740 ;
    LAYER M2 ;
      RECT 690 12880 7910 13160 ;
    LAYER M2 ;
      RECT 1550 22120 7050 22400 ;
    LAYER M2 ;
      RECT 3270 17920 5330 18200 ;
    LAYER M2 ;
      RECT 1550 18340 7050 18620 ;
    LAYER M2 ;
      RECT 690 18760 7910 19040 ;
    LAYER V1 ;
      RECT 6795 335 6965 505 ;
    LAYER V1 ;
      RECT 6795 4535 6965 4705 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 10415 6965 10585 ;
    LAYER V1 ;
      RECT 6795 12095 6965 12265 ;
    LAYER V1 ;
      RECT 6795 16295 6965 16465 ;
    LAYER V1 ;
      RECT 6795 18395 6965 18565 ;
    LAYER V1 ;
      RECT 6795 22175 6965 22345 ;
    LAYER V1 ;
      RECT 6795 24275 6965 24445 ;
    LAYER V1 ;
      RECT 1635 335 1805 505 ;
    LAYER V1 ;
      RECT 1635 4535 1805 4705 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 10415 1805 10585 ;
    LAYER V1 ;
      RECT 1635 12095 1805 12265 ;
    LAYER V1 ;
      RECT 1635 16295 1805 16465 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 22175 1805 22345 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 4535 5245 4705 ;
    LAYER V1 ;
      RECT 5075 6215 5245 6385 ;
    LAYER V1 ;
      RECT 5075 10415 5245 10585 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 16295 5245 16465 ;
    LAYER V1 ;
      RECT 5075 17975 5245 18145 ;
    LAYER V1 ;
      RECT 5075 22175 5245 22345 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 4535 3525 4705 ;
    LAYER V1 ;
      RECT 3355 6215 3525 6385 ;
    LAYER V1 ;
      RECT 3355 10415 3525 10585 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 16295 3525 16465 ;
    LAYER V1 ;
      RECT 3355 17975 3525 18145 ;
    LAYER V1 ;
      RECT 3355 22175 3525 22345 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 775 7055 945 7225 ;
    LAYER V1 ;
      RECT 775 12935 945 13105 ;
    LAYER V1 ;
      RECT 775 18815 945 18985 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 2495 7055 2665 7225 ;
    LAYER V1 ;
      RECT 2495 12935 2665 13105 ;
    LAYER V1 ;
      RECT 2495 18815 2665 18985 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 4215 7055 4385 7225 ;
    LAYER V1 ;
      RECT 4215 12935 4385 13105 ;
    LAYER V1 ;
      RECT 4215 18815 4385 18985 ;
    LAYER V1 ;
      RECT 5935 1175 6105 1345 ;
    LAYER V1 ;
      RECT 5935 7055 6105 7225 ;
    LAYER V1 ;
      RECT 5935 12935 6105 13105 ;
    LAYER V1 ;
      RECT 5935 18815 6105 18985 ;
    LAYER V1 ;
      RECT 7655 1175 7825 1345 ;
    LAYER V1 ;
      RECT 7655 7055 7825 7225 ;
    LAYER V1 ;
      RECT 7655 12935 7825 13105 ;
    LAYER V1 ;
      RECT 7655 18815 7825 18985 ;
    LAYER V2 ;
      RECT 3795 345 3945 495 ;
    LAYER V2 ;
      RECT 3795 4545 3945 4695 ;
    LAYER V2 ;
      RECT 3795 6225 3945 6375 ;
    LAYER V2 ;
      RECT 3795 10425 3945 10575 ;
    LAYER V2 ;
      RECT 3795 12105 3945 12255 ;
    LAYER V2 ;
      RECT 3795 16305 3945 16455 ;
    LAYER V2 ;
      RECT 3795 17985 3945 18135 ;
    LAYER V2 ;
      RECT 3795 22185 3945 22335 ;
    LAYER V2 ;
      RECT 4225 765 4375 915 ;
    LAYER V2 ;
      RECT 4225 6645 4375 6795 ;
    LAYER V2 ;
      RECT 4225 12525 4375 12675 ;
    LAYER V2 ;
      RECT 4225 18405 4375 18555 ;
    LAYER V2 ;
      RECT 4655 1185 4805 1335 ;
    LAYER V2 ;
      RECT 4655 7065 4805 7215 ;
    LAYER V2 ;
      RECT 4655 12945 4805 13095 ;
    LAYER V2 ;
      RECT 4655 18825 4805 18975 ;
  END
END SCM_NMOS_B_85279373_X2_Y4
