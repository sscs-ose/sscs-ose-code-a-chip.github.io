magic
tech sky130A
magscale 1 2
timestamp 1762074413
<< error_p >>
rect -29 60081 29 60087
rect -29 60047 -17 60081
rect -29 60041 29 60047
rect -29 -60047 29 -60041
rect -29 -60081 -17 -60047
rect -29 -60087 29 -60081
<< nwell >>
rect -211 -60219 211 60219
<< pmos >>
rect -15 -60000 15 60000
<< pdiff >>
rect -73 59988 -15 60000
rect -73 -59988 -61 59988
rect -27 -59988 -15 59988
rect -73 -60000 -15 -59988
rect 15 59988 73 60000
rect 15 -59988 27 59988
rect 61 -59988 73 59988
rect 15 -60000 73 -59988
<< pdiffc >>
rect -61 -59988 -27 59988
rect 27 -59988 61 59988
<< nsubdiff >>
rect -175 60149 -79 60183
rect 79 60149 175 60183
rect -175 60087 -141 60149
rect 141 60087 175 60149
rect -175 -60149 -141 -60087
rect 141 -60149 175 -60087
rect -175 -60183 -79 -60149
rect 79 -60183 175 -60149
<< nsubdiffcont >>
rect -79 60149 79 60183
rect -175 -60087 -141 60087
rect 141 -60087 175 60087
rect -79 -60183 79 -60149
<< poly >>
rect -33 60081 33 60097
rect -33 60047 -17 60081
rect 17 60047 33 60081
rect -33 60031 33 60047
rect -15 60000 15 60031
rect -15 -60031 15 -60000
rect -33 -60047 33 -60031
rect -33 -60081 -17 -60047
rect 17 -60081 33 -60047
rect -33 -60097 33 -60081
<< polycont >>
rect -17 60047 17 60081
rect -17 -60081 17 -60047
<< locali >>
rect -175 60149 -79 60183
rect 79 60149 175 60183
rect -175 60087 -141 60149
rect 141 60087 175 60149
rect -33 60047 -17 60081
rect 17 60047 33 60081
rect -61 59988 -27 60004
rect -61 -60004 -27 -59988
rect 27 59988 61 60004
rect 27 -60004 61 -59988
rect -33 -60081 -17 -60047
rect 17 -60081 33 -60047
rect -175 -60149 -141 -60087
rect 141 -60149 175 -60087
rect -175 -60183 -79 -60149
rect 79 -60183 175 -60149
<< viali >>
rect -17 60047 17 60081
rect -61 -59988 -27 59988
rect 27 -59988 61 59988
rect -17 -60081 17 -60047
<< metal1 >>
rect -29 60081 29 60087
rect -29 60047 -17 60081
rect 17 60047 29 60081
rect -29 60041 29 60047
rect -67 59988 -21 60000
rect -67 -59988 -61 59988
rect -27 -59988 -21 59988
rect -67 -60000 -21 -59988
rect 21 59988 67 60000
rect 21 -59988 27 59988
rect 61 -59988 67 59988
rect 21 -60000 67 -59988
rect -29 -60047 29 -60041
rect -29 -60081 -17 -60047
rect 17 -60081 29 -60047
rect -29 -60087 29 -60081
<< labels >>
rlabel nsubdiffcont 0 -60166 0 -60166 0 B
port 1 nsew
rlabel pdiffc -44 0 -44 0 0 D
port 2 nsew
rlabel pdiffc 44 0 44 0 0 S
port 3 nsew
rlabel polycont 0 60064 0 60064 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -60166 158 60166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 600 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
