* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 0
.param
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = 1.0050e+0
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = 1.0090e+0
.include "sky130_fd_pr__pfet_g5v0d10v5__tt.pm3.spice"
