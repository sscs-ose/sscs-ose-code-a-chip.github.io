# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__npn_11v0_W1p00L1p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__npn_11v0_W1p00L1p00 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.750000 BY  9.750000 ;
  PIN B
    ANTENNADIFFAREA  5.903200 ;
    ANTENNAGATEAREA  47.472099 ;
    PORT
      LAYER met1 ;
        RECT 1.680000 1.690000 8.060000 2.050000 ;
        RECT 1.680000 2.050000 2.040000 4.065000 ;
        RECT 1.680000 5.680000 2.040000 7.700000 ;
        RECT 1.680000 7.700000 8.060000 8.060000 ;
        RECT 7.700000 2.050000 8.060000 7.700000 ;
    END
  END B
  PIN C
    ANTENNADIFFAREA  13.07080 ;
    PORT
      LAYER met1 ;
        RECT 0.710000 0.710000 9.040000 1.070000 ;
        RECT 0.710000 1.070000 1.070000 8.685000 ;
        RECT 0.710000 8.685000 9.040000 9.045000 ;
        RECT 8.680000 1.070000 9.040000 8.685000 ;
    END
  END C
  PIN E
    ANTENNADIFFAREA  2.068700 ;
    ANTENNAGATEAREA  19.808849 ;
    PORT
      LAYER met1 ;
        RECT 1.445000 4.310000 2.395000 5.440000 ;
    END
  END E
  OBS
    LAYER li1 ;
      RECT 0.685000 0.685000 9.065000 1.095000 ;
      RECT 0.685000 1.095000 1.095000 8.655000 ;
      RECT 0.685000 8.655000 9.065000 9.065000 ;
      RECT 1.305000 4.370000 5.380000 5.380000 ;
      RECT 1.660000 1.670000 8.080000 2.070000 ;
      RECT 1.660000 2.070000 2.070000 4.065000 ;
      RECT 1.660000 5.680000 2.070000 7.680000 ;
      RECT 1.660000 7.680000 8.080000 8.080000 ;
      RECT 7.680000 2.070000 8.080000 7.680000 ;
      RECT 8.655000 1.095000 9.065000 8.655000 ;
    LAYER mcon ;
      RECT 0.805000 1.295000 0.975000 1.465000 ;
      RECT 0.805000 1.660000 0.975000 1.830000 ;
      RECT 0.805000 2.025000 0.975000 2.195000 ;
      RECT 0.805000 2.390000 0.975000 2.560000 ;
      RECT 0.805000 2.760000 0.975000 2.930000 ;
      RECT 0.805000 3.130000 0.975000 3.300000 ;
      RECT 0.805000 3.500000 0.975000 3.670000 ;
      RECT 0.805000 3.870000 0.975000 4.040000 ;
      RECT 0.805000 4.240000 0.975000 4.410000 ;
      RECT 0.805000 4.610000 0.975000 4.780000 ;
      RECT 0.805000 4.980000 0.975000 5.150000 ;
      RECT 0.805000 5.350000 0.975000 5.520000 ;
      RECT 0.805000 5.720000 0.975000 5.890000 ;
      RECT 0.805000 6.090000 0.975000 6.260000 ;
      RECT 0.805000 6.460000 0.975000 6.630000 ;
      RECT 0.805000 6.830000 0.975000 7.000000 ;
      RECT 0.805000 7.200000 0.975000 7.370000 ;
      RECT 0.805000 7.570000 0.975000 7.740000 ;
      RECT 0.805000 7.940000 0.975000 8.110000 ;
      RECT 0.805000 8.310000 0.975000 8.480000 ;
      RECT 1.295000 0.805000 1.465000 0.975000 ;
      RECT 1.295000 8.775000 1.465000 8.945000 ;
      RECT 1.475000 4.370000 1.645000 4.540000 ;
      RECT 1.475000 4.790000 1.645000 4.960000 ;
      RECT 1.475000 5.210000 1.645000 5.380000 ;
      RECT 1.660000 0.805000 1.830000 0.975000 ;
      RECT 1.660000 8.775000 1.830000 8.945000 ;
      RECT 1.775000 2.080000 1.945000 2.250000 ;
      RECT 1.775000 2.520000 1.945000 2.690000 ;
      RECT 1.775000 2.960000 1.945000 3.130000 ;
      RECT 1.775000 3.400000 1.945000 3.570000 ;
      RECT 1.775000 3.835000 1.945000 4.005000 ;
      RECT 1.775000 5.740000 1.945000 5.910000 ;
      RECT 1.775000 6.165000 1.945000 6.335000 ;
      RECT 1.775000 6.590000 1.945000 6.760000 ;
      RECT 1.775000 7.015000 1.945000 7.185000 ;
      RECT 1.775000 7.440000 1.945000 7.610000 ;
      RECT 1.835000 4.370000 2.005000 4.540000 ;
      RECT 1.835000 4.790000 2.005000 4.960000 ;
      RECT 1.835000 5.210000 2.005000 5.380000 ;
      RECT 2.025000 0.805000 2.195000 0.975000 ;
      RECT 2.025000 8.775000 2.195000 8.945000 ;
      RECT 2.070000 7.795000 2.240000 7.965000 ;
      RECT 2.195000 4.370000 2.365000 4.540000 ;
      RECT 2.195000 4.790000 2.365000 4.960000 ;
      RECT 2.195000 5.210000 2.365000 5.380000 ;
      RECT 2.390000 0.805000 2.560000 0.975000 ;
      RECT 2.390000 8.775000 2.560000 8.945000 ;
      RECT 2.430000 1.785000 2.600000 1.955000 ;
      RECT 2.435000 7.795000 2.605000 7.965000 ;
      RECT 2.755000 0.805000 2.925000 0.975000 ;
      RECT 2.755000 8.775000 2.925000 8.945000 ;
      RECT 2.790000 1.785000 2.960000 1.955000 ;
      RECT 2.800000 7.795000 2.970000 7.965000 ;
      RECT 3.125000 0.805000 3.295000 0.975000 ;
      RECT 3.125000 8.775000 3.295000 8.945000 ;
      RECT 3.150000 1.785000 3.320000 1.955000 ;
      RECT 3.165000 7.795000 3.335000 7.965000 ;
      RECT 3.495000 0.805000 3.665000 0.975000 ;
      RECT 3.495000 8.775000 3.665000 8.945000 ;
      RECT 3.510000 1.785000 3.680000 1.955000 ;
      RECT 3.530000 7.795000 3.700000 7.965000 ;
      RECT 3.865000 0.805000 4.035000 0.975000 ;
      RECT 3.865000 8.775000 4.035000 8.945000 ;
      RECT 3.870000 1.785000 4.040000 1.955000 ;
      RECT 3.895000 7.795000 4.065000 7.965000 ;
      RECT 4.230000 1.785000 4.400000 1.955000 ;
      RECT 4.235000 0.805000 4.405000 0.975000 ;
      RECT 4.235000 8.775000 4.405000 8.945000 ;
      RECT 4.260000 7.795000 4.430000 7.965000 ;
      RECT 4.590000 1.785000 4.760000 1.955000 ;
      RECT 4.605000 0.805000 4.775000 0.975000 ;
      RECT 4.605000 8.775000 4.775000 8.945000 ;
      RECT 4.620000 7.795000 4.790000 7.965000 ;
      RECT 4.950000 1.785000 5.120000 1.955000 ;
      RECT 4.975000 0.805000 5.145000 0.975000 ;
      RECT 4.975000 8.775000 5.145000 8.945000 ;
      RECT 4.980000 7.795000 5.150000 7.965000 ;
      RECT 5.310000 1.785000 5.480000 1.955000 ;
      RECT 5.340000 7.795000 5.510000 7.965000 ;
      RECT 5.345000 0.805000 5.515000 0.975000 ;
      RECT 5.345000 8.775000 5.515000 8.945000 ;
      RECT 5.675000 1.785000 5.845000 1.955000 ;
      RECT 5.700000 7.795000 5.870000 7.965000 ;
      RECT 5.715000 0.805000 5.885000 0.975000 ;
      RECT 5.715000 8.775000 5.885000 8.945000 ;
      RECT 6.040000 1.785000 6.210000 1.955000 ;
      RECT 6.060000 7.795000 6.230000 7.965000 ;
      RECT 6.085000 0.805000 6.255000 0.975000 ;
      RECT 6.085000 8.775000 6.255000 8.945000 ;
      RECT 6.405000 1.785000 6.575000 1.955000 ;
      RECT 6.420000 7.795000 6.590000 7.965000 ;
      RECT 6.455000 0.805000 6.625000 0.975000 ;
      RECT 6.455000 8.775000 6.625000 8.945000 ;
      RECT 6.770000 1.785000 6.940000 1.955000 ;
      RECT 6.780000 7.795000 6.950000 7.965000 ;
      RECT 6.825000 0.805000 6.995000 0.975000 ;
      RECT 6.825000 8.775000 6.995000 8.945000 ;
      RECT 7.135000 1.785000 7.305000 1.955000 ;
      RECT 7.140000 7.795000 7.310000 7.965000 ;
      RECT 7.195000 0.805000 7.365000 0.975000 ;
      RECT 7.195000 8.775000 7.365000 8.945000 ;
      RECT 7.500000 1.785000 7.670000 1.955000 ;
      RECT 7.565000 0.805000 7.735000 0.975000 ;
      RECT 7.565000 8.775000 7.735000 8.945000 ;
      RECT 7.795000 2.440000 7.965000 2.610000 ;
      RECT 7.795000 2.800000 7.965000 2.970000 ;
      RECT 7.795000 3.160000 7.965000 3.330000 ;
      RECT 7.795000 3.520000 7.965000 3.690000 ;
      RECT 7.795000 3.880000 7.965000 4.050000 ;
      RECT 7.795000 4.240000 7.965000 4.410000 ;
      RECT 7.795000 4.600000 7.965000 4.770000 ;
      RECT 7.795000 4.960000 7.965000 5.130000 ;
      RECT 7.795000 5.320000 7.965000 5.490000 ;
      RECT 7.795000 5.680000 7.965000 5.850000 ;
      RECT 7.795000 6.040000 7.965000 6.210000 ;
      RECT 7.795000 6.405000 7.965000 6.575000 ;
      RECT 7.795000 6.770000 7.965000 6.940000 ;
      RECT 7.795000 7.135000 7.965000 7.305000 ;
      RECT 7.795000 7.500000 7.965000 7.670000 ;
      RECT 7.935000 0.805000 8.105000 0.975000 ;
      RECT 7.935000 8.775000 8.105000 8.945000 ;
      RECT 8.305000 0.805000 8.475000 0.975000 ;
      RECT 8.305000 8.775000 8.475000 8.945000 ;
      RECT 8.775000 1.295000 8.945000 1.465000 ;
      RECT 8.775000 1.660000 8.945000 1.830000 ;
      RECT 8.775000 2.025000 8.945000 2.195000 ;
      RECT 8.775000 2.390000 8.945000 2.560000 ;
      RECT 8.775000 2.760000 8.945000 2.930000 ;
      RECT 8.775000 3.130000 8.945000 3.300000 ;
      RECT 8.775000 3.500000 8.945000 3.670000 ;
      RECT 8.775000 3.870000 8.945000 4.040000 ;
      RECT 8.775000 4.240000 8.945000 4.410000 ;
      RECT 8.775000 4.610000 8.945000 4.780000 ;
      RECT 8.775000 4.980000 8.945000 5.150000 ;
      RECT 8.775000 5.350000 8.945000 5.520000 ;
      RECT 8.775000 5.720000 8.945000 5.890000 ;
      RECT 8.775000 6.090000 8.945000 6.260000 ;
      RECT 8.775000 6.460000 8.945000 6.630000 ;
      RECT 8.775000 6.830000 8.945000 7.000000 ;
      RECT 8.775000 7.200000 8.945000 7.370000 ;
      RECT 8.775000 7.570000 8.945000 7.740000 ;
      RECT 8.775000 7.940000 8.945000 8.110000 ;
      RECT 8.775000 8.310000 8.945000 8.480000 ;
  END
END sky130_fd_pr__npn_11v0_W1p00L1p00
END LIBRARY
