magic
tech sky130A
magscale 1 2
timestamp 1762074413
<< error_p >>
rect -29 24072 29 24078
rect -29 24038 -17 24072
rect -29 24032 29 24038
rect -29 -24038 29 -24032
rect -29 -24072 -17 -24038
rect -29 -24078 29 -24072
<< pwell >>
rect -211 -24210 211 24210
<< nmos >>
rect -15 -24000 15 24000
<< ndiff >>
rect -73 23988 -15 24000
rect -73 -23988 -61 23988
rect -27 -23988 -15 23988
rect -73 -24000 -15 -23988
rect 15 23988 73 24000
rect 15 -23988 27 23988
rect 61 -23988 73 23988
rect 15 -24000 73 -23988
<< ndiffc >>
rect -61 -23988 -27 23988
rect 27 -23988 61 23988
<< psubdiff >>
rect -175 24140 -79 24174
rect 79 24140 175 24174
rect -175 24078 -141 24140
rect 141 24078 175 24140
rect -175 -24140 -141 -24078
rect 141 -24140 175 -24078
rect -175 -24174 -79 -24140
rect 79 -24174 175 -24140
<< psubdiffcont >>
rect -79 24140 79 24174
rect -175 -24078 -141 24078
rect 141 -24078 175 24078
rect -79 -24174 79 -24140
<< poly >>
rect -33 24072 33 24088
rect -33 24038 -17 24072
rect 17 24038 33 24072
rect -33 24022 33 24038
rect -15 24000 15 24022
rect -15 -24022 15 -24000
rect -33 -24038 33 -24022
rect -33 -24072 -17 -24038
rect 17 -24072 33 -24038
rect -33 -24088 33 -24072
<< polycont >>
rect -17 24038 17 24072
rect -17 -24072 17 -24038
<< locali >>
rect -175 24140 -79 24174
rect 79 24140 175 24174
rect -175 24078 -141 24140
rect 141 24078 175 24140
rect -33 24038 -17 24072
rect 17 24038 33 24072
rect -61 23988 -27 24004
rect -61 -24004 -27 -23988
rect 27 23988 61 24004
rect 27 -24004 61 -23988
rect -33 -24072 -17 -24038
rect 17 -24072 33 -24038
rect -175 -24140 -141 -24078
rect 141 -24140 175 -24078
rect -175 -24174 -79 -24140
rect 79 -24174 175 -24140
<< viali >>
rect -17 24038 17 24072
rect -61 -23988 -27 23988
rect 27 -23988 61 23988
rect -17 -24072 17 -24038
<< metal1 >>
rect -29 24072 29 24078
rect -29 24038 -17 24072
rect 17 24038 29 24072
rect -29 24032 29 24038
rect -67 23988 -21 24000
rect -67 -23988 -61 23988
rect -27 -23988 -21 23988
rect -67 -24000 -21 -23988
rect 21 23988 67 24000
rect 21 -23988 27 23988
rect 61 -23988 67 23988
rect 21 -24000 67 -23988
rect -29 -24038 29 -24032
rect -29 -24072 -17 -24038
rect 17 -24072 29 -24038
rect -29 -24078 29 -24072
<< labels >>
rlabel psubdiffcont 0 -24157 0 -24157 0 B
port 1 nsew
rlabel ndiffc -44 0 -44 0 0 D
port 2 nsew
rlabel ndiffc 44 0 44 0 0 S
port 3 nsew
rlabel polycont 0 24055 0 24055 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -24157 158 24157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 240 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
