# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25 ;
  ORIGIN -0.050000 -0.050000 ;
  SIZE  3.780000 BY  2.570000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 1.460000 3.830000 2.100000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.650000 ;
    PORT
      LAYER li1 ;
        RECT 0.925000 0.150000 2.955000 0.320000 ;
        RECT 0.925000 2.350000 2.955000 2.520000 ;
      LAYER mcon ;
        RECT 0.960000 0.150000 1.130000 0.320000 ;
        RECT 0.960000 2.350000 1.130000 2.520000 ;
        RECT 1.320000 0.150000 1.490000 0.320000 ;
        RECT 1.320000 2.350000 1.490000 2.520000 ;
        RECT 1.680000 0.150000 1.850000 0.320000 ;
        RECT 1.680000 2.350000 1.850000 2.520000 ;
        RECT 2.040000 0.150000 2.210000 0.320000 ;
        RECT 2.040000 2.350000 2.210000 2.520000 ;
        RECT 2.400000 0.150000 2.570000 0.320000 ;
        RECT 2.400000 2.350000 2.570000 2.520000 ;
        RECT 2.760000 0.150000 2.930000 0.320000 ;
        RECT 2.760000 2.350000 2.930000 2.520000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.900000 0.050000 2.990000 0.380000 ;
        RECT 0.900000 2.290000 2.990000 2.620000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.570000 3.830000 1.210000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.478500 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.570000 0.470000 2.100000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.410000 0.570000 3.700000 2.100000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.660000 0.410000 2.010000 ;
      RECT 0.795000 0.490000 0.965000 2.180000 ;
      RECT 1.325000 0.490000 1.495000 2.180000 ;
      RECT 1.855000 0.490000 2.025000 2.180000 ;
      RECT 2.385000 0.490000 2.555000 2.180000 ;
      RECT 2.915000 0.490000 3.085000 2.180000 ;
      RECT 3.470000 0.660000 3.640000 2.010000 ;
    LAYER mcon ;
      RECT 0.240000 0.710000 0.410000 0.880000 ;
      RECT 0.240000 1.070000 0.410000 1.240000 ;
      RECT 0.240000 1.430000 0.410000 1.600000 ;
      RECT 0.240000 1.790000 0.410000 1.960000 ;
      RECT 0.795000 0.710000 0.965000 0.880000 ;
      RECT 0.795000 1.070000 0.965000 1.240000 ;
      RECT 0.795000 1.430000 0.965000 1.600000 ;
      RECT 0.795000 1.790000 0.965000 1.960000 ;
      RECT 1.325000 0.710000 1.495000 0.880000 ;
      RECT 1.325000 1.070000 1.495000 1.240000 ;
      RECT 1.325000 1.430000 1.495000 1.600000 ;
      RECT 1.325000 1.790000 1.495000 1.960000 ;
      RECT 1.855000 0.710000 2.025000 0.880000 ;
      RECT 1.855000 1.070000 2.025000 1.240000 ;
      RECT 1.855000 1.430000 2.025000 1.600000 ;
      RECT 1.855000 1.790000 2.025000 1.960000 ;
      RECT 2.385000 0.710000 2.555000 0.880000 ;
      RECT 2.385000 1.070000 2.555000 1.240000 ;
      RECT 2.385000 1.430000 2.555000 1.600000 ;
      RECT 2.385000 1.790000 2.555000 1.960000 ;
      RECT 2.915000 0.710000 3.085000 0.880000 ;
      RECT 2.915000 1.070000 3.085000 1.240000 ;
      RECT 2.915000 1.430000 3.085000 1.600000 ;
      RECT 2.915000 1.790000 3.085000 1.960000 ;
      RECT 3.470000 0.710000 3.640000 0.880000 ;
      RECT 3.470000 1.070000 3.640000 1.240000 ;
      RECT 3.470000 1.430000 3.640000 1.600000 ;
      RECT 3.470000 1.790000 3.640000 1.960000 ;
    LAYER met1 ;
      RECT 0.750000 0.570000 1.010000 2.100000 ;
      RECT 1.280000 0.570000 1.540000 2.100000 ;
      RECT 1.810000 0.570000 2.070000 2.100000 ;
      RECT 2.340000 0.570000 2.600000 2.100000 ;
      RECT 2.870000 0.570000 3.130000 2.100000 ;
    LAYER via ;
      RECT 0.750000 0.600000 1.010000 0.860000 ;
      RECT 0.750000 0.920000 1.010000 1.180000 ;
      RECT 1.280000 1.490000 1.540000 1.750000 ;
      RECT 1.280000 1.810000 1.540000 2.070000 ;
      RECT 1.810000 0.600000 2.070000 0.860000 ;
      RECT 1.810000 0.920000 2.070000 1.180000 ;
      RECT 2.340000 1.490000 2.600000 1.750000 ;
      RECT 2.340000 1.810000 2.600000 2.070000 ;
      RECT 2.870000 0.600000 3.130000 0.860000 ;
      RECT 2.870000 0.920000 3.130000 1.180000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25
END LIBRARY
