* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+ sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult = 0.958
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult = 1.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult = 0.7713
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult = 9.5405e-1
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult = 9.6374e-1
+ sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff = 1.21275e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff = -2.252e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff = 1.21275e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff = -2.252e-8
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0 = -0.001863
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0 = 0.001058
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0 = -31427.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0 = 0.041954
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0 = -0.08688
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0 = 4.3035e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0 = -3.1175e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0 = 0.021424
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1 = 0.013438
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1 = -0.0020179
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1 = 0.0010444
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1 = -28354.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1 = 0.048874
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1 = -1.42e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1 = -0.065937
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1 = -2.3727e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2 = 0.017194
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2 = -0.0016532
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2 = 0.00075934
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2 = 0.051024
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2 = -7.6179e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2 = -27569.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2 = -0.094908
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2 = -2.0807e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3 = 0.018257
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3 = -0.0025581
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3 = 0.00124927
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3 = 0.044703
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3 = 7.5609e-12
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3 = -35289.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3 = -0.086391
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3 = -3.2769e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4 = 0.025977
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4 = -0.0013669
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4 = 0.00091382
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4 = 0.043787
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4 = 1.574e-10
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4 = -24808.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4 = 0.078325
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4 = -4.9963e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5 = 0.020181
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5 = -0.0021503
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5 = 0.0010663
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5 = 0.043391
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5 = -1.0798e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5 = -22995.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5 = -0.11963
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5 = -1.3111e-19
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6 = -1.868e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6 = 0.019337
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6 = -0.0018306
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6 = 0.00086193
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6 = 0.045188
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6 = -1.1042e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6 = -24982.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6 = -0.11297
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7 = -2.3793e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7 = 0.022032
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7 = -0.0019486
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7 = 0.00096865
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7 = 0.045761
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7 = -2.12e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7 = -21171.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7 = -0.13265
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7 = 0.0
.include "sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"
