magic
tech sky130A
magscale 1 2
timestamp 1762087944
<< error_p >>
rect -29 60045 29 60051
rect -29 60011 -17 60045
rect -29 60005 29 60011
<< nwell >>
rect -211 -60184 211 60184
<< pmos >>
rect -15 -60036 15 59964
<< pdiff >>
rect -73 59952 -15 59964
rect -73 -60024 -61 59952
rect -27 -60024 -15 59952
rect -73 -60036 -15 -60024
rect 15 59952 73 59964
rect 15 -60024 27 59952
rect 61 -60024 73 59952
rect 15 -60036 73 -60024
<< pdiffc >>
rect -61 -60024 -27 59952
rect 27 -60024 61 59952
<< nsubdiff >>
rect -175 60114 -79 60148
rect 79 60114 175 60148
rect -175 60051 -141 60114
rect 141 60051 175 60114
rect -175 -60114 -141 -60051
rect 141 -60114 175 -60051
rect -175 -60148 -79 -60114
rect 79 -60148 175 -60114
<< nsubdiffcont >>
rect -79 60114 79 60148
rect -175 -60051 -141 60051
rect 141 -60051 175 60051
rect -79 -60148 79 -60114
<< poly >>
rect -33 60045 33 60061
rect -33 60011 -17 60045
rect 17 60011 33 60045
rect -33 59995 33 60011
rect -15 59964 15 59995
rect -15 -60062 15 -60036
<< polycont >>
rect -17 60011 17 60045
<< locali >>
rect -175 60114 -79 60148
rect 79 60114 175 60148
rect -175 60051 -141 60114
rect 141 60051 175 60114
rect -33 60011 -17 60045
rect 17 60011 33 60045
rect -61 59952 -27 59968
rect -61 -60040 -27 -60024
rect 27 59952 61 59968
rect 27 -60040 61 -60024
rect -175 -60114 -141 -60051
rect 141 -60114 175 -60051
rect -175 -60148 -79 -60114
rect 79 -60148 175 -60114
<< viali >>
rect -17 60011 17 60045
rect -61 -60024 -27 59952
rect 27 -60024 61 59952
<< metal1 >>
rect -29 60045 29 60051
rect -29 60011 -17 60045
rect 17 60011 29 60045
rect -29 60005 29 60011
rect -67 59952 -21 59964
rect -67 -60024 -61 59952
rect -27 -60024 -21 59952
rect -67 -60036 -21 -60024
rect 21 59952 67 59964
rect 21 -60024 27 59952
rect 61 -60024 67 59952
rect 21 -60036 67 -60024
<< labels >>
rlabel nsubdiffcont 0 -60131 0 -60131 0 B
port 1 nsew
rlabel pdiffc -44 -36 -44 -36 0 D
port 2 nsew
rlabel pdiffc 44 -36 44 -36 0 S
port 3 nsew
rlabel polycont 0 60028 0 60028 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -60131 158 60131
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 600 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
