** sch_path: /home/evadeltor/VMA.sch
**.subckt VMA VIN+ VIN- VOUT IBIAS
*.ipin VIN+
*.ipin VIN-
*.opin VOUT
*.opin IBIAS
X2 net13 net12 VDD irf5305
X4 VOUT net11 net13 irf5305
X6 net12 net12 VDD irf5305
X8 net11 net11 net12 irf5305
X9 net8 VIN+ IBIAS irf5305
X10 net9 VIN- IBIAS irf5305
X11 VOUT net8 net7 irf540 m=1
X12 net9 net9 net2 irf540 m=1
X13 net8 net8 net4 irf540 m=1
X14 net11 net9 net10 irf540 m=1
X15 net10 net2 net1 irf540 m=1
X16 net1 net2 GND irf540 m=1
X17 net2 net2 net6 irf540 m=1
X18 net6 net2 GND irf540 m=1
X19 net6 net4 GND irf540 m=1
X20 net5 net2 GND irf540 m=1
X21 net5 net4 GND irf540 m=1
X22 net4 net4 net5 irf540 m=1
X23 net3 net4 GND irf540 m=1
X24 net7 net4 net3 irf540 m=1
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
