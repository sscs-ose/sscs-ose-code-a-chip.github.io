# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  1.140000 BY  4.110000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.840000 ;
    PORT
      LAYER met2 ;
        RECT 0.620000 2.440000 0.880000 3.080000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.900000 ;
    PORT
      LAYER met1 ;
        RECT 0.425000 3.355000 1.075000 3.645000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.680000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 1.295000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  3.105000 ;
        RECT 1.065000 -0.145000 1.295000  3.105000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.400000 3.200000 0.450000 3.285000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.235000 0.405000 3.105000 ;
      RECT 0.415000 3.335000 1.085000 3.665000 ;
      RECT 0.665000 0.255000 0.835000 3.105000 ;
      RECT 1.095000 0.255000 1.265000 3.105000 ;
    LAYER mcon ;
      RECT 0.235000 0.335000 0.405000 0.505000 ;
      RECT 0.235000 0.695000 0.405000 0.865000 ;
      RECT 0.235000 1.055000 0.405000 1.225000 ;
      RECT 0.235000 1.415000 0.405000 1.585000 ;
      RECT 0.235000 1.775000 0.405000 1.945000 ;
      RECT 0.235000 2.135000 0.405000 2.305000 ;
      RECT 0.235000 2.495000 0.405000 2.665000 ;
      RECT 0.235000 2.855000 0.405000 3.025000 ;
      RECT 0.485000 3.415000 0.655000 3.585000 ;
      RECT 0.665000 0.335000 0.835000 0.505000 ;
      RECT 0.665000 0.695000 0.835000 0.865000 ;
      RECT 0.665000 1.055000 0.835000 1.225000 ;
      RECT 0.665000 1.415000 0.835000 1.585000 ;
      RECT 0.665000 1.775000 0.835000 1.945000 ;
      RECT 0.665000 2.135000 0.835000 2.305000 ;
      RECT 0.665000 2.495000 0.835000 2.665000 ;
      RECT 0.665000 2.855000 0.835000 3.025000 ;
      RECT 0.845000 3.415000 1.015000 3.585000 ;
      RECT 1.095000 0.335000 1.265000 0.505000 ;
      RECT 1.095000 0.695000 1.265000 0.865000 ;
      RECT 1.095000 1.055000 1.265000 1.225000 ;
      RECT 1.095000 1.415000 1.265000 1.585000 ;
      RECT 1.095000 1.775000 1.265000 1.945000 ;
      RECT 1.095000 2.135000 1.265000 2.305000 ;
      RECT 1.095000 2.495000 1.265000 2.665000 ;
      RECT 1.095000 2.855000 1.265000 3.025000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 3.105000 ;
    LAYER via ;
      RECT 0.620000 2.470000 0.880000 2.730000 ;
      RECT 0.620000 2.790000 0.880000 3.050000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15
END LIBRARY
