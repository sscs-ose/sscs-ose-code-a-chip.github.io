# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_npn_05v5_W1p00L8p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_npn_05v5_W1p00L8p00 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  9.700000 BY  16.70000 ;
  OBS
    LAYER li1 ;
      RECT 0.170000  0.170000 9.790000  0.500000 ;
      RECT 0.170000  0.500000 0.500000 16.460000 ;
      RECT 0.170000 16.460000 9.790000 16.790000 ;
      RECT 1.300000  1.300000 8.660000  1.630000 ;
      RECT 1.300000  1.630000 1.630000 15.330000 ;
      RECT 1.300000 15.330000 8.660000 15.660000 ;
      RECT 3.310000  3.310000 6.650000  3.640000 ;
      RECT 3.310000  3.640000 3.640000 13.320000 ;
      RECT 3.310000 13.320000 6.650000 13.650000 ;
      RECT 4.475000  4.475000 5.485000 12.485000 ;
      RECT 6.320000  3.640000 6.650000 13.320000 ;
      RECT 8.330000  1.630000 8.660000 15.330000 ;
      RECT 9.460000  0.500000 9.790000 16.460000 ;
    LAYER mcon ;
      RECT 0.250000  0.250000 0.420000  0.420000 ;
      RECT 0.250000  0.655000 0.420000  0.825000 ;
      RECT 0.250000  1.015000 0.420000  1.185000 ;
      RECT 0.250000  1.375000 0.420000  1.545000 ;
      RECT 0.250000  1.735000 0.420000  1.905000 ;
      RECT 0.250000  2.095000 0.420000  2.265000 ;
      RECT 0.250000  2.455000 0.420000  2.625000 ;
      RECT 0.250000  2.815000 0.420000  2.985000 ;
      RECT 0.250000  3.175000 0.420000  3.345000 ;
      RECT 0.250000  3.535000 0.420000  3.705000 ;
      RECT 0.250000  3.895000 0.420000  4.065000 ;
      RECT 0.250000  4.255000 0.420000  4.425000 ;
      RECT 0.250000  4.615000 0.420000  4.785000 ;
      RECT 0.250000  4.975000 0.420000  5.145000 ;
      RECT 0.250000  5.335000 0.420000  5.505000 ;
      RECT 0.250000  5.695000 0.420000  5.865000 ;
      RECT 0.250000  6.055000 0.420000  6.225000 ;
      RECT 0.250000  6.415000 0.420000  6.585000 ;
      RECT 0.250000  6.775000 0.420000  6.945000 ;
      RECT 0.250000  7.135000 0.420000  7.305000 ;
      RECT 0.250000  7.495000 0.420000  7.665000 ;
      RECT 0.250000  7.855000 0.420000  8.025000 ;
      RECT 0.250000  8.215000 0.420000  8.385000 ;
      RECT 0.250000  8.575000 0.420000  8.745000 ;
      RECT 0.250000  8.935000 0.420000  9.105000 ;
      RECT 0.250000  9.295000 0.420000  9.465000 ;
      RECT 0.250000  9.655000 0.420000  9.825000 ;
      RECT 0.250000 10.015000 0.420000 10.185000 ;
      RECT 0.250000 10.375000 0.420000 10.545000 ;
      RECT 0.250000 10.735000 0.420000 10.905000 ;
      RECT 0.250000 11.095000 0.420000 11.265000 ;
      RECT 0.250000 11.455000 0.420000 11.625000 ;
      RECT 0.250000 11.815000 0.420000 11.985000 ;
      RECT 0.250000 12.175000 0.420000 12.345000 ;
      RECT 0.250000 12.535000 0.420000 12.705000 ;
      RECT 0.250000 12.895000 0.420000 13.065000 ;
      RECT 0.250000 13.255000 0.420000 13.425000 ;
      RECT 0.250000 13.615000 0.420000 13.785000 ;
      RECT 0.250000 13.975000 0.420000 14.145000 ;
      RECT 0.250000 14.335000 0.420000 14.505000 ;
      RECT 0.250000 14.695000 0.420000 14.865000 ;
      RECT 0.250000 15.055000 0.420000 15.225000 ;
      RECT 0.250000 15.415000 0.420000 15.585000 ;
      RECT 0.250000 15.775000 0.420000 15.945000 ;
      RECT 0.250000 16.135000 0.420000 16.305000 ;
      RECT 0.250000 16.540000 0.420000 16.710000 ;
      RECT 0.755000  0.250000 0.925000  0.420000 ;
      RECT 0.755000 16.540000 0.925000 16.710000 ;
      RECT 1.115000  0.250000 1.285000  0.420000 ;
      RECT 1.115000 16.540000 1.285000 16.710000 ;
      RECT 1.380000  1.380000 1.550000  1.550000 ;
      RECT 1.380000  1.915000 1.550000  2.085000 ;
      RECT 1.380000  2.275000 1.550000  2.445000 ;
      RECT 1.380000  2.635000 1.550000  2.805000 ;
      RECT 1.380000  2.995000 1.550000  3.165000 ;
      RECT 1.380000  3.355000 1.550000  3.525000 ;
      RECT 1.380000  3.715000 1.550000  3.885000 ;
      RECT 1.380000  4.075000 1.550000  4.245000 ;
      RECT 1.380000  4.435000 1.550000  4.605000 ;
      RECT 1.380000  4.795000 1.550000  4.965000 ;
      RECT 1.380000  5.155000 1.550000  5.325000 ;
      RECT 1.380000  5.515000 1.550000  5.685000 ;
      RECT 1.380000  5.875000 1.550000  6.045000 ;
      RECT 1.380000  6.235000 1.550000  6.405000 ;
      RECT 1.380000  6.595000 1.550000  6.765000 ;
      RECT 1.380000  6.955000 1.550000  7.125000 ;
      RECT 1.380000  7.315000 1.550000  7.485000 ;
      RECT 1.380000  7.675000 1.550000  7.845000 ;
      RECT 1.380000  8.035000 1.550000  8.205000 ;
      RECT 1.380000  8.395000 1.550000  8.565000 ;
      RECT 1.380000  8.755000 1.550000  8.925000 ;
      RECT 1.380000  9.115000 1.550000  9.285000 ;
      RECT 1.380000  9.475000 1.550000  9.645000 ;
      RECT 1.380000  9.835000 1.550000 10.005000 ;
      RECT 1.380000 10.195000 1.550000 10.365000 ;
      RECT 1.380000 10.555000 1.550000 10.725000 ;
      RECT 1.380000 10.915000 1.550000 11.085000 ;
      RECT 1.380000 11.275000 1.550000 11.445000 ;
      RECT 1.380000 11.635000 1.550000 11.805000 ;
      RECT 1.380000 11.995000 1.550000 12.165000 ;
      RECT 1.380000 12.355000 1.550000 12.525000 ;
      RECT 1.380000 12.715000 1.550000 12.885000 ;
      RECT 1.380000 13.075000 1.550000 13.245000 ;
      RECT 1.380000 13.435000 1.550000 13.605000 ;
      RECT 1.380000 13.795000 1.550000 13.965000 ;
      RECT 1.380000 14.155000 1.550000 14.325000 ;
      RECT 1.380000 14.515000 1.550000 14.685000 ;
      RECT 1.380000 14.875000 1.550000 15.045000 ;
      RECT 1.380000 15.410000 1.550000 15.580000 ;
      RECT 1.475000  0.250000 1.645000  0.420000 ;
      RECT 1.475000 16.540000 1.645000 16.710000 ;
      RECT 1.835000  0.250000 2.005000  0.420000 ;
      RECT 1.835000  1.380000 2.005000  1.550000 ;
      RECT 1.835000 15.410000 2.005000 15.580000 ;
      RECT 1.835000 16.540000 2.005000 16.710000 ;
      RECT 2.195000  0.250000 2.365000  0.420000 ;
      RECT 2.195000  1.380000 2.365000  1.550000 ;
      RECT 2.195000 15.410000 2.365000 15.580000 ;
      RECT 2.195000 16.540000 2.365000 16.710000 ;
      RECT 2.555000  0.250000 2.725000  0.420000 ;
      RECT 2.555000  1.380000 2.725000  1.550000 ;
      RECT 2.555000 15.410000 2.725000 15.580000 ;
      RECT 2.555000 16.540000 2.725000 16.710000 ;
      RECT 2.915000  0.250000 3.085000  0.420000 ;
      RECT 2.915000  1.380000 3.085000  1.550000 ;
      RECT 2.915000 15.410000 3.085000 15.580000 ;
      RECT 2.915000 16.540000 3.085000 16.710000 ;
      RECT 3.275000  0.250000 3.445000  0.420000 ;
      RECT 3.275000  1.380000 3.445000  1.550000 ;
      RECT 3.275000 15.410000 3.445000 15.580000 ;
      RECT 3.275000 16.540000 3.445000 16.710000 ;
      RECT 3.390000  3.390000 3.560000  3.560000 ;
      RECT 3.390000  3.895000 3.560000  4.065000 ;
      RECT 3.390000  4.255000 3.560000  4.425000 ;
      RECT 3.390000  4.615000 3.560000  4.785000 ;
      RECT 3.390000  4.975000 3.560000  5.145000 ;
      RECT 3.390000  5.335000 3.560000  5.505000 ;
      RECT 3.390000  5.695000 3.560000  5.865000 ;
      RECT 3.390000  6.055000 3.560000  6.225000 ;
      RECT 3.390000  6.415000 3.560000  6.585000 ;
      RECT 3.390000  6.775000 3.560000  6.945000 ;
      RECT 3.390000  7.135000 3.560000  7.305000 ;
      RECT 3.390000  7.495000 3.560000  7.665000 ;
      RECT 3.390000  7.855000 3.560000  8.025000 ;
      RECT 3.390000  8.215000 3.560000  8.385000 ;
      RECT 3.390000  8.575000 3.560000  8.745000 ;
      RECT 3.390000  8.935000 3.560000  9.105000 ;
      RECT 3.390000  9.295000 3.560000  9.465000 ;
      RECT 3.390000  9.655000 3.560000  9.825000 ;
      RECT 3.390000 10.015000 3.560000 10.185000 ;
      RECT 3.390000 10.375000 3.560000 10.545000 ;
      RECT 3.390000 10.735000 3.560000 10.905000 ;
      RECT 3.390000 11.095000 3.560000 11.265000 ;
      RECT 3.390000 11.455000 3.560000 11.625000 ;
      RECT 3.390000 11.815000 3.560000 11.985000 ;
      RECT 3.390000 12.175000 3.560000 12.345000 ;
      RECT 3.390000 12.535000 3.560000 12.705000 ;
      RECT 3.390000 12.895000 3.560000 13.065000 ;
      RECT 3.390000 13.400000 3.560000 13.570000 ;
      RECT 3.635000  0.250000 3.805000  0.420000 ;
      RECT 3.635000  1.380000 3.805000  1.550000 ;
      RECT 3.635000 15.410000 3.805000 15.580000 ;
      RECT 3.635000 16.540000 3.805000 16.710000 ;
      RECT 3.815000  3.390000 3.985000  3.560000 ;
      RECT 3.815000 13.400000 3.985000 13.570000 ;
      RECT 3.995000  0.250000 4.165000  0.420000 ;
      RECT 3.995000  1.380000 4.165000  1.550000 ;
      RECT 3.995000 15.410000 4.165000 15.580000 ;
      RECT 3.995000 16.540000 4.165000 16.710000 ;
      RECT 4.175000  3.390000 4.345000  3.560000 ;
      RECT 4.175000 13.400000 4.345000 13.570000 ;
      RECT 4.355000  0.250000 4.525000  0.420000 ;
      RECT 4.355000  1.380000 4.525000  1.550000 ;
      RECT 4.355000 15.410000 4.525000 15.580000 ;
      RECT 4.355000 16.540000 4.525000 16.710000 ;
      RECT 4.535000  3.390000 4.705000  3.560000 ;
      RECT 4.535000  4.615000 5.425000 12.345000 ;
      RECT 4.535000 13.400000 4.705000 13.570000 ;
      RECT 4.715000  0.250000 4.885000  0.420000 ;
      RECT 4.715000  1.380000 4.885000  1.550000 ;
      RECT 4.715000 15.410000 4.885000 15.580000 ;
      RECT 4.715000 16.540000 4.885000 16.710000 ;
      RECT 4.895000  3.390000 5.065000  3.560000 ;
      RECT 4.895000 13.400000 5.065000 13.570000 ;
      RECT 5.075000  0.250000 5.245000  0.420000 ;
      RECT 5.075000  1.380000 5.245000  1.550000 ;
      RECT 5.075000 15.410000 5.245000 15.580000 ;
      RECT 5.075000 16.540000 5.245000 16.710000 ;
      RECT 5.255000  3.390000 5.425000  3.560000 ;
      RECT 5.255000 13.400000 5.425000 13.570000 ;
      RECT 5.435000  0.250000 5.605000  0.420000 ;
      RECT 5.435000  1.380000 5.605000  1.550000 ;
      RECT 5.435000 15.410000 5.605000 15.580000 ;
      RECT 5.435000 16.540000 5.605000 16.710000 ;
      RECT 5.615000  3.390000 5.785000  3.560000 ;
      RECT 5.615000 13.400000 5.785000 13.570000 ;
      RECT 5.795000  0.250000 5.965000  0.420000 ;
      RECT 5.795000  1.380000 5.965000  1.550000 ;
      RECT 5.795000 15.410000 5.965000 15.580000 ;
      RECT 5.795000 16.540000 5.965000 16.710000 ;
      RECT 5.975000  3.390000 6.145000  3.560000 ;
      RECT 5.975000 13.400000 6.145000 13.570000 ;
      RECT 6.155000  0.250000 6.325000  0.420000 ;
      RECT 6.155000  1.380000 6.325000  1.550000 ;
      RECT 6.155000 15.410000 6.325000 15.580000 ;
      RECT 6.155000 16.540000 6.325000 16.710000 ;
      RECT 6.400000  3.390000 6.570000  3.560000 ;
      RECT 6.400000  3.895000 6.570000  4.065000 ;
      RECT 6.400000  4.255000 6.570000  4.425000 ;
      RECT 6.400000  4.615000 6.570000  4.785000 ;
      RECT 6.400000  4.975000 6.570000  5.145000 ;
      RECT 6.400000  5.335000 6.570000  5.505000 ;
      RECT 6.400000  5.695000 6.570000  5.865000 ;
      RECT 6.400000  6.055000 6.570000  6.225000 ;
      RECT 6.400000  6.415000 6.570000  6.585000 ;
      RECT 6.400000  6.775000 6.570000  6.945000 ;
      RECT 6.400000  7.135000 6.570000  7.305000 ;
      RECT 6.400000  7.495000 6.570000  7.665000 ;
      RECT 6.400000  7.855000 6.570000  8.025000 ;
      RECT 6.400000  8.215000 6.570000  8.385000 ;
      RECT 6.400000  8.575000 6.570000  8.745000 ;
      RECT 6.400000  8.935000 6.570000  9.105000 ;
      RECT 6.400000  9.295000 6.570000  9.465000 ;
      RECT 6.400000  9.655000 6.570000  9.825000 ;
      RECT 6.400000 10.015000 6.570000 10.185000 ;
      RECT 6.400000 10.375000 6.570000 10.545000 ;
      RECT 6.400000 10.735000 6.570000 10.905000 ;
      RECT 6.400000 11.095000 6.570000 11.265000 ;
      RECT 6.400000 11.455000 6.570000 11.625000 ;
      RECT 6.400000 11.815000 6.570000 11.985000 ;
      RECT 6.400000 12.175000 6.570000 12.345000 ;
      RECT 6.400000 12.535000 6.570000 12.705000 ;
      RECT 6.400000 12.895000 6.570000 13.065000 ;
      RECT 6.400000 13.400000 6.570000 13.570000 ;
      RECT 6.515000  0.250000 6.685000  0.420000 ;
      RECT 6.515000  1.380000 6.685000  1.550000 ;
      RECT 6.515000 15.410000 6.685000 15.580000 ;
      RECT 6.515000 16.540000 6.685000 16.710000 ;
      RECT 6.875000  0.250000 7.045000  0.420000 ;
      RECT 6.875000  1.380000 7.045000  1.550000 ;
      RECT 6.875000 15.410000 7.045000 15.580000 ;
      RECT 6.875000 16.540000 7.045000 16.710000 ;
      RECT 7.235000  0.250000 7.405000  0.420000 ;
      RECT 7.235000  1.380000 7.405000  1.550000 ;
      RECT 7.235000 15.410000 7.405000 15.580000 ;
      RECT 7.235000 16.540000 7.405000 16.710000 ;
      RECT 7.595000  0.250000 7.765000  0.420000 ;
      RECT 7.595000  1.380000 7.765000  1.550000 ;
      RECT 7.595000 15.410000 7.765000 15.580000 ;
      RECT 7.595000 16.540000 7.765000 16.710000 ;
      RECT 7.955000  0.250000 8.125000  0.420000 ;
      RECT 7.955000  1.380000 8.125000  1.550000 ;
      RECT 7.955000 15.410000 8.125000 15.580000 ;
      RECT 7.955000 16.540000 8.125000 16.710000 ;
      RECT 8.315000  0.250000 8.485000  0.420000 ;
      RECT 8.315000 16.540000 8.485000 16.710000 ;
      RECT 8.410000  1.380000 8.580000  1.550000 ;
      RECT 8.410000  1.915000 8.580000  2.085000 ;
      RECT 8.410000  2.275000 8.580000  2.445000 ;
      RECT 8.410000  2.635000 8.580000  2.805000 ;
      RECT 8.410000  2.995000 8.580000  3.165000 ;
      RECT 8.410000  3.355000 8.580000  3.525000 ;
      RECT 8.410000  3.715000 8.580000  3.885000 ;
      RECT 8.410000  4.075000 8.580000  4.245000 ;
      RECT 8.410000  4.435000 8.580000  4.605000 ;
      RECT 8.410000  4.795000 8.580000  4.965000 ;
      RECT 8.410000  5.155000 8.580000  5.325000 ;
      RECT 8.410000  5.515000 8.580000  5.685000 ;
      RECT 8.410000  5.875000 8.580000  6.045000 ;
      RECT 8.410000  6.235000 8.580000  6.405000 ;
      RECT 8.410000  6.595000 8.580000  6.765000 ;
      RECT 8.410000  6.955000 8.580000  7.125000 ;
      RECT 8.410000  7.315000 8.580000  7.485000 ;
      RECT 8.410000  7.675000 8.580000  7.845000 ;
      RECT 8.410000  8.035000 8.580000  8.205000 ;
      RECT 8.410000  8.395000 8.580000  8.565000 ;
      RECT 8.410000  8.755000 8.580000  8.925000 ;
      RECT 8.410000  9.115000 8.580000  9.285000 ;
      RECT 8.410000  9.475000 8.580000  9.645000 ;
      RECT 8.410000  9.835000 8.580000 10.005000 ;
      RECT 8.410000 10.195000 8.580000 10.365000 ;
      RECT 8.410000 10.555000 8.580000 10.725000 ;
      RECT 8.410000 10.915000 8.580000 11.085000 ;
      RECT 8.410000 11.275000 8.580000 11.445000 ;
      RECT 8.410000 11.635000 8.580000 11.805000 ;
      RECT 8.410000 11.995000 8.580000 12.165000 ;
      RECT 8.410000 12.355000 8.580000 12.525000 ;
      RECT 8.410000 12.715000 8.580000 12.885000 ;
      RECT 8.410000 13.075000 8.580000 13.245000 ;
      RECT 8.410000 13.435000 8.580000 13.605000 ;
      RECT 8.410000 13.795000 8.580000 13.965000 ;
      RECT 8.410000 14.155000 8.580000 14.325000 ;
      RECT 8.410000 14.515000 8.580000 14.685000 ;
      RECT 8.410000 14.875000 8.580000 15.045000 ;
      RECT 8.410000 15.410000 8.580000 15.580000 ;
      RECT 8.675000  0.250000 8.845000  0.420000 ;
      RECT 8.675000 16.540000 8.845000 16.710000 ;
      RECT 9.035000  0.250000 9.205000  0.420000 ;
      RECT 9.035000 16.540000 9.205000 16.710000 ;
      RECT 9.540000  0.250000 9.710000  0.420000 ;
      RECT 9.540000  0.655000 9.710000  0.825000 ;
      RECT 9.540000  1.015000 9.710000  1.185000 ;
      RECT 9.540000  1.375000 9.710000  1.545000 ;
      RECT 9.540000  1.735000 9.710000  1.905000 ;
      RECT 9.540000  2.095000 9.710000  2.265000 ;
      RECT 9.540000  2.455000 9.710000  2.625000 ;
      RECT 9.540000  2.815000 9.710000  2.985000 ;
      RECT 9.540000  3.175000 9.710000  3.345000 ;
      RECT 9.540000  3.535000 9.710000  3.705000 ;
      RECT 9.540000  3.895000 9.710000  4.065000 ;
      RECT 9.540000  4.255000 9.710000  4.425000 ;
      RECT 9.540000  4.615000 9.710000  4.785000 ;
      RECT 9.540000  4.975000 9.710000  5.145000 ;
      RECT 9.540000  5.335000 9.710000  5.505000 ;
      RECT 9.540000  5.695000 9.710000  5.865000 ;
      RECT 9.540000  6.055000 9.710000  6.225000 ;
      RECT 9.540000  6.415000 9.710000  6.585000 ;
      RECT 9.540000  6.775000 9.710000  6.945000 ;
      RECT 9.540000  7.135000 9.710000  7.305000 ;
      RECT 9.540000  7.495000 9.710000  7.665000 ;
      RECT 9.540000  7.855000 9.710000  8.025000 ;
      RECT 9.540000  8.215000 9.710000  8.385000 ;
      RECT 9.540000  8.575000 9.710000  8.745000 ;
      RECT 9.540000  8.935000 9.710000  9.105000 ;
      RECT 9.540000  9.295000 9.710000  9.465000 ;
      RECT 9.540000  9.655000 9.710000  9.825000 ;
      RECT 9.540000 10.015000 9.710000 10.185000 ;
      RECT 9.540000 10.375000 9.710000 10.545000 ;
      RECT 9.540000 10.735000 9.710000 10.905000 ;
      RECT 9.540000 11.095000 9.710000 11.265000 ;
      RECT 9.540000 11.455000 9.710000 11.625000 ;
      RECT 9.540000 11.815000 9.710000 11.985000 ;
      RECT 9.540000 12.175000 9.710000 12.345000 ;
      RECT 9.540000 12.535000 9.710000 12.705000 ;
      RECT 9.540000 12.895000 9.710000 13.065000 ;
      RECT 9.540000 13.255000 9.710000 13.425000 ;
      RECT 9.540000 13.615000 9.710000 13.785000 ;
      RECT 9.540000 13.975000 9.710000 14.145000 ;
      RECT 9.540000 14.335000 9.710000 14.505000 ;
      RECT 9.540000 14.695000 9.710000 14.865000 ;
      RECT 9.540000 15.055000 9.710000 15.225000 ;
      RECT 9.540000 15.415000 9.710000 15.585000 ;
      RECT 9.540000 15.775000 9.710000 15.945000 ;
      RECT 9.540000 16.135000 9.710000 16.305000 ;
      RECT 9.540000 16.540000 9.710000 16.710000 ;
    LAYER met1 ;
      RECT 0.190000  0.190000 9.770000  0.480000 ;
      RECT 0.190000  0.480000 0.480000 16.480000 ;
      RECT 0.190000 16.480000 9.770000 16.770000 ;
      RECT 1.320000  1.320000 8.640000  1.610000 ;
      RECT 1.320000  1.610000 1.610000 15.350000 ;
      RECT 1.320000 15.350000 8.640000 15.640000 ;
      RECT 3.330000  3.330000 6.630000  3.620000 ;
      RECT 3.330000  3.620000 3.620000 13.340000 ;
      RECT 3.330000 13.340000 6.630000 13.630000 ;
      RECT 4.475000  4.555000 5.485000 12.405000 ;
      RECT 6.340000  3.620000 6.630000 13.340000 ;
      RECT 8.350000  1.610000 8.640000 15.350000 ;
      RECT 9.480000  0.480000 9.770000 16.480000 ;
  END
END sky130_fd_pr__rf_npn_05v5_W1p00L8p00
END LIBRARY
