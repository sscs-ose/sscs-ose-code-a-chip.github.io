# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  1.500000 BY  1.960000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.235200 ;
    PORT
      LAYER met2 ;
        RECT 0.635000 0.280000 0.895000 0.920000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.252000 ;
    PORT
      LAYER met1 ;
        RECT 0.440000 1.205000 1.090000 1.495000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.445200 ;
    PORT
      LAYER met1 ;
        RECT 0.220000 -0.445000 1.310000 -0.145000 ;
        RECT 0.220000 -0.145000 0.450000  0.945000 ;
        RECT 1.080000 -0.145000 1.310000  0.945000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.250000 0.255000 0.420000 0.945000 ;
      RECT 0.430000 1.175000 1.100000 1.515000 ;
      RECT 0.680000 0.255000 0.850000 0.945000 ;
      RECT 1.110000 0.255000 1.280000 0.945000 ;
    LAYER mcon ;
      RECT 0.250000 0.335000 0.420000 0.505000 ;
      RECT 0.250000 0.695000 0.420000 0.865000 ;
      RECT 0.500000 1.265000 0.670000 1.435000 ;
      RECT 0.680000 0.335000 0.850000 0.505000 ;
      RECT 0.680000 0.695000 0.850000 0.865000 ;
      RECT 0.860000 1.265000 1.030000 1.435000 ;
      RECT 1.110000 0.335000 1.280000 0.505000 ;
      RECT 1.110000 0.695000 1.280000 0.865000 ;
    LAYER met1 ;
      RECT 0.635000 0.255000 0.895000 0.945000 ;
    LAYER via ;
      RECT 0.635000 0.310000 0.895000 0.570000 ;
      RECT 0.635000 0.630000 0.895000 0.890000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15
END LIBRARY
