# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield ;
  ORIGIN  0.440000  0.000000 ;
  SIZE  8.580000 BY  7.840000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT -0.440000 0.000000  8.140000 0.320000 ;
        RECT -0.440000 0.320000 -0.170000 7.380000 ;
        RECT  0.280000 0.320000  0.420000 7.380000 ;
        RECT  0.840000 0.320000  0.980000 7.380000 ;
        RECT  1.400000 0.320000  1.540000 7.380000 ;
        RECT  1.960000 0.320000  2.100000 7.380000 ;
        RECT  2.520000 0.320000  2.660000 7.380000 ;
        RECT  3.080000 0.320000  3.220000 7.380000 ;
        RECT  3.640000 0.320000  3.780000 7.380000 ;
        RECT  4.200000 0.320000  4.340000 7.380000 ;
        RECT  4.760000 0.320000  4.900000 7.380000 ;
        RECT  5.320000 0.320000  5.460000 7.380000 ;
        RECT  5.880000 0.320000  6.020000 7.380000 ;
        RECT  6.440000 0.320000  6.580000 7.380000 ;
        RECT  7.000000 0.320000  7.140000 7.380000 ;
        RECT  7.560000 0.320000  7.700000 7.380000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT -0.440000 7.520000 8.140000 7.840000 ;
        RECT  0.000000 0.460000 0.140000 7.520000 ;
        RECT  0.560000 0.460000 0.700000 7.520000 ;
        RECT  1.120000 0.460000 1.260000 7.520000 ;
        RECT  1.680000 0.460000 1.820000 7.520000 ;
        RECT  2.240000 0.460000 2.380000 7.520000 ;
        RECT  2.800000 0.460000 2.940000 7.520000 ;
        RECT  3.360000 0.460000 3.500000 7.520000 ;
        RECT  3.920000 0.460000 4.060000 7.520000 ;
        RECT  4.480000 0.460000 4.620000 7.520000 ;
        RECT  5.040000 0.460000 5.180000 7.520000 ;
        RECT  5.600000 0.460000 5.740000 7.520000 ;
        RECT  6.160000 0.460000 6.300000 7.520000 ;
        RECT  6.720000 0.460000 6.860000 7.520000 ;
        RECT  7.280000 0.460000 7.420000 7.520000 ;
        RECT  7.870000 0.460000 8.140000 7.520000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 3.805000 3.825000 3.880000 3.915000 ;
    END
  END SUB
  OBS
    LAYER met1 ;
      RECT -0.440000 0.000000  8.140000 0.320000 ;
      RECT -0.440000 0.320000 -0.170000 7.380000 ;
      RECT -0.440000 7.520000  8.140000 7.840000 ;
      RECT  0.000000 0.320000  0.140000 7.380000 ;
      RECT  0.280000 0.460000  0.420000 7.520000 ;
      RECT  0.560000 0.320000  0.700000 7.380000 ;
      RECT  0.840000 0.460000  0.980000 7.520000 ;
      RECT  1.120000 0.320000  1.260000 7.380000 ;
      RECT  1.400000 0.460000  1.540000 7.520000 ;
      RECT  1.680000 0.320000  1.820000 7.380000 ;
      RECT  1.960000 0.460000  2.100000 7.520000 ;
      RECT  2.240000 0.320000  2.380000 7.380000 ;
      RECT  2.520000 0.460000  2.660000 7.520000 ;
      RECT  2.800000 0.320000  2.940000 7.380000 ;
      RECT  3.080000 0.460000  3.220000 7.520000 ;
      RECT  3.360000 0.320000  3.500000 7.380000 ;
      RECT  3.640000 0.460000  3.780000 7.520000 ;
      RECT  3.920000 0.320000  4.060000 7.380000 ;
      RECT  4.200000 0.460000  4.340000 7.520000 ;
      RECT  4.480000 0.320000  4.620000 7.380000 ;
      RECT  4.760000 0.460000  4.900000 7.520000 ;
      RECT  5.040000 0.320000  5.180000 7.380000 ;
      RECT  5.320000 0.460000  5.460000 7.520000 ;
      RECT  5.600000 0.320000  5.740000 7.380000 ;
      RECT  5.880000 0.460000  6.020000 7.520000 ;
      RECT  6.160000 0.320000  6.300000 7.380000 ;
      RECT  6.440000 0.460000  6.580000 7.520000 ;
      RECT  6.720000 0.320000  6.860000 7.380000 ;
      RECT  7.000000 0.460000  7.140000 7.520000 ;
      RECT  7.280000 0.320000  7.420000 7.380000 ;
      RECT  7.560000 0.460000  7.700000 7.520000 ;
      RECT  7.870000 0.460000  8.140000 7.520000 ;
    LAYER via ;
      RECT -0.435000 0.265000 -0.175000 0.525000 ;
      RECT -0.435000 0.585000 -0.175000 0.845000 ;
      RECT -0.435000 0.905000 -0.175000 1.165000 ;
      RECT -0.435000 1.225000 -0.175000 1.485000 ;
      RECT -0.435000 1.545000 -0.175000 1.805000 ;
      RECT -0.435000 1.865000 -0.175000 2.125000 ;
      RECT -0.435000 2.185000 -0.175000 2.445000 ;
      RECT -0.435000 2.505000 -0.175000 2.765000 ;
      RECT -0.435000 2.825000 -0.175000 3.085000 ;
      RECT -0.435000 3.145000 -0.175000 3.405000 ;
      RECT -0.435000 3.465000 -0.175000 3.725000 ;
      RECT -0.435000 3.785000 -0.175000 4.045000 ;
      RECT -0.435000 4.105000 -0.175000 4.365000 ;
      RECT -0.435000 4.425000 -0.175000 4.685000 ;
      RECT -0.435000 4.745000 -0.175000 5.005000 ;
      RECT -0.435000 5.065000 -0.175000 5.325000 ;
      RECT -0.435000 5.385000 -0.175000 5.645000 ;
      RECT -0.435000 5.705000 -0.175000 5.965000 ;
      RECT -0.435000 6.025000 -0.175000 6.285000 ;
      RECT -0.435000 6.345000 -0.175000 6.605000 ;
      RECT -0.435000 6.665000 -0.175000 6.925000 ;
      RECT -0.435000 6.985000 -0.175000 7.245000 ;
      RECT -0.060000 0.030000  0.200000 0.290000 ;
      RECT -0.060000 7.550000  0.200000 7.810000 ;
      RECT  0.260000 0.030000  0.520000 0.290000 ;
      RECT  0.260000 7.550000  0.520000 7.810000 ;
      RECT  0.580000 0.030000  0.840000 0.290000 ;
      RECT  0.580000 7.550000  0.840000 7.810000 ;
      RECT  0.900000 0.030000  1.160000 0.290000 ;
      RECT  0.900000 7.550000  1.160000 7.810000 ;
      RECT  1.220000 0.030000  1.480000 0.290000 ;
      RECT  1.220000 7.550000  1.480000 7.810000 ;
      RECT  1.540000 0.030000  1.800000 0.290000 ;
      RECT  1.540000 7.550000  1.800000 7.810000 ;
      RECT  1.860000 0.030000  2.120000 0.290000 ;
      RECT  1.860000 7.550000  2.120000 7.810000 ;
      RECT  2.180000 0.030000  2.440000 0.290000 ;
      RECT  2.180000 7.550000  2.440000 7.810000 ;
      RECT  2.500000 0.030000  2.760000 0.290000 ;
      RECT  2.500000 7.550000  2.760000 7.810000 ;
      RECT  2.820000 0.030000  3.080000 0.290000 ;
      RECT  2.820000 7.550000  3.080000 7.810000 ;
      RECT  3.140000 0.030000  3.400000 0.290000 ;
      RECT  3.140000 7.550000  3.400000 7.810000 ;
      RECT  3.460000 0.030000  3.720000 0.290000 ;
      RECT  3.460000 7.550000  3.720000 7.810000 ;
      RECT  3.780000 0.030000  4.040000 0.290000 ;
      RECT  3.780000 7.550000  4.040000 7.810000 ;
      RECT  4.100000 0.030000  4.360000 0.290000 ;
      RECT  4.100000 7.550000  4.360000 7.810000 ;
      RECT  4.420000 0.030000  4.680000 0.290000 ;
      RECT  4.420000 7.550000  4.680000 7.810000 ;
      RECT  4.740000 0.030000  5.000000 0.290000 ;
      RECT  4.740000 7.550000  5.000000 7.810000 ;
      RECT  5.060000 0.030000  5.320000 0.290000 ;
      RECT  5.060000 7.550000  5.320000 7.810000 ;
      RECT  5.380000 0.030000  5.640000 0.290000 ;
      RECT  5.380000 7.550000  5.640000 7.810000 ;
      RECT  5.700000 0.030000  5.960000 0.290000 ;
      RECT  5.700000 7.550000  5.960000 7.810000 ;
      RECT  6.020000 0.030000  6.280000 0.290000 ;
      RECT  6.020000 7.550000  6.280000 7.810000 ;
      RECT  6.340000 0.030000  6.600000 0.290000 ;
      RECT  6.340000 7.550000  6.600000 7.810000 ;
      RECT  6.660000 0.030000  6.920000 0.290000 ;
      RECT  6.660000 7.550000  6.920000 7.810000 ;
      RECT  6.980000 0.030000  7.240000 0.290000 ;
      RECT  6.980000 7.550000  7.240000 7.810000 ;
      RECT  7.300000 0.030000  7.560000 0.290000 ;
      RECT  7.300000 7.550000  7.560000 7.810000 ;
      RECT  7.620000 0.030000  7.880000 0.290000 ;
      RECT  7.620000 7.550000  7.880000 7.810000 ;
      RECT  7.875000 0.490000  8.135000 0.750000 ;
      RECT  7.875000 0.810000  8.135000 1.070000 ;
      RECT  7.875000 1.130000  8.135000 1.390000 ;
      RECT  7.875000 1.450000  8.135000 1.710000 ;
      RECT  7.875000 1.770000  8.135000 2.030000 ;
      RECT  7.875000 2.090000  8.135000 2.350000 ;
      RECT  7.875000 2.410000  8.135000 2.670000 ;
      RECT  7.875000 2.730000  8.135000 2.990000 ;
      RECT  7.875000 3.050000  8.135000 3.310000 ;
      RECT  7.875000 3.370000  8.135000 3.630000 ;
      RECT  7.875000 3.690000  8.135000 3.950000 ;
      RECT  7.875000 4.010000  8.135000 4.270000 ;
      RECT  7.875000 4.330000  8.135000 4.590000 ;
      RECT  7.875000 4.650000  8.135000 4.910000 ;
      RECT  7.875000 4.970000  8.135000 5.230000 ;
      RECT  7.875000 5.290000  8.135000 5.550000 ;
      RECT  7.875000 5.610000  8.135000 5.870000 ;
      RECT  7.875000 5.930000  8.135000 6.190000 ;
      RECT  7.875000 6.250000  8.135000 6.510000 ;
      RECT  7.875000 6.570000  8.135000 6.830000 ;
      RECT  7.875000 6.890000  8.135000 7.150000 ;
      RECT  7.875000 7.210000  8.135000 7.470000 ;
  END
END sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield
END LIBRARY
