* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


* Top level circuit sky130_fd_pr__esd_rf_nfet_20v0_iec_21vW60p00
X0 dw_n700_n714# SUBS SUBS SUBS sky130_fd_pr__nfet_20v0 w=3e+07u l=1.5e+06u
X1 dw_n700_n714# SUBS SUBS SUBS sky130_fd_pr__nfet_20v0 w=3e+07u l=1.5e+06u
.end
