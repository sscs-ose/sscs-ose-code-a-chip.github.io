# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50 ;
  ORIGIN -0.050000  0.000000 ;
  SIZE  5.020000 BY  5.970000 ;
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 3.110000 5.070000 5.470000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  10.099999 ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.100000 4.085000 0.270000 ;
        RECT 1.035000 5.700000 4.085000 5.870000 ;
      LAYER mcon ;
        RECT 1.215000 0.100000 1.385000 0.270000 ;
        RECT 1.215000 5.700000 1.385000 5.870000 ;
        RECT 1.575000 0.100000 1.745000 0.270000 ;
        RECT 1.575000 5.700000 1.745000 5.870000 ;
        RECT 1.935000 0.100000 2.105000 0.270000 ;
        RECT 1.935000 5.700000 2.105000 5.870000 ;
        RECT 2.295000 0.100000 2.465000 0.270000 ;
        RECT 2.295000 5.700000 2.465000 5.870000 ;
        RECT 2.655000 0.100000 2.825000 0.270000 ;
        RECT 2.655000 5.700000 2.825000 5.870000 ;
        RECT 3.015000 0.100000 3.185000 0.270000 ;
        RECT 3.015000 5.700000 3.185000 5.870000 ;
        RECT 3.375000 0.100000 3.545000 0.270000 ;
        RECT 3.375000 5.700000 3.545000 5.870000 ;
        RECT 3.735000 0.100000 3.905000 0.270000 ;
        RECT 3.735000 5.700000 3.905000 5.870000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.155000 0.000000 3.965000 0.330000 ;
        RECT 1.155000 5.640000 3.965000 5.970000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.500000 5.070000 2.860000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.464500 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.500000 0.475000 5.470000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.650000 0.500000 4.945000 5.470000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.560000 0.410000 5.410000 ;
      RECT 0.915000 0.440000 1.085000 5.530000 ;
      RECT 1.695000 0.440000 1.865000 5.530000 ;
      RECT 2.475000 0.440000 2.645000 5.530000 ;
      RECT 3.255000 0.440000 3.425000 5.530000 ;
      RECT 4.035000 0.440000 4.205000 5.530000 ;
      RECT 4.710000 0.560000 4.880000 5.410000 ;
    LAYER mcon ;
      RECT 0.240000 0.920000 0.410000 1.090000 ;
      RECT 0.240000 1.280000 0.410000 1.450000 ;
      RECT 0.240000 1.640000 0.410000 1.810000 ;
      RECT 0.240000 2.000000 0.410000 2.170000 ;
      RECT 0.240000 2.360000 0.410000 2.530000 ;
      RECT 0.240000 2.720000 0.410000 2.890000 ;
      RECT 0.240000 3.080000 0.410000 3.250000 ;
      RECT 0.240000 3.440000 0.410000 3.610000 ;
      RECT 0.240000 3.800000 0.410000 3.970000 ;
      RECT 0.240000 4.160000 0.410000 4.330000 ;
      RECT 0.240000 4.520000 0.410000 4.690000 ;
      RECT 0.240000 4.880000 0.410000 5.050000 ;
      RECT 0.240000 5.240000 0.410000 5.410000 ;
      RECT 0.915000 0.560000 1.085000 0.730000 ;
      RECT 0.915000 0.920000 1.085000 1.090000 ;
      RECT 0.915000 1.280000 1.085000 1.450000 ;
      RECT 0.915000 1.640000 1.085000 1.810000 ;
      RECT 0.915000 2.000000 1.085000 2.170000 ;
      RECT 0.915000 2.360000 1.085000 2.530000 ;
      RECT 0.915000 2.720000 1.085000 2.890000 ;
      RECT 0.915000 3.080000 1.085000 3.250000 ;
      RECT 0.915000 3.440000 1.085000 3.610000 ;
      RECT 0.915000 3.800000 1.085000 3.970000 ;
      RECT 0.915000 4.160000 1.085000 4.330000 ;
      RECT 0.915000 4.520000 1.085000 4.690000 ;
      RECT 0.915000 4.880000 1.085000 5.050000 ;
      RECT 0.915000 5.240000 1.085000 5.410000 ;
      RECT 1.695000 0.560000 1.865000 0.730000 ;
      RECT 1.695000 0.920000 1.865000 1.090000 ;
      RECT 1.695000 1.280000 1.865000 1.450000 ;
      RECT 1.695000 1.640000 1.865000 1.810000 ;
      RECT 1.695000 2.000000 1.865000 2.170000 ;
      RECT 1.695000 2.360000 1.865000 2.530000 ;
      RECT 1.695000 2.720000 1.865000 2.890000 ;
      RECT 1.695000 3.080000 1.865000 3.250000 ;
      RECT 1.695000 3.440000 1.865000 3.610000 ;
      RECT 1.695000 3.800000 1.865000 3.970000 ;
      RECT 1.695000 4.160000 1.865000 4.330000 ;
      RECT 1.695000 4.520000 1.865000 4.690000 ;
      RECT 1.695000 4.880000 1.865000 5.050000 ;
      RECT 1.695000 5.240000 1.865000 5.410000 ;
      RECT 2.475000 0.560000 2.645000 0.730000 ;
      RECT 2.475000 0.920000 2.645000 1.090000 ;
      RECT 2.475000 1.280000 2.645000 1.450000 ;
      RECT 2.475000 1.640000 2.645000 1.810000 ;
      RECT 2.475000 2.000000 2.645000 2.170000 ;
      RECT 2.475000 2.360000 2.645000 2.530000 ;
      RECT 2.475000 2.720000 2.645000 2.890000 ;
      RECT 2.475000 3.080000 2.645000 3.250000 ;
      RECT 2.475000 3.440000 2.645000 3.610000 ;
      RECT 2.475000 3.800000 2.645000 3.970000 ;
      RECT 2.475000 4.160000 2.645000 4.330000 ;
      RECT 2.475000 4.520000 2.645000 4.690000 ;
      RECT 2.475000 4.880000 2.645000 5.050000 ;
      RECT 2.475000 5.240000 2.645000 5.410000 ;
      RECT 3.255000 0.560000 3.425000 0.730000 ;
      RECT 3.255000 0.920000 3.425000 1.090000 ;
      RECT 3.255000 1.280000 3.425000 1.450000 ;
      RECT 3.255000 1.640000 3.425000 1.810000 ;
      RECT 3.255000 2.000000 3.425000 2.170000 ;
      RECT 3.255000 2.360000 3.425000 2.530000 ;
      RECT 3.255000 2.720000 3.425000 2.890000 ;
      RECT 3.255000 3.080000 3.425000 3.250000 ;
      RECT 3.255000 3.440000 3.425000 3.610000 ;
      RECT 3.255000 3.800000 3.425000 3.970000 ;
      RECT 3.255000 4.160000 3.425000 4.330000 ;
      RECT 3.255000 4.520000 3.425000 4.690000 ;
      RECT 3.255000 4.880000 3.425000 5.050000 ;
      RECT 3.255000 5.240000 3.425000 5.410000 ;
      RECT 4.035000 0.560000 4.205000 0.730000 ;
      RECT 4.035000 0.920000 4.205000 1.090000 ;
      RECT 4.035000 1.280000 4.205000 1.450000 ;
      RECT 4.035000 1.640000 4.205000 1.810000 ;
      RECT 4.035000 2.000000 4.205000 2.170000 ;
      RECT 4.035000 2.360000 4.205000 2.530000 ;
      RECT 4.035000 2.720000 4.205000 2.890000 ;
      RECT 4.035000 3.080000 4.205000 3.250000 ;
      RECT 4.035000 3.440000 4.205000 3.610000 ;
      RECT 4.035000 3.800000 4.205000 3.970000 ;
      RECT 4.035000 4.160000 4.205000 4.330000 ;
      RECT 4.035000 4.520000 4.205000 4.690000 ;
      RECT 4.035000 4.880000 4.205000 5.050000 ;
      RECT 4.035000 5.240000 4.205000 5.410000 ;
      RECT 4.710000 0.920000 4.880000 1.090000 ;
      RECT 4.710000 1.280000 4.880000 1.450000 ;
      RECT 4.710000 1.640000 4.880000 1.810000 ;
      RECT 4.710000 2.000000 4.880000 2.170000 ;
      RECT 4.710000 2.360000 4.880000 2.530000 ;
      RECT 4.710000 2.720000 4.880000 2.890000 ;
      RECT 4.710000 3.080000 4.880000 3.250000 ;
      RECT 4.710000 3.440000 4.880000 3.610000 ;
      RECT 4.710000 3.800000 4.880000 3.970000 ;
      RECT 4.710000 4.160000 4.880000 4.330000 ;
      RECT 4.710000 4.520000 4.880000 4.690000 ;
      RECT 4.710000 4.880000 4.880000 5.050000 ;
      RECT 4.710000 5.240000 4.880000 5.410000 ;
    LAYER met1 ;
      RECT 0.870000 0.500000 1.130000 5.470000 ;
      RECT 1.650000 0.500000 1.910000 5.470000 ;
      RECT 2.430000 0.500000 2.690000 5.470000 ;
      RECT 3.210000 0.500000 3.470000 5.470000 ;
      RECT 3.990000 0.500000 4.250000 5.470000 ;
    LAYER via ;
      RECT 0.870000 0.530000 1.130000 0.790000 ;
      RECT 0.870000 0.850000 1.130000 1.110000 ;
      RECT 0.870000 1.170000 1.130000 1.430000 ;
      RECT 0.870000 1.490000 1.130000 1.750000 ;
      RECT 0.870000 1.810000 1.130000 2.070000 ;
      RECT 0.870000 2.130000 1.130000 2.390000 ;
      RECT 0.870000 2.450000 1.130000 2.710000 ;
      RECT 1.650000 3.260000 1.910000 3.520000 ;
      RECT 1.650000 3.580000 1.910000 3.840000 ;
      RECT 1.650000 3.900000 1.910000 4.160000 ;
      RECT 1.650000 4.220000 1.910000 4.480000 ;
      RECT 1.650000 4.540000 1.910000 4.800000 ;
      RECT 1.650000 4.860000 1.910000 5.120000 ;
      RECT 1.650000 5.180000 1.910000 5.440000 ;
      RECT 2.430000 0.530000 2.690000 0.790000 ;
      RECT 2.430000 0.850000 2.690000 1.110000 ;
      RECT 2.430000 1.170000 2.690000 1.430000 ;
      RECT 2.430000 1.490000 2.690000 1.750000 ;
      RECT 2.430000 1.810000 2.690000 2.070000 ;
      RECT 2.430000 2.130000 2.690000 2.390000 ;
      RECT 2.430000 2.450000 2.690000 2.710000 ;
      RECT 3.210000 3.260000 3.470000 3.520000 ;
      RECT 3.210000 3.580000 3.470000 3.840000 ;
      RECT 3.210000 3.900000 3.470000 4.160000 ;
      RECT 3.210000 4.220000 3.470000 4.480000 ;
      RECT 3.210000 4.540000 3.470000 4.800000 ;
      RECT 3.210000 4.860000 3.470000 5.120000 ;
      RECT 3.210000 5.180000 3.470000 5.440000 ;
      RECT 3.990000 0.530000 4.250000 0.790000 ;
      RECT 3.990000 0.850000 4.250000 1.110000 ;
      RECT 3.990000 1.170000 4.250000 1.430000 ;
      RECT 3.990000 1.490000 4.250000 1.750000 ;
      RECT 3.990000 1.810000 4.250000 2.070000 ;
      RECT 3.990000 2.130000 4.250000 2.390000 ;
      RECT 3.990000 2.450000 4.250000 2.710000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50
END LIBRARY
