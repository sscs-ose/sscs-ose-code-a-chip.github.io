# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF06W2p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF06W2p00L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  3.190000 BY  3.120000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.680000 ;
    PORT
      LAYER met3 ;
        RECT 0.570000 1.375000 0.900000 1.815000 ;
        RECT 0.570000 1.815000 2.620000 2.145000 ;
        RECT 1.430000 1.375000 1.760000 1.815000 ;
        RECT 2.290000 1.375000 2.620000 1.815000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.800000 ;
    PORT
      LAYER met1 ;
        RECT 0.550000 2.365000 2.640000 2.655000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.180000 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.445000 3.000000 -0.145000 ;
        RECT 0.190000 -0.145000 0.420000  2.105000 ;
        RECT 1.050000 -0.145000 1.280000  2.105000 ;
        RECT 1.910000 -0.145000 2.140000  2.105000 ;
        RECT 2.770000 -0.145000 3.000000  2.105000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.255000 0.390000 2.105000 ;
      RECT 0.580000 2.335000 2.610000 2.675000 ;
      RECT 0.650000 0.255000 0.820000 2.105000 ;
      RECT 1.080000 0.255000 1.250000 2.105000 ;
      RECT 1.510000 0.255000 1.680000 2.105000 ;
      RECT 1.940000 0.255000 2.110000 2.105000 ;
      RECT 2.370000 0.255000 2.540000 2.105000 ;
      RECT 2.800000 0.255000 2.970000 2.105000 ;
    LAYER mcon ;
      RECT 0.220000 0.375000 0.390000 0.545000 ;
      RECT 0.220000 0.735000 0.390000 0.905000 ;
      RECT 0.220000 1.095000 0.390000 1.265000 ;
      RECT 0.220000 1.455000 0.390000 1.625000 ;
      RECT 0.220000 1.815000 0.390000 1.985000 ;
      RECT 0.610000 2.425000 0.780000 2.595000 ;
      RECT 0.650000 0.375000 0.820000 0.545000 ;
      RECT 0.650000 0.735000 0.820000 0.905000 ;
      RECT 0.650000 1.095000 0.820000 1.265000 ;
      RECT 0.650000 1.455000 0.820000 1.625000 ;
      RECT 0.650000 1.815000 0.820000 1.985000 ;
      RECT 0.970000 2.425000 1.140000 2.595000 ;
      RECT 1.080000 0.375000 1.250000 0.545000 ;
      RECT 1.080000 0.735000 1.250000 0.905000 ;
      RECT 1.080000 1.095000 1.250000 1.265000 ;
      RECT 1.080000 1.455000 1.250000 1.625000 ;
      RECT 1.080000 1.815000 1.250000 1.985000 ;
      RECT 1.330000 2.425000 1.500000 2.595000 ;
      RECT 1.510000 0.375000 1.680000 0.545000 ;
      RECT 1.510000 0.735000 1.680000 0.905000 ;
      RECT 1.510000 1.095000 1.680000 1.265000 ;
      RECT 1.510000 1.455000 1.680000 1.625000 ;
      RECT 1.510000 1.815000 1.680000 1.985000 ;
      RECT 1.690000 2.425000 1.860000 2.595000 ;
      RECT 1.940000 0.375000 2.110000 0.545000 ;
      RECT 1.940000 0.735000 2.110000 0.905000 ;
      RECT 1.940000 1.095000 2.110000 1.265000 ;
      RECT 1.940000 1.455000 2.110000 1.625000 ;
      RECT 1.940000 1.815000 2.110000 1.985000 ;
      RECT 2.050000 2.425000 2.220000 2.595000 ;
      RECT 2.370000 0.375000 2.540000 0.545000 ;
      RECT 2.370000 0.735000 2.540000 0.905000 ;
      RECT 2.370000 1.095000 2.540000 1.265000 ;
      RECT 2.370000 1.455000 2.540000 1.625000 ;
      RECT 2.370000 1.815000 2.540000 1.985000 ;
      RECT 2.410000 2.425000 2.580000 2.595000 ;
      RECT 2.800000 0.375000 2.970000 0.545000 ;
      RECT 2.800000 0.735000 2.970000 0.905000 ;
      RECT 2.800000 1.095000 2.970000 1.265000 ;
      RECT 2.800000 1.455000 2.970000 1.625000 ;
      RECT 2.800000 1.815000 2.970000 1.985000 ;
    LAYER met1 ;
      RECT 0.605000 0.255000 0.865000 2.105000 ;
      RECT 1.465000 0.255000 1.725000 2.105000 ;
      RECT 2.325000 0.255000 2.585000 2.105000 ;
    LAYER met2 ;
      RECT 0.570000 1.375000 0.900000 2.145000 ;
      RECT 1.430000 1.375000 1.760000 2.145000 ;
      RECT 2.290000 1.375000 2.620000 2.145000 ;
    LAYER via ;
      RECT 0.605000 1.470000 0.865000 1.730000 ;
      RECT 0.605000 1.790000 0.865000 2.050000 ;
      RECT 1.465000 1.470000 1.725000 1.730000 ;
      RECT 1.465000 1.790000 1.725000 2.050000 ;
      RECT 2.325000 1.470000 2.585000 1.730000 ;
      RECT 2.325000 1.790000 2.585000 2.050000 ;
    LAYER via2 ;
      RECT 0.595000 1.420000 0.875000 1.700000 ;
      RECT 0.595000 1.820000 0.875000 2.100000 ;
      RECT 1.455000 1.420000 1.735000 1.700000 ;
      RECT 1.455000 1.820000 1.735000 2.100000 ;
      RECT 2.315000 1.420000 2.595000 1.700000 ;
      RECT 2.315000 1.820000 2.595000 2.100000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF06W2p00L0p15
END LIBRARY
