** sch_path: /home/evadeltor/half_Miyahara.sch
**.subckt half_Miyahara
M5 net1 Vin- net2 M2N7002 m=1
M1 net1 Vb net2 M2N7002 m=1
M6 GND net2 net3 M2N7002 m=1
M7 GND net4 net3 M2N7002 m=1
M10 GND net2 net5 M2N7002 m=1
M13 net5 net2 VDD DMP2035U m=1
M14 net3 net4 net5 DMP2035U m=1
M16 net2 CLK VDD DMP2035U m=1
**.ends
.GLOBAL GND
.end
