magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< error_p >>
rect -29 62323 29 62329
rect -29 62289 -17 62323
rect -29 62283 29 62289
rect -29 56195 29 56201
rect -29 56161 -17 56195
rect -29 56155 29 56161
rect -29 56087 29 56093
rect -29 56053 -17 56087
rect -29 56047 29 56053
rect -29 49959 29 49965
rect -29 49925 -17 49959
rect -29 49919 29 49925
rect -29 49851 29 49857
rect -29 49817 -17 49851
rect -29 49811 29 49817
rect -29 43723 29 43729
rect -29 43689 -17 43723
rect -29 43683 29 43689
rect -29 43615 29 43621
rect -29 43581 -17 43615
rect -29 43575 29 43581
rect -29 37487 29 37493
rect -29 37453 -17 37487
rect -29 37447 29 37453
rect -29 37379 29 37385
rect -29 37345 -17 37379
rect -29 37339 29 37345
rect -29 31251 29 31257
rect -29 31217 -17 31251
rect -29 31211 29 31217
rect -29 31143 29 31149
rect -29 31109 -17 31143
rect -29 31103 29 31109
rect -29 25015 29 25021
rect -29 24981 -17 25015
rect -29 24975 29 24981
rect -29 24907 29 24913
rect -29 24873 -17 24907
rect -29 24867 29 24873
rect -29 18779 29 18785
rect -29 18745 -17 18779
rect -29 18739 29 18745
rect -29 18671 29 18677
rect -29 18637 -17 18671
rect -29 18631 29 18637
rect -29 12543 29 12549
rect -29 12509 -17 12543
rect -29 12503 29 12509
rect -29 12435 29 12441
rect -29 12401 -17 12435
rect -29 12395 29 12401
rect -29 6307 29 6313
rect -29 6273 -17 6307
rect -29 6267 29 6273
rect -29 6199 29 6205
rect -29 6165 -17 6199
rect -29 6159 29 6165
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -6165 29 -6159
rect -29 -6199 -17 -6165
rect -29 -6205 29 -6199
rect -29 -6273 29 -6267
rect -29 -6307 -17 -6273
rect -29 -6313 29 -6307
rect -29 -12401 29 -12395
rect -29 -12435 -17 -12401
rect -29 -12441 29 -12435
rect -29 -12509 29 -12503
rect -29 -12543 -17 -12509
rect -29 -12549 29 -12543
rect -29 -18637 29 -18631
rect -29 -18671 -17 -18637
rect -29 -18677 29 -18671
rect -29 -18745 29 -18739
rect -29 -18779 -17 -18745
rect -29 -18785 29 -18779
rect -29 -24873 29 -24867
rect -29 -24907 -17 -24873
rect -29 -24913 29 -24907
rect -29 -24981 29 -24975
rect -29 -25015 -17 -24981
rect -29 -25021 29 -25015
rect -29 -31109 29 -31103
rect -29 -31143 -17 -31109
rect -29 -31149 29 -31143
rect -29 -31217 29 -31211
rect -29 -31251 -17 -31217
rect -29 -31257 29 -31251
rect -29 -37345 29 -37339
rect -29 -37379 -17 -37345
rect -29 -37385 29 -37379
rect -29 -37453 29 -37447
rect -29 -37487 -17 -37453
rect -29 -37493 29 -37487
rect -29 -43581 29 -43575
rect -29 -43615 -17 -43581
rect -29 -43621 29 -43615
rect -29 -43689 29 -43683
rect -29 -43723 -17 -43689
rect -29 -43729 29 -43723
rect -29 -49817 29 -49811
rect -29 -49851 -17 -49817
rect -29 -49857 29 -49851
rect -29 -49925 29 -49919
rect -29 -49959 -17 -49925
rect -29 -49965 29 -49959
rect -29 -56053 29 -56047
rect -29 -56087 -17 -56053
rect -29 -56093 29 -56087
rect -29 -56161 29 -56155
rect -29 -56195 -17 -56161
rect -29 -56201 29 -56195
rect -29 -62289 29 -62283
rect -29 -62323 -17 -62289
rect -29 -62329 29 -62323
<< nwell >>
rect -211 -62461 211 62461
<< pmos >>
rect -15 56242 15 62242
rect -15 50006 15 56006
rect -15 43770 15 49770
rect -15 37534 15 43534
rect -15 31298 15 37298
rect -15 25062 15 31062
rect -15 18826 15 24826
rect -15 12590 15 18590
rect -15 6354 15 12354
rect -15 118 15 6118
rect -15 -6118 15 -118
rect -15 -12354 15 -6354
rect -15 -18590 15 -12590
rect -15 -24826 15 -18826
rect -15 -31062 15 -25062
rect -15 -37298 15 -31298
rect -15 -43534 15 -37534
rect -15 -49770 15 -43770
rect -15 -56006 15 -50006
rect -15 -62242 15 -56242
<< pdiff >>
rect -73 62230 -15 62242
rect -73 56254 -61 62230
rect -27 56254 -15 62230
rect -73 56242 -15 56254
rect 15 62230 73 62242
rect 15 56254 27 62230
rect 61 56254 73 62230
rect 15 56242 73 56254
rect -73 55994 -15 56006
rect -73 50018 -61 55994
rect -27 50018 -15 55994
rect -73 50006 -15 50018
rect 15 55994 73 56006
rect 15 50018 27 55994
rect 61 50018 73 55994
rect 15 50006 73 50018
rect -73 49758 -15 49770
rect -73 43782 -61 49758
rect -27 43782 -15 49758
rect -73 43770 -15 43782
rect 15 49758 73 49770
rect 15 43782 27 49758
rect 61 43782 73 49758
rect 15 43770 73 43782
rect -73 43522 -15 43534
rect -73 37546 -61 43522
rect -27 37546 -15 43522
rect -73 37534 -15 37546
rect 15 43522 73 43534
rect 15 37546 27 43522
rect 61 37546 73 43522
rect 15 37534 73 37546
rect -73 37286 -15 37298
rect -73 31310 -61 37286
rect -27 31310 -15 37286
rect -73 31298 -15 31310
rect 15 37286 73 37298
rect 15 31310 27 37286
rect 61 31310 73 37286
rect 15 31298 73 31310
rect -73 31050 -15 31062
rect -73 25074 -61 31050
rect -27 25074 -15 31050
rect -73 25062 -15 25074
rect 15 31050 73 31062
rect 15 25074 27 31050
rect 61 25074 73 31050
rect 15 25062 73 25074
rect -73 24814 -15 24826
rect -73 18838 -61 24814
rect -27 18838 -15 24814
rect -73 18826 -15 18838
rect 15 24814 73 24826
rect 15 18838 27 24814
rect 61 18838 73 24814
rect 15 18826 73 18838
rect -73 18578 -15 18590
rect -73 12602 -61 18578
rect -27 12602 -15 18578
rect -73 12590 -15 12602
rect 15 18578 73 18590
rect 15 12602 27 18578
rect 61 12602 73 18578
rect 15 12590 73 12602
rect -73 12342 -15 12354
rect -73 6366 -61 12342
rect -27 6366 -15 12342
rect -73 6354 -15 6366
rect 15 12342 73 12354
rect 15 6366 27 12342
rect 61 6366 73 12342
rect 15 6354 73 6366
rect -73 6106 -15 6118
rect -73 130 -61 6106
rect -27 130 -15 6106
rect -73 118 -15 130
rect 15 6106 73 6118
rect 15 130 27 6106
rect 61 130 73 6106
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -6106 -61 -130
rect -27 -6106 -15 -130
rect -73 -6118 -15 -6106
rect 15 -130 73 -118
rect 15 -6106 27 -130
rect 61 -6106 73 -130
rect 15 -6118 73 -6106
rect -73 -6366 -15 -6354
rect -73 -12342 -61 -6366
rect -27 -12342 -15 -6366
rect -73 -12354 -15 -12342
rect 15 -6366 73 -6354
rect 15 -12342 27 -6366
rect 61 -12342 73 -6366
rect 15 -12354 73 -12342
rect -73 -12602 -15 -12590
rect -73 -18578 -61 -12602
rect -27 -18578 -15 -12602
rect -73 -18590 -15 -18578
rect 15 -12602 73 -12590
rect 15 -18578 27 -12602
rect 61 -18578 73 -12602
rect 15 -18590 73 -18578
rect -73 -18838 -15 -18826
rect -73 -24814 -61 -18838
rect -27 -24814 -15 -18838
rect -73 -24826 -15 -24814
rect 15 -18838 73 -18826
rect 15 -24814 27 -18838
rect 61 -24814 73 -18838
rect 15 -24826 73 -24814
rect -73 -25074 -15 -25062
rect -73 -31050 -61 -25074
rect -27 -31050 -15 -25074
rect -73 -31062 -15 -31050
rect 15 -25074 73 -25062
rect 15 -31050 27 -25074
rect 61 -31050 73 -25074
rect 15 -31062 73 -31050
rect -73 -31310 -15 -31298
rect -73 -37286 -61 -31310
rect -27 -37286 -15 -31310
rect -73 -37298 -15 -37286
rect 15 -31310 73 -31298
rect 15 -37286 27 -31310
rect 61 -37286 73 -31310
rect 15 -37298 73 -37286
rect -73 -37546 -15 -37534
rect -73 -43522 -61 -37546
rect -27 -43522 -15 -37546
rect -73 -43534 -15 -43522
rect 15 -37546 73 -37534
rect 15 -43522 27 -37546
rect 61 -43522 73 -37546
rect 15 -43534 73 -43522
rect -73 -43782 -15 -43770
rect -73 -49758 -61 -43782
rect -27 -49758 -15 -43782
rect -73 -49770 -15 -49758
rect 15 -43782 73 -43770
rect 15 -49758 27 -43782
rect 61 -49758 73 -43782
rect 15 -49770 73 -49758
rect -73 -50018 -15 -50006
rect -73 -55994 -61 -50018
rect -27 -55994 -15 -50018
rect -73 -56006 -15 -55994
rect 15 -50018 73 -50006
rect 15 -55994 27 -50018
rect 61 -55994 73 -50018
rect 15 -56006 73 -55994
rect -73 -56254 -15 -56242
rect -73 -62230 -61 -56254
rect -27 -62230 -15 -56254
rect -73 -62242 -15 -62230
rect 15 -56254 73 -56242
rect 15 -62230 27 -56254
rect 61 -62230 73 -56254
rect 15 -62242 73 -62230
<< pdiffc >>
rect -61 56254 -27 62230
rect 27 56254 61 62230
rect -61 50018 -27 55994
rect 27 50018 61 55994
rect -61 43782 -27 49758
rect 27 43782 61 49758
rect -61 37546 -27 43522
rect 27 37546 61 43522
rect -61 31310 -27 37286
rect 27 31310 61 37286
rect -61 25074 -27 31050
rect 27 25074 61 31050
rect -61 18838 -27 24814
rect 27 18838 61 24814
rect -61 12602 -27 18578
rect 27 12602 61 18578
rect -61 6366 -27 12342
rect 27 6366 61 12342
rect -61 130 -27 6106
rect 27 130 61 6106
rect -61 -6106 -27 -130
rect 27 -6106 61 -130
rect -61 -12342 -27 -6366
rect 27 -12342 61 -6366
rect -61 -18578 -27 -12602
rect 27 -18578 61 -12602
rect -61 -24814 -27 -18838
rect 27 -24814 61 -18838
rect -61 -31050 -27 -25074
rect 27 -31050 61 -25074
rect -61 -37286 -27 -31310
rect 27 -37286 61 -31310
rect -61 -43522 -27 -37546
rect 27 -43522 61 -37546
rect -61 -49758 -27 -43782
rect 27 -49758 61 -43782
rect -61 -55994 -27 -50018
rect 27 -55994 61 -50018
rect -61 -62230 -27 -56254
rect 27 -62230 61 -56254
<< nsubdiff >>
rect -175 62391 -79 62425
rect 79 62391 175 62425
rect -175 62329 -141 62391
rect 141 62329 175 62391
rect -175 -62391 -141 -62329
rect 141 -62391 175 -62329
rect -175 -62425 -79 -62391
rect 79 -62425 175 -62391
<< nsubdiffcont >>
rect -79 62391 79 62425
rect -175 -62329 -141 62329
rect 141 -62329 175 62329
rect -79 -62425 79 -62391
<< poly >>
rect -33 62323 33 62339
rect -33 62289 -17 62323
rect 17 62289 33 62323
rect -33 62273 33 62289
rect -15 62242 15 62273
rect -15 56211 15 56242
rect -33 56195 33 56211
rect -33 56161 -17 56195
rect 17 56161 33 56195
rect -33 56145 33 56161
rect -33 56087 33 56103
rect -33 56053 -17 56087
rect 17 56053 33 56087
rect -33 56037 33 56053
rect -15 56006 15 56037
rect -15 49975 15 50006
rect -33 49959 33 49975
rect -33 49925 -17 49959
rect 17 49925 33 49959
rect -33 49909 33 49925
rect -33 49851 33 49867
rect -33 49817 -17 49851
rect 17 49817 33 49851
rect -33 49801 33 49817
rect -15 49770 15 49801
rect -15 43739 15 43770
rect -33 43723 33 43739
rect -33 43689 -17 43723
rect 17 43689 33 43723
rect -33 43673 33 43689
rect -33 43615 33 43631
rect -33 43581 -17 43615
rect 17 43581 33 43615
rect -33 43565 33 43581
rect -15 43534 15 43565
rect -15 37503 15 37534
rect -33 37487 33 37503
rect -33 37453 -17 37487
rect 17 37453 33 37487
rect -33 37437 33 37453
rect -33 37379 33 37395
rect -33 37345 -17 37379
rect 17 37345 33 37379
rect -33 37329 33 37345
rect -15 37298 15 37329
rect -15 31267 15 31298
rect -33 31251 33 31267
rect -33 31217 -17 31251
rect 17 31217 33 31251
rect -33 31201 33 31217
rect -33 31143 33 31159
rect -33 31109 -17 31143
rect 17 31109 33 31143
rect -33 31093 33 31109
rect -15 31062 15 31093
rect -15 25031 15 25062
rect -33 25015 33 25031
rect -33 24981 -17 25015
rect 17 24981 33 25015
rect -33 24965 33 24981
rect -33 24907 33 24923
rect -33 24873 -17 24907
rect 17 24873 33 24907
rect -33 24857 33 24873
rect -15 24826 15 24857
rect -15 18795 15 18826
rect -33 18779 33 18795
rect -33 18745 -17 18779
rect 17 18745 33 18779
rect -33 18729 33 18745
rect -33 18671 33 18687
rect -33 18637 -17 18671
rect 17 18637 33 18671
rect -33 18621 33 18637
rect -15 18590 15 18621
rect -15 12559 15 12590
rect -33 12543 33 12559
rect -33 12509 -17 12543
rect 17 12509 33 12543
rect -33 12493 33 12509
rect -33 12435 33 12451
rect -33 12401 -17 12435
rect 17 12401 33 12435
rect -33 12385 33 12401
rect -15 12354 15 12385
rect -15 6323 15 6354
rect -33 6307 33 6323
rect -33 6273 -17 6307
rect 17 6273 33 6307
rect -33 6257 33 6273
rect -33 6199 33 6215
rect -33 6165 -17 6199
rect 17 6165 33 6199
rect -33 6149 33 6165
rect -15 6118 15 6149
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -6149 15 -6118
rect -33 -6165 33 -6149
rect -33 -6199 -17 -6165
rect 17 -6199 33 -6165
rect -33 -6215 33 -6199
rect -33 -6273 33 -6257
rect -33 -6307 -17 -6273
rect 17 -6307 33 -6273
rect -33 -6323 33 -6307
rect -15 -6354 15 -6323
rect -15 -12385 15 -12354
rect -33 -12401 33 -12385
rect -33 -12435 -17 -12401
rect 17 -12435 33 -12401
rect -33 -12451 33 -12435
rect -33 -12509 33 -12493
rect -33 -12543 -17 -12509
rect 17 -12543 33 -12509
rect -33 -12559 33 -12543
rect -15 -12590 15 -12559
rect -15 -18621 15 -18590
rect -33 -18637 33 -18621
rect -33 -18671 -17 -18637
rect 17 -18671 33 -18637
rect -33 -18687 33 -18671
rect -33 -18745 33 -18729
rect -33 -18779 -17 -18745
rect 17 -18779 33 -18745
rect -33 -18795 33 -18779
rect -15 -18826 15 -18795
rect -15 -24857 15 -24826
rect -33 -24873 33 -24857
rect -33 -24907 -17 -24873
rect 17 -24907 33 -24873
rect -33 -24923 33 -24907
rect -33 -24981 33 -24965
rect -33 -25015 -17 -24981
rect 17 -25015 33 -24981
rect -33 -25031 33 -25015
rect -15 -25062 15 -25031
rect -15 -31093 15 -31062
rect -33 -31109 33 -31093
rect -33 -31143 -17 -31109
rect 17 -31143 33 -31109
rect -33 -31159 33 -31143
rect -33 -31217 33 -31201
rect -33 -31251 -17 -31217
rect 17 -31251 33 -31217
rect -33 -31267 33 -31251
rect -15 -31298 15 -31267
rect -15 -37329 15 -37298
rect -33 -37345 33 -37329
rect -33 -37379 -17 -37345
rect 17 -37379 33 -37345
rect -33 -37395 33 -37379
rect -33 -37453 33 -37437
rect -33 -37487 -17 -37453
rect 17 -37487 33 -37453
rect -33 -37503 33 -37487
rect -15 -37534 15 -37503
rect -15 -43565 15 -43534
rect -33 -43581 33 -43565
rect -33 -43615 -17 -43581
rect 17 -43615 33 -43581
rect -33 -43631 33 -43615
rect -33 -43689 33 -43673
rect -33 -43723 -17 -43689
rect 17 -43723 33 -43689
rect -33 -43739 33 -43723
rect -15 -43770 15 -43739
rect -15 -49801 15 -49770
rect -33 -49817 33 -49801
rect -33 -49851 -17 -49817
rect 17 -49851 33 -49817
rect -33 -49867 33 -49851
rect -33 -49925 33 -49909
rect -33 -49959 -17 -49925
rect 17 -49959 33 -49925
rect -33 -49975 33 -49959
rect -15 -50006 15 -49975
rect -15 -56037 15 -56006
rect -33 -56053 33 -56037
rect -33 -56087 -17 -56053
rect 17 -56087 33 -56053
rect -33 -56103 33 -56087
rect -33 -56161 33 -56145
rect -33 -56195 -17 -56161
rect 17 -56195 33 -56161
rect -33 -56211 33 -56195
rect -15 -56242 15 -56211
rect -15 -62273 15 -62242
rect -33 -62289 33 -62273
rect -33 -62323 -17 -62289
rect 17 -62323 33 -62289
rect -33 -62339 33 -62323
<< polycont >>
rect -17 62289 17 62323
rect -17 56161 17 56195
rect -17 56053 17 56087
rect -17 49925 17 49959
rect -17 49817 17 49851
rect -17 43689 17 43723
rect -17 43581 17 43615
rect -17 37453 17 37487
rect -17 37345 17 37379
rect -17 31217 17 31251
rect -17 31109 17 31143
rect -17 24981 17 25015
rect -17 24873 17 24907
rect -17 18745 17 18779
rect -17 18637 17 18671
rect -17 12509 17 12543
rect -17 12401 17 12435
rect -17 6273 17 6307
rect -17 6165 17 6199
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -6199 17 -6165
rect -17 -6307 17 -6273
rect -17 -12435 17 -12401
rect -17 -12543 17 -12509
rect -17 -18671 17 -18637
rect -17 -18779 17 -18745
rect -17 -24907 17 -24873
rect -17 -25015 17 -24981
rect -17 -31143 17 -31109
rect -17 -31251 17 -31217
rect -17 -37379 17 -37345
rect -17 -37487 17 -37453
rect -17 -43615 17 -43581
rect -17 -43723 17 -43689
rect -17 -49851 17 -49817
rect -17 -49959 17 -49925
rect -17 -56087 17 -56053
rect -17 -56195 17 -56161
rect -17 -62323 17 -62289
<< locali >>
rect -175 62391 -79 62425
rect 79 62391 175 62425
rect -175 62329 -141 62391
rect 141 62329 175 62391
rect -33 62289 -17 62323
rect 17 62289 33 62323
rect -61 62230 -27 62246
rect -61 56238 -27 56254
rect 27 62230 61 62246
rect 27 56238 61 56254
rect -33 56161 -17 56195
rect 17 56161 33 56195
rect -33 56053 -17 56087
rect 17 56053 33 56087
rect -61 55994 -27 56010
rect -61 50002 -27 50018
rect 27 55994 61 56010
rect 27 50002 61 50018
rect -33 49925 -17 49959
rect 17 49925 33 49959
rect -33 49817 -17 49851
rect 17 49817 33 49851
rect -61 49758 -27 49774
rect -61 43766 -27 43782
rect 27 49758 61 49774
rect 27 43766 61 43782
rect -33 43689 -17 43723
rect 17 43689 33 43723
rect -33 43581 -17 43615
rect 17 43581 33 43615
rect -61 43522 -27 43538
rect -61 37530 -27 37546
rect 27 43522 61 43538
rect 27 37530 61 37546
rect -33 37453 -17 37487
rect 17 37453 33 37487
rect -33 37345 -17 37379
rect 17 37345 33 37379
rect -61 37286 -27 37302
rect -61 31294 -27 31310
rect 27 37286 61 37302
rect 27 31294 61 31310
rect -33 31217 -17 31251
rect 17 31217 33 31251
rect -33 31109 -17 31143
rect 17 31109 33 31143
rect -61 31050 -27 31066
rect -61 25058 -27 25074
rect 27 31050 61 31066
rect 27 25058 61 25074
rect -33 24981 -17 25015
rect 17 24981 33 25015
rect -33 24873 -17 24907
rect 17 24873 33 24907
rect -61 24814 -27 24830
rect -61 18822 -27 18838
rect 27 24814 61 24830
rect 27 18822 61 18838
rect -33 18745 -17 18779
rect 17 18745 33 18779
rect -33 18637 -17 18671
rect 17 18637 33 18671
rect -61 18578 -27 18594
rect -61 12586 -27 12602
rect 27 18578 61 18594
rect 27 12586 61 12602
rect -33 12509 -17 12543
rect 17 12509 33 12543
rect -33 12401 -17 12435
rect 17 12401 33 12435
rect -61 12342 -27 12358
rect -61 6350 -27 6366
rect 27 12342 61 12358
rect 27 6350 61 6366
rect -33 6273 -17 6307
rect 17 6273 33 6307
rect -33 6165 -17 6199
rect 17 6165 33 6199
rect -61 6106 -27 6122
rect -61 114 -27 130
rect 27 6106 61 6122
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -6122 -27 -6106
rect 27 -130 61 -114
rect 27 -6122 61 -6106
rect -33 -6199 -17 -6165
rect 17 -6199 33 -6165
rect -33 -6307 -17 -6273
rect 17 -6307 33 -6273
rect -61 -6366 -27 -6350
rect -61 -12358 -27 -12342
rect 27 -6366 61 -6350
rect 27 -12358 61 -12342
rect -33 -12435 -17 -12401
rect 17 -12435 33 -12401
rect -33 -12543 -17 -12509
rect 17 -12543 33 -12509
rect -61 -12602 -27 -12586
rect -61 -18594 -27 -18578
rect 27 -12602 61 -12586
rect 27 -18594 61 -18578
rect -33 -18671 -17 -18637
rect 17 -18671 33 -18637
rect -33 -18779 -17 -18745
rect 17 -18779 33 -18745
rect -61 -18838 -27 -18822
rect -61 -24830 -27 -24814
rect 27 -18838 61 -18822
rect 27 -24830 61 -24814
rect -33 -24907 -17 -24873
rect 17 -24907 33 -24873
rect -33 -25015 -17 -24981
rect 17 -25015 33 -24981
rect -61 -25074 -27 -25058
rect -61 -31066 -27 -31050
rect 27 -25074 61 -25058
rect 27 -31066 61 -31050
rect -33 -31143 -17 -31109
rect 17 -31143 33 -31109
rect -33 -31251 -17 -31217
rect 17 -31251 33 -31217
rect -61 -31310 -27 -31294
rect -61 -37302 -27 -37286
rect 27 -31310 61 -31294
rect 27 -37302 61 -37286
rect -33 -37379 -17 -37345
rect 17 -37379 33 -37345
rect -33 -37487 -17 -37453
rect 17 -37487 33 -37453
rect -61 -37546 -27 -37530
rect -61 -43538 -27 -43522
rect 27 -37546 61 -37530
rect 27 -43538 61 -43522
rect -33 -43615 -17 -43581
rect 17 -43615 33 -43581
rect -33 -43723 -17 -43689
rect 17 -43723 33 -43689
rect -61 -43782 -27 -43766
rect -61 -49774 -27 -49758
rect 27 -43782 61 -43766
rect 27 -49774 61 -49758
rect -33 -49851 -17 -49817
rect 17 -49851 33 -49817
rect -33 -49959 -17 -49925
rect 17 -49959 33 -49925
rect -61 -50018 -27 -50002
rect -61 -56010 -27 -55994
rect 27 -50018 61 -50002
rect 27 -56010 61 -55994
rect -33 -56087 -17 -56053
rect 17 -56087 33 -56053
rect -33 -56195 -17 -56161
rect 17 -56195 33 -56161
rect -61 -56254 -27 -56238
rect -61 -62246 -27 -62230
rect 27 -56254 61 -56238
rect 27 -62246 61 -62230
rect -33 -62323 -17 -62289
rect 17 -62323 33 -62289
rect -175 -62391 -141 -62329
rect 141 -62391 175 -62329
rect -175 -62425 -79 -62391
rect 79 -62425 175 -62391
<< viali >>
rect -17 62289 17 62323
rect -61 56254 -27 62230
rect 27 56254 61 62230
rect -17 56161 17 56195
rect -17 56053 17 56087
rect -61 50018 -27 55994
rect 27 50018 61 55994
rect -17 49925 17 49959
rect -17 49817 17 49851
rect -61 43782 -27 49758
rect 27 43782 61 49758
rect -17 43689 17 43723
rect -17 43581 17 43615
rect -61 37546 -27 43522
rect 27 37546 61 43522
rect -17 37453 17 37487
rect -17 37345 17 37379
rect -61 31310 -27 37286
rect 27 31310 61 37286
rect -17 31217 17 31251
rect -17 31109 17 31143
rect -61 25074 -27 31050
rect 27 25074 61 31050
rect -17 24981 17 25015
rect -17 24873 17 24907
rect -61 18838 -27 24814
rect 27 18838 61 24814
rect -17 18745 17 18779
rect -17 18637 17 18671
rect -61 12602 -27 18578
rect 27 12602 61 18578
rect -17 12509 17 12543
rect -17 12401 17 12435
rect -61 6366 -27 12342
rect 27 6366 61 12342
rect -17 6273 17 6307
rect -17 6165 17 6199
rect -61 130 -27 6106
rect 27 130 61 6106
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -6106 -27 -130
rect 27 -6106 61 -130
rect -17 -6199 17 -6165
rect -17 -6307 17 -6273
rect -61 -12342 -27 -6366
rect 27 -12342 61 -6366
rect -17 -12435 17 -12401
rect -17 -12543 17 -12509
rect -61 -18578 -27 -12602
rect 27 -18578 61 -12602
rect -17 -18671 17 -18637
rect -17 -18779 17 -18745
rect -61 -24814 -27 -18838
rect 27 -24814 61 -18838
rect -17 -24907 17 -24873
rect -17 -25015 17 -24981
rect -61 -31050 -27 -25074
rect 27 -31050 61 -25074
rect -17 -31143 17 -31109
rect -17 -31251 17 -31217
rect -61 -37286 -27 -31310
rect 27 -37286 61 -31310
rect -17 -37379 17 -37345
rect -17 -37487 17 -37453
rect -61 -43522 -27 -37546
rect 27 -43522 61 -37546
rect -17 -43615 17 -43581
rect -17 -43723 17 -43689
rect -61 -49758 -27 -43782
rect 27 -49758 61 -43782
rect -17 -49851 17 -49817
rect -17 -49959 17 -49925
rect -61 -55994 -27 -50018
rect 27 -55994 61 -50018
rect -17 -56087 17 -56053
rect -17 -56195 17 -56161
rect -61 -62230 -27 -56254
rect 27 -62230 61 -56254
rect -17 -62323 17 -62289
<< metal1 >>
rect -29 62323 29 62329
rect -29 62289 -17 62323
rect 17 62289 29 62323
rect -29 62283 29 62289
rect -67 62230 -21 62242
rect -67 56254 -61 62230
rect -27 56254 -21 62230
rect -67 56242 -21 56254
rect 21 62230 67 62242
rect 21 56254 27 62230
rect 61 56254 67 62230
rect 21 56242 67 56254
rect -29 56195 29 56201
rect -29 56161 -17 56195
rect 17 56161 29 56195
rect -29 56155 29 56161
rect -29 56087 29 56093
rect -29 56053 -17 56087
rect 17 56053 29 56087
rect -29 56047 29 56053
rect -67 55994 -21 56006
rect -67 50018 -61 55994
rect -27 50018 -21 55994
rect -67 50006 -21 50018
rect 21 55994 67 56006
rect 21 50018 27 55994
rect 61 50018 67 55994
rect 21 50006 67 50018
rect -29 49959 29 49965
rect -29 49925 -17 49959
rect 17 49925 29 49959
rect -29 49919 29 49925
rect -29 49851 29 49857
rect -29 49817 -17 49851
rect 17 49817 29 49851
rect -29 49811 29 49817
rect -67 49758 -21 49770
rect -67 43782 -61 49758
rect -27 43782 -21 49758
rect -67 43770 -21 43782
rect 21 49758 67 49770
rect 21 43782 27 49758
rect 61 43782 67 49758
rect 21 43770 67 43782
rect -29 43723 29 43729
rect -29 43689 -17 43723
rect 17 43689 29 43723
rect -29 43683 29 43689
rect -29 43615 29 43621
rect -29 43581 -17 43615
rect 17 43581 29 43615
rect -29 43575 29 43581
rect -67 43522 -21 43534
rect -67 37546 -61 43522
rect -27 37546 -21 43522
rect -67 37534 -21 37546
rect 21 43522 67 43534
rect 21 37546 27 43522
rect 61 37546 67 43522
rect 21 37534 67 37546
rect -29 37487 29 37493
rect -29 37453 -17 37487
rect 17 37453 29 37487
rect -29 37447 29 37453
rect -29 37379 29 37385
rect -29 37345 -17 37379
rect 17 37345 29 37379
rect -29 37339 29 37345
rect -67 37286 -21 37298
rect -67 31310 -61 37286
rect -27 31310 -21 37286
rect -67 31298 -21 31310
rect 21 37286 67 37298
rect 21 31310 27 37286
rect 61 31310 67 37286
rect 21 31298 67 31310
rect -29 31251 29 31257
rect -29 31217 -17 31251
rect 17 31217 29 31251
rect -29 31211 29 31217
rect -29 31143 29 31149
rect -29 31109 -17 31143
rect 17 31109 29 31143
rect -29 31103 29 31109
rect -67 31050 -21 31062
rect -67 25074 -61 31050
rect -27 25074 -21 31050
rect -67 25062 -21 25074
rect 21 31050 67 31062
rect 21 25074 27 31050
rect 61 25074 67 31050
rect 21 25062 67 25074
rect -29 25015 29 25021
rect -29 24981 -17 25015
rect 17 24981 29 25015
rect -29 24975 29 24981
rect -29 24907 29 24913
rect -29 24873 -17 24907
rect 17 24873 29 24907
rect -29 24867 29 24873
rect -67 24814 -21 24826
rect -67 18838 -61 24814
rect -27 18838 -21 24814
rect -67 18826 -21 18838
rect 21 24814 67 24826
rect 21 18838 27 24814
rect 61 18838 67 24814
rect 21 18826 67 18838
rect -29 18779 29 18785
rect -29 18745 -17 18779
rect 17 18745 29 18779
rect -29 18739 29 18745
rect -29 18671 29 18677
rect -29 18637 -17 18671
rect 17 18637 29 18671
rect -29 18631 29 18637
rect -67 18578 -21 18590
rect -67 12602 -61 18578
rect -27 12602 -21 18578
rect -67 12590 -21 12602
rect 21 18578 67 18590
rect 21 12602 27 18578
rect 61 12602 67 18578
rect 21 12590 67 12602
rect -29 12543 29 12549
rect -29 12509 -17 12543
rect 17 12509 29 12543
rect -29 12503 29 12509
rect -29 12435 29 12441
rect -29 12401 -17 12435
rect 17 12401 29 12435
rect -29 12395 29 12401
rect -67 12342 -21 12354
rect -67 6366 -61 12342
rect -27 6366 -21 12342
rect -67 6354 -21 6366
rect 21 12342 67 12354
rect 21 6366 27 12342
rect 61 6366 67 12342
rect 21 6354 67 6366
rect -29 6307 29 6313
rect -29 6273 -17 6307
rect 17 6273 29 6307
rect -29 6267 29 6273
rect -29 6199 29 6205
rect -29 6165 -17 6199
rect 17 6165 29 6199
rect -29 6159 29 6165
rect -67 6106 -21 6118
rect -67 130 -61 6106
rect -27 130 -21 6106
rect -67 118 -21 130
rect 21 6106 67 6118
rect 21 130 27 6106
rect 61 130 67 6106
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -6106 -61 -130
rect -27 -6106 -21 -130
rect -67 -6118 -21 -6106
rect 21 -130 67 -118
rect 21 -6106 27 -130
rect 61 -6106 67 -130
rect 21 -6118 67 -6106
rect -29 -6165 29 -6159
rect -29 -6199 -17 -6165
rect 17 -6199 29 -6165
rect -29 -6205 29 -6199
rect -29 -6273 29 -6267
rect -29 -6307 -17 -6273
rect 17 -6307 29 -6273
rect -29 -6313 29 -6307
rect -67 -6366 -21 -6354
rect -67 -12342 -61 -6366
rect -27 -12342 -21 -6366
rect -67 -12354 -21 -12342
rect 21 -6366 67 -6354
rect 21 -12342 27 -6366
rect 61 -12342 67 -6366
rect 21 -12354 67 -12342
rect -29 -12401 29 -12395
rect -29 -12435 -17 -12401
rect 17 -12435 29 -12401
rect -29 -12441 29 -12435
rect -29 -12509 29 -12503
rect -29 -12543 -17 -12509
rect 17 -12543 29 -12509
rect -29 -12549 29 -12543
rect -67 -12602 -21 -12590
rect -67 -18578 -61 -12602
rect -27 -18578 -21 -12602
rect -67 -18590 -21 -18578
rect 21 -12602 67 -12590
rect 21 -18578 27 -12602
rect 61 -18578 67 -12602
rect 21 -18590 67 -18578
rect -29 -18637 29 -18631
rect -29 -18671 -17 -18637
rect 17 -18671 29 -18637
rect -29 -18677 29 -18671
rect -29 -18745 29 -18739
rect -29 -18779 -17 -18745
rect 17 -18779 29 -18745
rect -29 -18785 29 -18779
rect -67 -18838 -21 -18826
rect -67 -24814 -61 -18838
rect -27 -24814 -21 -18838
rect -67 -24826 -21 -24814
rect 21 -18838 67 -18826
rect 21 -24814 27 -18838
rect 61 -24814 67 -18838
rect 21 -24826 67 -24814
rect -29 -24873 29 -24867
rect -29 -24907 -17 -24873
rect 17 -24907 29 -24873
rect -29 -24913 29 -24907
rect -29 -24981 29 -24975
rect -29 -25015 -17 -24981
rect 17 -25015 29 -24981
rect -29 -25021 29 -25015
rect -67 -25074 -21 -25062
rect -67 -31050 -61 -25074
rect -27 -31050 -21 -25074
rect -67 -31062 -21 -31050
rect 21 -25074 67 -25062
rect 21 -31050 27 -25074
rect 61 -31050 67 -25074
rect 21 -31062 67 -31050
rect -29 -31109 29 -31103
rect -29 -31143 -17 -31109
rect 17 -31143 29 -31109
rect -29 -31149 29 -31143
rect -29 -31217 29 -31211
rect -29 -31251 -17 -31217
rect 17 -31251 29 -31217
rect -29 -31257 29 -31251
rect -67 -31310 -21 -31298
rect -67 -37286 -61 -31310
rect -27 -37286 -21 -31310
rect -67 -37298 -21 -37286
rect 21 -31310 67 -31298
rect 21 -37286 27 -31310
rect 61 -37286 67 -31310
rect 21 -37298 67 -37286
rect -29 -37345 29 -37339
rect -29 -37379 -17 -37345
rect 17 -37379 29 -37345
rect -29 -37385 29 -37379
rect -29 -37453 29 -37447
rect -29 -37487 -17 -37453
rect 17 -37487 29 -37453
rect -29 -37493 29 -37487
rect -67 -37546 -21 -37534
rect -67 -43522 -61 -37546
rect -27 -43522 -21 -37546
rect -67 -43534 -21 -43522
rect 21 -37546 67 -37534
rect 21 -43522 27 -37546
rect 61 -43522 67 -37546
rect 21 -43534 67 -43522
rect -29 -43581 29 -43575
rect -29 -43615 -17 -43581
rect 17 -43615 29 -43581
rect -29 -43621 29 -43615
rect -29 -43689 29 -43683
rect -29 -43723 -17 -43689
rect 17 -43723 29 -43689
rect -29 -43729 29 -43723
rect -67 -43782 -21 -43770
rect -67 -49758 -61 -43782
rect -27 -49758 -21 -43782
rect -67 -49770 -21 -49758
rect 21 -43782 67 -43770
rect 21 -49758 27 -43782
rect 61 -49758 67 -43782
rect 21 -49770 67 -49758
rect -29 -49817 29 -49811
rect -29 -49851 -17 -49817
rect 17 -49851 29 -49817
rect -29 -49857 29 -49851
rect -29 -49925 29 -49919
rect -29 -49959 -17 -49925
rect 17 -49959 29 -49925
rect -29 -49965 29 -49959
rect -67 -50018 -21 -50006
rect -67 -55994 -61 -50018
rect -27 -55994 -21 -50018
rect -67 -56006 -21 -55994
rect 21 -50018 67 -50006
rect 21 -55994 27 -50018
rect 61 -55994 67 -50018
rect 21 -56006 67 -55994
rect -29 -56053 29 -56047
rect -29 -56087 -17 -56053
rect 17 -56087 29 -56053
rect -29 -56093 29 -56087
rect -29 -56161 29 -56155
rect -29 -56195 -17 -56161
rect 17 -56195 29 -56161
rect -29 -56201 29 -56195
rect -67 -56254 -21 -56242
rect -67 -62230 -61 -56254
rect -27 -62230 -21 -56254
rect -67 -62242 -21 -62230
rect 21 -56254 67 -56242
rect 21 -62230 27 -56254
rect 61 -62230 67 -56254
rect 21 -62242 67 -62230
rect -29 -62289 29 -62283
rect -29 -62323 -17 -62289
rect 17 -62323 29 -62289
rect -29 -62329 29 -62323
<< labels >>
rlabel nsubdiffcont 0 -62408 0 -62408 0 B
port 1 nsew
rlabel pdiffc -44 -59242 -44 -59242 0 D0
port 2 nsew
rlabel pdiffc 44 -59242 44 -59242 0 S0
port 3 nsew
rlabel polycont 0 -56178 0 -56178 0 G0
port 4 nsew
rlabel pdiffc -44 -53006 -44 -53006 0 D1
port 5 nsew
rlabel pdiffc 44 -53006 44 -53006 0 S1
port 6 nsew
rlabel polycont 0 -49942 0 -49942 0 G1
port 7 nsew
rlabel pdiffc -44 -46770 -44 -46770 0 D2
port 8 nsew
rlabel pdiffc 44 -46770 44 -46770 0 S2
port 9 nsew
rlabel polycont 0 -43706 0 -43706 0 G2
port 10 nsew
rlabel pdiffc -44 -40534 -44 -40534 0 D3
port 11 nsew
rlabel pdiffc 44 -40534 44 -40534 0 S3
port 12 nsew
rlabel polycont 0 -37470 0 -37470 0 G3
port 13 nsew
rlabel pdiffc -44 -34298 -44 -34298 0 D4
port 14 nsew
rlabel pdiffc 44 -34298 44 -34298 0 S4
port 15 nsew
rlabel polycont 0 -31234 0 -31234 0 G4
port 16 nsew
rlabel pdiffc -44 -28062 -44 -28062 0 D5
port 17 nsew
rlabel pdiffc 44 -28062 44 -28062 0 S5
port 18 nsew
rlabel polycont 0 -24998 0 -24998 0 G5
port 19 nsew
rlabel pdiffc -44 -21826 -44 -21826 0 D6
port 20 nsew
rlabel pdiffc 44 -21826 44 -21826 0 S6
port 21 nsew
rlabel polycont 0 -18762 0 -18762 0 G6
port 22 nsew
rlabel pdiffc -44 -15590 -44 -15590 0 D7
port 23 nsew
rlabel pdiffc 44 -15590 44 -15590 0 S7
port 24 nsew
rlabel polycont 0 -12526 0 -12526 0 G7
port 25 nsew
rlabel pdiffc -44 -9354 -44 -9354 0 D8
port 26 nsew
rlabel pdiffc 44 -9354 44 -9354 0 S8
port 27 nsew
rlabel polycont 0 -6290 0 -6290 0 G8
port 28 nsew
rlabel pdiffc -44 -3118 -44 -3118 0 D9
port 29 nsew
rlabel pdiffc 44 -3118 44 -3118 0 S9
port 30 nsew
rlabel polycont 0 -54 0 -54 0 G9
port 31 nsew
rlabel pdiffc -44 3118 -44 3118 0 D10
port 32 nsew
rlabel pdiffc 44 3118 44 3118 0 S10
port 33 nsew
rlabel polycont 0 6182 0 6182 0 G10
port 34 nsew
rlabel pdiffc -44 9354 -44 9354 0 D11
port 35 nsew
rlabel pdiffc 44 9354 44 9354 0 S11
port 36 nsew
rlabel polycont 0 12418 0 12418 0 G11
port 37 nsew
rlabel pdiffc -44 15590 -44 15590 0 D12
port 38 nsew
rlabel pdiffc 44 15590 44 15590 0 S12
port 39 nsew
rlabel polycont 0 18654 0 18654 0 G12
port 40 nsew
rlabel pdiffc -44 21826 -44 21826 0 D13
port 41 nsew
rlabel pdiffc 44 21826 44 21826 0 S13
port 42 nsew
rlabel polycont 0 24890 0 24890 0 G13
port 43 nsew
rlabel pdiffc -44 28062 -44 28062 0 D14
port 44 nsew
rlabel pdiffc 44 28062 44 28062 0 S14
port 45 nsew
rlabel polycont 0 31126 0 31126 0 G14
port 46 nsew
rlabel pdiffc -44 34298 -44 34298 0 D15
port 47 nsew
rlabel pdiffc 44 34298 44 34298 0 S15
port 48 nsew
rlabel polycont 0 37362 0 37362 0 G15
port 49 nsew
rlabel pdiffc -44 40534 -44 40534 0 D16
port 50 nsew
rlabel pdiffc 44 40534 44 40534 0 S16
port 51 nsew
rlabel polycont 0 43598 0 43598 0 G16
port 52 nsew
rlabel pdiffc -44 46770 -44 46770 0 D17
port 53 nsew
rlabel pdiffc 44 46770 44 46770 0 S17
port 54 nsew
rlabel polycont 0 49834 0 49834 0 G17
port 55 nsew
rlabel pdiffc -44 53006 -44 53006 0 D18
port 56 nsew
rlabel pdiffc 44 53006 44 53006 0 S18
port 57 nsew
rlabel polycont 0 56070 0 56070 0 G18
port 58 nsew
rlabel pdiffc -44 59242 -44 59242 0 D19
port 59 nsew
rlabel pdiffc 44 59242 44 59242 0 S19
port 60 nsew
rlabel polycont 0 62306 0 62306 0 G19
port 61 nsew
<< properties >>
string FIXED_BBOX -158 -62408 158 62408
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 30.0 l 0.15 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1 ad 8.7 as 8.7 pd 60.58 ps 60.58 nrd 0.00966666666666667 nrs 0.00966666666666667 sa 0 sb 0 sd 0 mult 20
<< end >>
