* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff = -0.010
* Number of bins: 49
.param
+ sky130_fd_pr__nfet_g5v0d10v5__toxe_mult = 1.0
+ sky130_fd_pr__nfet_g5v0d10v5__rshn_mult = 1.0
+ sky130_fd_pr__nfet_g5v0d10v5__overlap_mult = 0.89805
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = 9.9505e-1
+ sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult = 1.0144e+0
+ sky130_fd_pr__nfet_g5v0d10v5__lint_diff = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__wint_diff = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__dlc_diff = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__dwc_diff = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 000, W = 10.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0 = -0.0040673
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0 = 0.004518
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0 = ' -0.029667 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0 = -4.0229e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0 = -3454.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0 = 0.20809
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0 = 8.9403e-19
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 001, W = 15.0, L = 1.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1 = 0.0041381
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1 = 0.00081984
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1 = ' -0.027418 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1 = -0.0019156
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1 = -4.0807e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1 = -0.0021526
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1 = 0.28834
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1 = -1.9191e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 002, W = 15.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2 = 0.19886
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2 = 9.4919e-19
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2 = -0.004621
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2 = 0.0057526
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2 = ' -0.019002 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2 = -3.3871e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2 = -240.09
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 003, W = 1.5, L = 1.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3 = 0.40503
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3 = -1.1047e-19
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3 = -0.003457
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3 = -0.0018906
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3 = ' -0.047528 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3 = -0.0025502
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3 = 2.07e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3 = -0.0029411
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 004, W = 1.5, L = 2.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4 = -0.0069981
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4 = 0.40977
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4 = -7.7364e-20
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4 = -0.012669
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4 = -0.0013003
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4 = ' -0.036138 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4 = 0.016072
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4 = 1.3854e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 005, W = 1.5, L = 4.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5 = 1.5709e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5 = -0.0027239
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5 = 1.4396e-20
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5 = 0.44344
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5 = -0.016401
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5 = -0.00065178
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5 = ' -0.022464 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5 = 0.0092656
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 006, W = 1.5, L = 0.5
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6 = 4.4758e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6 = -5802.9
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6 = 4.799e-19
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6 = 0.46614
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6 = 0.0026935
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6 = 0.00056839
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6 = ' -0.047902 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 007, W = 1.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7 = 0.0024141
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7 = 7.1734e-13
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7 = -0.0071612
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7 = 2.3936e-19
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7 = 0.44078
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7 = 0.0066427
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7 = 6.4698e-5
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7 = ' -0.037156 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 008, W = 1.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8 = 0.0017771
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8 = 2.7032e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8 = -0.0034746
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8 = 1.6905e-19
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8 = 0.45085
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8 = -0.016086
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8 = -0.00022984
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8 = ' -0.031099 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 009, W = 1.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9 = -6.9939e-5
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9 = 0.0095036
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9 = 2.3937e-12
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9 = -0.0033641
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9 = 2.0697e-19
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9 = 0.475
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9 = -0.0097819
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9 = ' -0.023728 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 010, W = 1.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10 = -0.00043688
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10 = -0.00030286
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10 = -0.0012863
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10 = ' -0.025384 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10 = -0.011768
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10 = 0.54261
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10 = 1.3166e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10 = 1.0118e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 011, W = 1.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11 = 9.1925e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11 = 0.00050158
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11 = -5029.3
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11 = ' -0.029992 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11 = 0.0057524
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11 = 0.50711
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11 = 1.0295e-11
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 012, W = 1.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12 = 0.45674
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12 = 5.6764e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12 = 6.4202e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12 = 0.00099605
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12 = -5703.7
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12 = ' -0.038872 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12 = -0.00058493
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 013, W = 1.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13 = -0.0040079
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13 = 0.45136
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13 = 5.7016e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13 = 3.3811e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13 = -0.00056411
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13 = -4336.2
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13 = ' -0.018352 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 014, W = 20.0, L = 1.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14 = ' -0.023854 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14 = 0.0038916
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14 = 0.28785
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14 = -1.3826e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14 = -1.5094e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14 = -0.024639
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14 = 0.001071
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14 = 0.04329
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 015, W = 20.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15 = ' -0.018147 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15 = -0.0050434
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15 = 0.16952
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15 = 2.1478e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15 = 1.1465e-18
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15 = 0.0042157
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15 = -2329.7
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 016, W = 3.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16 = ' -0.030154 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16 = -0.0054809
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16 = 0.33488
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16 = 2.0355e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16 = -7.105e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16 = -0.0049461
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16 = -0.0010575
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16 = 0.0069932
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 017, W = 3.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17 = 0.0030754
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17 = ' -0.029897 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17 = -0.013966
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17 = 0.35229
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17 = 1.2012e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17 = -6.5305e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17 = -0.0035995
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17 = -0.00070267
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 018, W = 3.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18 = -0.00091243
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18 = 0.015143
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18 = ' -0.027618 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18 = -0.018565
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18 = 0.39546
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18 = 1.8827e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18 = -4.0537e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18 = -0.0053012
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 019, W = 3.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19 = -0.00099573
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19 = 0.0034779
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19 = ' -0.030559 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19 = -0.02028
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19 = 0.44945
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19 = 1.8294e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19 = -5.1199e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19 = -0.0029181
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 020, W = 3.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20 = 0.0020465
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20 = -2130.8
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20 = ' -0.027277 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20 = -0.0011535
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20 = 0.32846
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20 = 2.9889e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20 = 6.9218e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 021, W = 3.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21 = 0.0012316
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21 = -3422.1
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21 = ' -0.018699 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21 = -0.0042518
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21 = 0.29677
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21 = 3.0882e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21 = 5.1269e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 022, W = 5.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22 = -3.4186e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22 = -0.01089
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22 = 4.7233e-5
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22 = 0.021221
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22 = ' -0.033499 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22 = 0.0050875
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22 = 0.3001
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22 = -5.02e-14
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 023, W = 5.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23 = 0.34333
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23 = 2.4666e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23 = -1.8273e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23 = -0.0082333
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23 = -0.0016627
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23 = 0.022524
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23 = ' -0.032779 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23 = -0.004773
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 024, W = 5.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24 = -0.0091071
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24 = 0.38706
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24 = 2.7814e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24 = -2.6555e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24 = -0.0060983
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24 = -0.0021546
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24 = 0.0099201
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24 = ' -0.031205 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 025, W = 5.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25 = ' -0.025773 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25 = -0.010755
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25 = 0.44696
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25 = 3.0981e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25 = -2.833e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25 = -0.0037504
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25 = -0.0024975
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25 = 0.0057792
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 026, W = 5.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26 = ' -0.037535 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26 = -0.0025585
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26 = 0.26088
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26 = 7.055e-13
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26 = 7.9652e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26 = 0.0034079
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26 = -3120.9
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 027, W = 5.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27 = ' -0.015876 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27 = 0.0028301
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27 = 0.27216
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27 = 2.3477e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27 = 5.7387e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27 = 0.0017998
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27 = -2096.9
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 028, W = 5.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28 = ' -0.03154 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28 = 0.0074722
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28 = 0.29717
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28 = 2.27e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28 = 1.9698e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28 = 0.00015867
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28 = -546.93
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 029, W = 7.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29 = -0.0012422
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29 = 0.0055211
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29 = ' -0.038036 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29 = 0.0051679
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29 = 0.28552
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29 = 1.1207e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29 = -2.2129e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29 = -0.0053554
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 030, W = 7.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30 = -0.0024147
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30 = 0.015899
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30 = ' -0.034674 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30 = -0.0044554
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30 = 0.3274
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30 = 3.371e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30 = -3.0344e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30 = -0.0067289
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 031, W = 7.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31 = -0.0049034
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31 = -0.002325
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31 = 0.005644
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31 = ' -0.03154 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31 = -0.0091003
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31 = 0.37561
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31 = 2.7784e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31 = -3.1676e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 032, W = 7.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32 = -0.0027511
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32 = -0.0028978
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32 = 0.0019878
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32 = ' -0.02821 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32 = -0.010488
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32 = 0.42418
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32 = 3.6729e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32 = -3.6459e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 033, W = 7.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33 = 8.3637e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33 = 0.0040296
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33 = -793.31
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33 = ' -0.035485 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33 = -0.0039041
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33 = 0.22979
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33 = -4.3508e-13
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 034, W = 7.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34 = 0.28064
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34 = 1.5857e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34 = -1.4752e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34 = -0.0011477
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34 = -3415.9
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34 = ' -0.029606 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34 = 0.0072429
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 035, W = 0.42, L = 1.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35 = -0.0044332
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35 = 0.44964
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35 = 1.162e-11
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35 = 1.8897e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35 = -0.003158
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35 = 3.9516e-8
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35 = 5.7202e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35 = ' -0.050123 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 036, W = 0.42, L = 20.0
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36 = ' -0.032204 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36 = -0.0076473
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36 = 0.72918
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36 = 7.145e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36 = -5.0938e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36 = -0.0032011
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36 = -1.4304e-9
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36 = -6.5705e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 037, W = 0.42, L = 2.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37 = ' -0.029618 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37 = -0.0060614
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37 = 0.48503
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37 = 8.8917e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37 = 5.4941e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37 = -0.0029838
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37 = -1.1296e-8
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37 = 2.3412e-9
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 038, W = 0.42, L = 4.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38 = -2.7666e-11
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38 = ' -0.029893 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38 = -0.0052776
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38 = 0.54516
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38 = 8.9623e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38 = 8.5149e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38 = -0.0029895
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38 = -1.6462e-8
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 039, W = 0.42, L = 8.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39 = 1.6548e-9
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39 = 3.4708e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39 = ' -0.03647 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39 = -0.0080677
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39 = 0.61884
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39 = 8.5232e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39 = -3.7718e-20
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39 = -0.0032385
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 040, W = 0.42, L = 0.5
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40 = ' -0.017851 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40 = -0.00065333
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40 = 0.50807
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40 = 2.3883e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40 = 7.4268e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40 = -0.0010841
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40 = -12629.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 041, W = 0.42, L = 0.6
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41 = -0.0027932
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41 = -10499.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41 = ' -0.044571 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41 = -0.0065553
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41 = 0.44784
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41 = 4.3026e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41 = 5.537e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 042, W = 0.42, L = 0.8
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42 = -0.0030568
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42 = -5745.7
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42 = ' -0.072824 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42 = -0.010628
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42 = 0.46794
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42 = 2.7005e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42 = 5.4519e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 043, W = 0.75, L = 1.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43 = -0.0012026
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43 = -3.1092e-8
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43 = 1.5248e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43 = ' -0.023219 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43 = -0.0023873
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43 = 0.46747
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43 = 5.9725e-12
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43 = 2.3384e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 044, W = 0.75, L = 2.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44 = 1.3655e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44 = -0.00095313
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44 = -7.733e-9
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44 = 7.1418e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44 = ' -0.043616 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44 = -0.0091521
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44 = 0.49252
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44 = 4.467e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 045, W = 0.75, L = 4.0
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45 = 0.52792
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45 = 3.7257e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45 = 1.5093e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45 = -0.00093771
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45 = -4.2402e-8
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45 = 3.4216e-10
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45 = ' -0.020684 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45 = -0.013079
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 046, W = 0.75, L = 0.5
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46 = -0.00090328
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46 = 0.5267
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46 = 1.221e-11
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46 = 1.0027e-18
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46 = 0.00020174
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46 = -5377.6
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46 = ' -0.028684 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 047, W = 0.75, L = 0.8
* -------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47 = ' -0.022451 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47 = 0.00054712
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47 = 0.48306
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47 = 6.0929e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47 = 2.6833e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47 = -0.0010186
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47 = -6456.0
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47 = 0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 048, W = 0.7, L = 0.6
* ------------------------------
+ sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48 = ' -0.032032 + sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff'
+ sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48 = 0.0018639
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48 = 0.50359
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48 = 7.1767e-12
+ sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48 = 4.2917e-19
+ sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48 = -0.00059541
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48 = -9162.3
+ sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48 = 0.0
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48 = 0.0
.include "sky130_fd_pr__nfet_g5v0d10v5.pm3.spice"
