# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  22.49000 BY  23.05000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT  0.000000  0.000000 22.490000  0.330000 ;
        RECT  0.000000  0.330000  0.330000 11.360000 ;
        RECT  0.000000 11.360000 22.490000 11.690000 ;
        RECT  0.000000 11.690000  0.330000 22.720000 ;
        RECT  0.000000 22.720000 22.490000 23.050000 ;
        RECT  1.230000  0.330000  1.530000  5.380000 ;
        RECT  1.230000  6.310000  1.530000 11.360000 ;
        RECT  1.230000 11.690000  1.530000 16.740000 ;
        RECT  1.230000 17.670000  1.530000 22.720000 ;
        RECT  2.430000  0.330000  2.730000  5.380000 ;
        RECT  2.430000  6.310000  2.730000 11.360000 ;
        RECT  2.430000 11.690000  2.730000 16.740000 ;
        RECT  2.430000 17.670000  2.730000 22.720000 ;
        RECT  3.630000  0.330000  3.930000  5.380000 ;
        RECT  3.630000  6.310000  3.930000 11.360000 ;
        RECT  3.630000 11.690000  3.930000 16.740000 ;
        RECT  3.630000 17.670000  3.930000 22.720000 ;
        RECT  4.830000  0.330000  5.240000  5.380000 ;
        RECT  4.830000  6.310000  5.240000 11.360000 ;
        RECT  4.830000 11.690000  5.240000 16.740000 ;
        RECT  4.830000 17.670000  5.240000 22.720000 ;
        RECT  6.170000  0.330000  6.580000  5.380000 ;
        RECT  6.170000  6.310000  6.580000 11.360000 ;
        RECT  6.170000 11.690000  6.580000 16.740000 ;
        RECT  6.170000 17.670000  6.580000 22.720000 ;
        RECT  7.480000  0.330000  7.780000  5.380000 ;
        RECT  7.480000  6.310000  7.780000 11.360000 ;
        RECT  7.480000 11.690000  7.780000 16.740000 ;
        RECT  7.480000 17.670000  7.780000 22.720000 ;
        RECT  8.680000  0.330000  8.980000  5.380000 ;
        RECT  8.680000  6.310000  8.980000 11.360000 ;
        RECT  8.680000 11.690000  8.980000 16.740000 ;
        RECT  8.680000 17.670000  8.980000 22.720000 ;
        RECT  9.880000  0.330000 10.180000  5.380000 ;
        RECT  9.880000  6.310000 10.180000 11.360000 ;
        RECT  9.880000 11.690000 10.180000 16.740000 ;
        RECT  9.880000 17.670000 10.180000 22.720000 ;
        RECT 11.080000  0.330000 11.410000 11.360000 ;
        RECT 11.080000 11.690000 11.410000 22.720000 ;
        RECT 12.310000  0.330000 12.610000  5.380000 ;
        RECT 12.310000  6.310000 12.610000 11.360000 ;
        RECT 12.310000 11.690000 12.610000 16.740000 ;
        RECT 12.310000 17.670000 12.610000 22.720000 ;
        RECT 13.510000  0.330000 13.810000  5.380000 ;
        RECT 13.510000  6.310000 13.810000 11.360000 ;
        RECT 13.510000 11.690000 13.810000 16.740000 ;
        RECT 13.510000 17.670000 13.810000 22.720000 ;
        RECT 14.710000  0.330000 15.010000  5.380000 ;
        RECT 14.710000  6.310000 15.010000 11.360000 ;
        RECT 14.710000 11.690000 15.010000 16.740000 ;
        RECT 14.710000 17.670000 15.010000 22.720000 ;
        RECT 15.910000  0.330000 16.320000  5.380000 ;
        RECT 15.910000  6.310000 16.320000 11.360000 ;
        RECT 15.910000 11.690000 16.320000 16.740000 ;
        RECT 15.910000 17.670000 16.320000 22.720000 ;
        RECT 17.250000  0.330000 17.660000  5.380000 ;
        RECT 17.250000  6.310000 17.660000 11.360000 ;
        RECT 17.250000 11.690000 17.660000 16.740000 ;
        RECT 17.250000 17.670000 17.660000 22.720000 ;
        RECT 18.560000  0.330000 18.860000  5.380000 ;
        RECT 18.560000  6.310000 18.860000 11.360000 ;
        RECT 18.560000 11.690000 18.860000 16.740000 ;
        RECT 18.560000 17.670000 18.860000 22.720000 ;
        RECT 19.760000  0.330000 20.060000  5.380000 ;
        RECT 19.760000  6.310000 20.060000 11.360000 ;
        RECT 19.760000 11.690000 20.060000 16.740000 ;
        RECT 19.760000 17.670000 20.060000 22.720000 ;
        RECT 20.960000  0.330000 21.260000  5.380000 ;
        RECT 20.960000  6.310000 21.260000 11.360000 ;
        RECT 20.960000 11.690000 21.260000 16.740000 ;
        RECT 20.960000 17.670000 21.260000 22.720000 ;
        RECT 22.160000  0.330000 22.490000 11.360000 ;
        RECT 22.160000 11.690000 22.490000 22.720000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT  0.630000  0.630000  0.930000  5.680000 ;
        RECT  0.630000  5.680000 10.780000  6.010000 ;
        RECT  0.630000  6.010000  0.930000 11.060000 ;
        RECT  0.630000 11.990000  0.930000 17.040000 ;
        RECT  0.630000 17.040000 10.780000 17.370000 ;
        RECT  0.630000 17.370000  0.930000 22.420000 ;
        RECT  1.830000  0.630000  2.130000  5.680000 ;
        RECT  1.830000  6.010000  2.130000 11.060000 ;
        RECT  1.830000 11.990000  2.130000 17.040000 ;
        RECT  1.830000 17.370000  2.130000 22.420000 ;
        RECT  3.030000  0.630000  3.330000  5.680000 ;
        RECT  3.030000  6.010000  3.330000 11.060000 ;
        RECT  3.030000 11.990000  3.330000 17.040000 ;
        RECT  3.030000 17.370000  3.330000 22.420000 ;
        RECT  4.230000  0.630000  4.530000  5.680000 ;
        RECT  4.230000  6.010000  4.530000 11.060000 ;
        RECT  4.230000 11.990000  4.530000 17.040000 ;
        RECT  4.230000 17.370000  4.530000 22.420000 ;
        RECT  5.540000  0.630000  5.870000  5.680000 ;
        RECT  5.540000  6.010000  5.870000 11.060000 ;
        RECT  5.540000 11.990000  5.870000 17.040000 ;
        RECT  5.540000 17.370000  5.870000 22.420000 ;
        RECT  6.880000  0.630000  7.180000  5.680000 ;
        RECT  6.880000  6.010000  7.180000 11.060000 ;
        RECT  6.880000 11.990000  7.180000 17.040000 ;
        RECT  6.880000 17.370000  7.180000 22.420000 ;
        RECT  8.080000  0.630000  8.380000  5.680000 ;
        RECT  8.080000  6.010000  8.380000 11.060000 ;
        RECT  8.080000 11.990000  8.380000 17.040000 ;
        RECT  8.080000 17.370000  8.380000 22.420000 ;
        RECT  9.280000  0.630000  9.580000  5.680000 ;
        RECT  9.280000  6.010000  9.580000 11.060000 ;
        RECT  9.280000 11.990000  9.580000 17.040000 ;
        RECT  9.280000 17.370000  9.580000 22.420000 ;
        RECT 10.480000  0.630000 10.780000  5.680000 ;
        RECT 10.480000  6.010000 10.780000 11.060000 ;
        RECT 10.480000 11.990000 10.780000 17.040000 ;
        RECT 10.480000 17.370000 10.780000 22.420000 ;
        RECT 11.710000  0.630000 12.010000  5.680000 ;
        RECT 11.710000  5.680000 21.860000  6.010000 ;
        RECT 11.710000  6.010000 12.010000 11.060000 ;
        RECT 11.710000 11.990000 12.010000 17.040000 ;
        RECT 11.710000 17.040000 21.860000 17.370000 ;
        RECT 11.710000 17.370000 12.010000 22.420000 ;
        RECT 12.910000  0.630000 13.210000  5.680000 ;
        RECT 12.910000  6.010000 13.210000 11.060000 ;
        RECT 12.910000 11.990000 13.210000 17.040000 ;
        RECT 12.910000 17.370000 13.210000 22.420000 ;
        RECT 14.110000  0.630000 14.410000  5.680000 ;
        RECT 14.110000  6.010000 14.410000 11.060000 ;
        RECT 14.110000 11.990000 14.410000 17.040000 ;
        RECT 14.110000 17.370000 14.410000 22.420000 ;
        RECT 15.310000  0.630000 15.610000  5.680000 ;
        RECT 15.310000  6.010000 15.610000 11.060000 ;
        RECT 15.310000 11.990000 15.610000 17.040000 ;
        RECT 15.310000 17.370000 15.610000 22.420000 ;
        RECT 16.620000  0.630000 16.950000  5.680000 ;
        RECT 16.620000  6.010000 16.950000 11.060000 ;
        RECT 16.620000 11.990000 16.950000 17.040000 ;
        RECT 16.620000 17.370000 16.950000 22.420000 ;
        RECT 17.960000  0.630000 18.260000  5.680000 ;
        RECT 17.960000  6.010000 18.260000 11.060000 ;
        RECT 17.960000 11.990000 18.260000 17.040000 ;
        RECT 17.960000 17.370000 18.260000 22.420000 ;
        RECT 19.160000  0.630000 19.460000  5.680000 ;
        RECT 19.160000  6.010000 19.460000 11.060000 ;
        RECT 19.160000 11.990000 19.460000 17.040000 ;
        RECT 19.160000 17.370000 19.460000 22.420000 ;
        RECT 20.360000  0.630000 20.660000  5.680000 ;
        RECT 20.360000  6.010000 20.660000 11.060000 ;
        RECT 20.360000 11.990000 20.660000 17.040000 ;
        RECT 20.360000 17.370000 20.660000 22.420000 ;
        RECT 21.560000  0.630000 21.860000  5.680000 ;
        RECT 21.560000  6.010000 21.860000 11.060000 ;
        RECT 21.560000 11.990000 21.860000 17.040000 ;
        RECT 21.560000 17.370000 21.860000 22.420000 ;
    END
  END C1
  PIN M4
    PORT
      LAYER met4 ;
        RECT 0.000000 0.000000 22.490000 23.050000 ;
    END
  END M4
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 5.895000 6.345000 5.945000 6.395000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT  0.000000  0.000000 22.490000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.860000 ;
      RECT  0.000000  0.860000  5.400000  1.030000 ;
      RECT  0.000000  1.030000  0.330000  1.560000 ;
      RECT  0.000000  1.560000  5.400000  1.730000 ;
      RECT  0.000000  1.730000  0.330000  2.260000 ;
      RECT  0.000000  2.260000  5.400000  2.430000 ;
      RECT  0.000000  2.430000  0.330000  2.960000 ;
      RECT  0.000000  2.960000  5.400000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.660000 ;
      RECT  0.000000  3.660000  5.400000  3.830000 ;
      RECT  0.000000  3.830000  0.330000  4.360000 ;
      RECT  0.000000  4.360000  5.400000  4.530000 ;
      RECT  0.000000  4.530000  0.330000  5.060000 ;
      RECT  0.000000  5.060000  5.400000  5.230000 ;
      RECT  0.000000  5.230000  0.330000  5.760000 ;
      RECT  0.000000  5.760000  5.400000  5.930000 ;
      RECT  0.000000  5.930000  0.330000  6.460000 ;
      RECT  0.000000  6.460000  5.400000  6.630000 ;
      RECT  0.000000  6.630000  0.330000  7.150000 ;
      RECT  0.000000  7.150000  5.400000  7.330000 ;
      RECT  0.000000  7.330000  0.330000  7.860000 ;
      RECT  0.000000  7.860000  5.400000  8.030000 ;
      RECT  0.000000  8.030000  0.330000  8.560000 ;
      RECT  0.000000  8.560000  5.400000  8.730000 ;
      RECT  0.000000  8.730000  0.330000  9.260000 ;
      RECT  0.000000  9.260000  5.400000  9.430000 ;
      RECT  0.000000  9.430000  0.330000  9.960000 ;
      RECT  0.000000  9.960000  5.400000 10.130000 ;
      RECT  0.000000 10.130000  0.330000 10.660000 ;
      RECT  0.000000 10.660000  5.400000 10.830000 ;
      RECT  0.000000 10.830000  0.330000 11.360000 ;
      RECT  0.000000 11.360000 22.490000 11.690000 ;
      RECT  0.000000 11.690000  0.330000 12.220000 ;
      RECT  0.000000 12.220000  5.400000 12.390000 ;
      RECT  0.000000 12.390000  0.330000 12.920000 ;
      RECT  0.000000 12.920000  5.400000 13.090000 ;
      RECT  0.000000 13.090000  0.330000 13.620000 ;
      RECT  0.000000 13.620000  5.400000 13.790000 ;
      RECT  0.000000 13.790000  0.330000 14.320000 ;
      RECT  0.000000 14.320000  5.400000 14.490000 ;
      RECT  0.000000 14.490000  0.330000 15.020000 ;
      RECT  0.000000 15.020000  5.400000 15.190000 ;
      RECT  0.000000 15.190000  0.330000 15.720000 ;
      RECT  0.000000 15.720000  5.400000 15.890000 ;
      RECT  0.000000 15.890000  0.330000 16.420000 ;
      RECT  0.000000 16.420000  5.400000 16.590000 ;
      RECT  0.000000 16.590000  0.330000 17.120000 ;
      RECT  0.000000 17.120000  5.400000 17.290000 ;
      RECT  0.000000 17.290000  0.330000 17.820000 ;
      RECT  0.000000 17.820000  5.400000 17.990000 ;
      RECT  0.000000 17.990000  0.330000 18.510000 ;
      RECT  0.000000 18.510000  5.400000 18.690000 ;
      RECT  0.000000 18.690000  0.330000 19.220000 ;
      RECT  0.000000 19.220000  5.400000 19.390000 ;
      RECT  0.000000 19.390000  0.330000 19.920000 ;
      RECT  0.000000 19.920000  5.400000 20.090000 ;
      RECT  0.000000 20.090000  0.330000 20.620000 ;
      RECT  0.000000 20.620000  5.400000 20.790000 ;
      RECT  0.000000 20.790000  0.330000 21.320000 ;
      RECT  0.000000 21.320000  5.400000 21.490000 ;
      RECT  0.000000 21.490000  0.330000 22.020000 ;
      RECT  0.000000 22.020000  5.400000 22.190000 ;
      RECT  0.000000 22.190000  0.330000 22.720000 ;
      RECT  0.000000 22.720000 22.490000 23.050000 ;
      RECT  0.500000  0.500000 10.905000  0.690000 ;
      RECT  0.500000  1.200000 10.905000  1.390000 ;
      RECT  0.500000  1.900000 10.905000  2.090000 ;
      RECT  0.500000  2.600000 10.905000  2.790000 ;
      RECT  0.500000  3.300000 10.905000  3.490000 ;
      RECT  0.500000  4.000000 10.905000  4.190000 ;
      RECT  0.500000  4.700000 10.905000  4.890000 ;
      RECT  0.500000  5.400000 10.905000  5.590000 ;
      RECT  0.500000  6.100000 10.905000  6.290000 ;
      RECT  0.500000  6.800000 10.905000  6.980000 ;
      RECT  0.500000  7.500000 10.905000  7.690000 ;
      RECT  0.500000  8.200000 10.905000  8.390000 ;
      RECT  0.500000  8.900000 10.905000  9.090000 ;
      RECT  0.500000  9.600000 10.905000  9.790000 ;
      RECT  0.500000 10.300000 10.905000 10.490000 ;
      RECT  0.500000 11.000000 10.905000 11.190000 ;
      RECT  0.500000 11.860000 10.905000 12.050000 ;
      RECT  0.500000 12.560000 10.905000 12.750000 ;
      RECT  0.500000 13.260000 10.905000 13.450000 ;
      RECT  0.500000 13.960000 10.905000 14.150000 ;
      RECT  0.500000 14.660000 10.905000 14.850000 ;
      RECT  0.500000 15.360000 10.905000 15.550000 ;
      RECT  0.500000 16.060000 10.905000 16.250000 ;
      RECT  0.500000 16.760000 10.905000 16.950000 ;
      RECT  0.500000 17.460000 10.905000 17.650000 ;
      RECT  0.500000 18.160000 10.905000 18.340000 ;
      RECT  0.500000 18.860000 10.905000 19.050000 ;
      RECT  0.500000 19.560000 10.905000 19.750000 ;
      RECT  0.500000 20.260000 10.905000 20.450000 ;
      RECT  0.500000 20.960000 10.905000 21.150000 ;
      RECT  0.500000 21.660000 10.905000 21.850000 ;
      RECT  0.500000 22.360000 10.905000 22.550000 ;
      RECT  5.570000  0.690000  5.840000  1.200000 ;
      RECT  5.570000  1.390000  5.840000  1.900000 ;
      RECT  5.570000  2.090000  5.840000  2.600000 ;
      RECT  5.570000  2.790000  5.840000  3.300000 ;
      RECT  5.570000  3.490000  5.840000  4.000000 ;
      RECT  5.570000  4.190000  5.840000  4.700000 ;
      RECT  5.570000  4.890000  5.840000  5.400000 ;
      RECT  5.570000  5.590000  5.840000  6.100000 ;
      RECT  5.570000  6.290000  5.840000  6.800000 ;
      RECT  5.570000  6.980000 10.905000  6.990000 ;
      RECT  5.570000  6.990000  5.840000  7.500000 ;
      RECT  5.570000  7.690000  5.840000  8.200000 ;
      RECT  5.570000  8.390000  5.840000  8.900000 ;
      RECT  5.570000  9.090000  5.840000  9.600000 ;
      RECT  5.570000  9.790000  5.840000 10.300000 ;
      RECT  5.570000 10.490000  5.840000 11.000000 ;
      RECT  5.570000 12.050000  5.840000 12.560000 ;
      RECT  5.570000 12.750000  5.840000 13.260000 ;
      RECT  5.570000 13.450000  5.840000 13.960000 ;
      RECT  5.570000 14.150000  5.840000 14.660000 ;
      RECT  5.570000 14.850000  5.840000 15.360000 ;
      RECT  5.570000 15.550000  5.840000 16.060000 ;
      RECT  5.570000 16.250000  5.840000 16.760000 ;
      RECT  5.570000 16.950000  5.840000 17.460000 ;
      RECT  5.570000 17.650000  5.840000 18.160000 ;
      RECT  5.570000 18.340000 10.905000 18.350000 ;
      RECT  5.570000 18.350000  5.840000 18.860000 ;
      RECT  5.570000 19.050000  5.840000 19.560000 ;
      RECT  5.570000 19.750000  5.840000 20.260000 ;
      RECT  5.570000 20.450000  5.840000 20.960000 ;
      RECT  5.570000 21.150000  5.840000 21.660000 ;
      RECT  5.570000 21.850000  5.840000 22.360000 ;
      RECT  6.010000  0.860000 16.480000  1.030000 ;
      RECT  6.010000  1.560000 16.480000  1.730000 ;
      RECT  6.010000  2.260000 16.480000  2.430000 ;
      RECT  6.010000  2.960000 16.480000  3.130000 ;
      RECT  6.010000  3.660000 16.480000  3.830000 ;
      RECT  6.010000  4.360000 16.480000  4.530000 ;
      RECT  6.010000  5.060000 16.480000  5.230000 ;
      RECT  6.010000  5.760000 16.480000  5.930000 ;
      RECT  6.010000  6.460000 16.480000  6.630000 ;
      RECT  6.010000  7.160000 16.480000  7.330000 ;
      RECT  6.010000  7.860000 16.480000  8.030000 ;
      RECT  6.010000  8.560000 16.480000  8.730000 ;
      RECT  6.010000  9.260000 16.480000  9.430000 ;
      RECT  6.010000  9.960000 16.480000 10.130000 ;
      RECT  6.010000 10.660000 16.480000 10.830000 ;
      RECT  6.010000 12.220000 16.480000 12.390000 ;
      RECT  6.010000 12.920000 16.480000 13.090000 ;
      RECT  6.010000 13.620000 16.480000 13.790000 ;
      RECT  6.010000 14.320000 16.480000 14.490000 ;
      RECT  6.010000 15.020000 16.480000 15.190000 ;
      RECT  6.010000 15.720000 16.480000 15.890000 ;
      RECT  6.010000 16.420000 16.480000 16.590000 ;
      RECT  6.010000 17.120000 16.480000 17.290000 ;
      RECT  6.010000 17.820000 16.480000 17.990000 ;
      RECT  6.010000 18.520000 16.480000 18.690000 ;
      RECT  6.010000 19.220000 16.480000 19.390000 ;
      RECT  6.010000 19.920000 16.480000 20.090000 ;
      RECT  6.010000 20.620000 16.480000 20.790000 ;
      RECT  6.010000 21.320000 16.480000 21.490000 ;
      RECT  6.010000 22.020000 16.480000 22.190000 ;
      RECT 11.080000  0.330000 11.410000  0.860000 ;
      RECT 11.080000  1.030000 11.410000  1.560000 ;
      RECT 11.080000  1.730000 11.410000  2.260000 ;
      RECT 11.080000  2.430000 11.410000  2.960000 ;
      RECT 11.080000  3.130000 11.410000  3.660000 ;
      RECT 11.080000  3.830000 11.410000  4.360000 ;
      RECT 11.080000  4.530000 11.410000  5.060000 ;
      RECT 11.080000  5.230000 11.410000  5.760000 ;
      RECT 11.080000  5.930000 11.410000  6.460000 ;
      RECT 11.080000  6.630000 11.410000  7.150000 ;
      RECT 11.080000  7.150000 16.480000  7.160000 ;
      RECT 11.080000  7.330000 11.410000  7.860000 ;
      RECT 11.080000  8.030000 11.410000  8.560000 ;
      RECT 11.080000  8.730000 11.410000  9.260000 ;
      RECT 11.080000  9.430000 11.410000  9.960000 ;
      RECT 11.080000 10.130000 11.410000 10.660000 ;
      RECT 11.080000 10.830000 11.410000 11.360000 ;
      RECT 11.080000 11.690000 11.410000 12.220000 ;
      RECT 11.080000 12.390000 11.410000 12.920000 ;
      RECT 11.080000 13.090000 11.410000 13.620000 ;
      RECT 11.080000 13.790000 11.410000 14.320000 ;
      RECT 11.080000 14.490000 11.410000 15.020000 ;
      RECT 11.080000 15.190000 11.410000 15.720000 ;
      RECT 11.080000 15.890000 11.410000 16.420000 ;
      RECT 11.080000 16.590000 11.410000 17.120000 ;
      RECT 11.080000 17.290000 11.410000 17.820000 ;
      RECT 11.080000 17.990000 11.410000 18.510000 ;
      RECT 11.080000 18.510000 16.480000 18.520000 ;
      RECT 11.080000 18.690000 11.410000 19.220000 ;
      RECT 11.080000 19.390000 11.410000 19.920000 ;
      RECT 11.080000 20.090000 11.410000 20.620000 ;
      RECT 11.080000 20.790000 11.410000 21.320000 ;
      RECT 11.080000 21.490000 11.410000 22.020000 ;
      RECT 11.080000 22.190000 11.410000 22.720000 ;
      RECT 11.580000  0.500000 21.985000  0.690000 ;
      RECT 11.580000  1.200000 21.985000  1.390000 ;
      RECT 11.580000  1.900000 21.985000  2.090000 ;
      RECT 11.580000  2.600000 21.985000  2.790000 ;
      RECT 11.580000  3.300000 21.985000  3.490000 ;
      RECT 11.580000  4.000000 21.985000  4.190000 ;
      RECT 11.580000  4.700000 21.985000  4.890000 ;
      RECT 11.580000  5.400000 21.985000  5.590000 ;
      RECT 11.580000  6.100000 21.985000  6.290000 ;
      RECT 11.580000  6.800000 21.985000  6.980000 ;
      RECT 11.580000  7.500000 21.985000  7.690000 ;
      RECT 11.580000  8.200000 21.985000  8.390000 ;
      RECT 11.580000  8.900000 21.985000  9.090000 ;
      RECT 11.580000  9.600000 21.985000  9.790000 ;
      RECT 11.580000 10.300000 21.985000 10.490000 ;
      RECT 11.580000 11.000000 21.985000 11.190000 ;
      RECT 11.580000 11.860000 21.985000 12.050000 ;
      RECT 11.580000 12.560000 21.985000 12.750000 ;
      RECT 11.580000 13.260000 21.985000 13.450000 ;
      RECT 11.580000 13.960000 21.985000 14.150000 ;
      RECT 11.580000 14.660000 21.985000 14.850000 ;
      RECT 11.580000 15.360000 21.985000 15.550000 ;
      RECT 11.580000 16.060000 21.985000 16.250000 ;
      RECT 11.580000 16.760000 21.985000 16.950000 ;
      RECT 11.580000 17.460000 21.985000 17.650000 ;
      RECT 11.580000 18.160000 21.985000 18.340000 ;
      RECT 11.580000 18.860000 21.985000 19.050000 ;
      RECT 11.580000 19.560000 21.985000 19.750000 ;
      RECT 11.580000 20.260000 21.985000 20.450000 ;
      RECT 11.580000 20.960000 21.985000 21.150000 ;
      RECT 11.580000 21.660000 21.985000 21.850000 ;
      RECT 11.580000 22.360000 21.985000 22.550000 ;
      RECT 16.650000  0.690000 16.920000  1.200000 ;
      RECT 16.650000  1.390000 16.920000  1.900000 ;
      RECT 16.650000  2.090000 16.920000  2.600000 ;
      RECT 16.650000  2.790000 16.920000  3.300000 ;
      RECT 16.650000  3.490000 16.920000  4.000000 ;
      RECT 16.650000  4.190000 16.920000  4.700000 ;
      RECT 16.650000  4.890000 16.920000  5.400000 ;
      RECT 16.650000  5.590000 16.920000  6.100000 ;
      RECT 16.650000  6.290000 16.920000  6.800000 ;
      RECT 16.650000  6.980000 21.985000  6.990000 ;
      RECT 16.650000  6.990000 16.920000  7.500000 ;
      RECT 16.650000  7.690000 16.920000  8.200000 ;
      RECT 16.650000  8.390000 16.920000  8.900000 ;
      RECT 16.650000  9.090000 16.920000  9.600000 ;
      RECT 16.650000  9.790000 16.920000 10.300000 ;
      RECT 16.650000 10.490000 16.920000 11.000000 ;
      RECT 16.650000 12.050000 16.920000 12.560000 ;
      RECT 16.650000 12.750000 16.920000 13.260000 ;
      RECT 16.650000 13.450000 16.920000 13.960000 ;
      RECT 16.650000 14.150000 16.920000 14.660000 ;
      RECT 16.650000 14.850000 16.920000 15.360000 ;
      RECT 16.650000 15.550000 16.920000 16.060000 ;
      RECT 16.650000 16.250000 16.920000 16.760000 ;
      RECT 16.650000 16.950000 16.920000 17.460000 ;
      RECT 16.650000 17.650000 16.920000 18.160000 ;
      RECT 16.650000 18.340000 21.985000 18.350000 ;
      RECT 16.650000 18.350000 16.920000 18.860000 ;
      RECT 16.650000 19.050000 16.920000 19.560000 ;
      RECT 16.650000 19.750000 16.920000 20.260000 ;
      RECT 16.650000 20.450000 16.920000 20.960000 ;
      RECT 16.650000 21.150000 16.920000 21.660000 ;
      RECT 16.650000 21.850000 16.920000 22.360000 ;
      RECT 17.090000  0.860000 22.490000  1.030000 ;
      RECT 17.090000  1.560000 22.490000  1.730000 ;
      RECT 17.090000  2.260000 22.490000  2.430000 ;
      RECT 17.090000  2.960000 22.490000  3.130000 ;
      RECT 17.090000  3.660000 22.490000  3.830000 ;
      RECT 17.090000  4.360000 22.490000  4.530000 ;
      RECT 17.090000  5.060000 22.490000  5.230000 ;
      RECT 17.090000  5.760000 22.490000  5.930000 ;
      RECT 17.090000  6.460000 22.490000  6.630000 ;
      RECT 17.090000  7.160000 22.490000  7.330000 ;
      RECT 17.090000  7.860000 22.490000  8.030000 ;
      RECT 17.090000  8.560000 22.490000  8.730000 ;
      RECT 17.090000  9.260000 22.490000  9.430000 ;
      RECT 17.090000  9.960000 22.490000 10.130000 ;
      RECT 17.090000 10.660000 22.490000 10.830000 ;
      RECT 17.090000 12.220000 22.490000 12.390000 ;
      RECT 17.090000 12.920000 22.490000 13.090000 ;
      RECT 17.090000 13.620000 22.490000 13.790000 ;
      RECT 17.090000 14.320000 22.490000 14.490000 ;
      RECT 17.090000 15.020000 22.490000 15.190000 ;
      RECT 17.090000 15.720000 22.490000 15.890000 ;
      RECT 17.090000 16.420000 22.490000 16.590000 ;
      RECT 17.090000 17.120000 22.490000 17.290000 ;
      RECT 17.090000 17.820000 22.490000 17.990000 ;
      RECT 17.090000 18.520000 22.490000 18.690000 ;
      RECT 17.090000 19.220000 22.490000 19.390000 ;
      RECT 17.090000 19.920000 22.490000 20.090000 ;
      RECT 17.090000 20.620000 22.490000 20.790000 ;
      RECT 17.090000 21.320000 22.490000 21.490000 ;
      RECT 17.090000 22.020000 22.490000 22.190000 ;
      RECT 22.160000  0.330000 22.490000  0.860000 ;
      RECT 22.160000  1.030000 22.490000  1.560000 ;
      RECT 22.160000  1.730000 22.490000  2.260000 ;
      RECT 22.160000  2.430000 22.490000  2.960000 ;
      RECT 22.160000  3.130000 22.490000  3.660000 ;
      RECT 22.160000  3.830000 22.490000  4.360000 ;
      RECT 22.160000  4.530000 22.490000  5.060000 ;
      RECT 22.160000  5.230000 22.490000  5.760000 ;
      RECT 22.160000  5.930000 22.490000  6.460000 ;
      RECT 22.160000  6.630000 22.490000  7.160000 ;
      RECT 22.160000  7.330000 22.490000  7.860000 ;
      RECT 22.160000  8.030000 22.490000  8.560000 ;
      RECT 22.160000  8.730000 22.490000  9.260000 ;
      RECT 22.160000  9.430000 22.490000  9.960000 ;
      RECT 22.160000 10.130000 22.490000 10.660000 ;
      RECT 22.160000 10.830000 22.490000 11.360000 ;
      RECT 22.160000 11.690000 22.490000 12.220000 ;
      RECT 22.160000 12.390000 22.490000 12.920000 ;
      RECT 22.160000 13.090000 22.490000 13.620000 ;
      RECT 22.160000 13.790000 22.490000 14.320000 ;
      RECT 22.160000 14.490000 22.490000 15.020000 ;
      RECT 22.160000 15.190000 22.490000 15.720000 ;
      RECT 22.160000 15.890000 22.490000 16.420000 ;
      RECT 22.160000 16.590000 22.490000 17.120000 ;
      RECT 22.160000 17.290000 22.490000 17.820000 ;
      RECT 22.160000 17.990000 22.490000 18.520000 ;
      RECT 22.160000 18.690000 22.490000 19.220000 ;
      RECT 22.160000 19.390000 22.490000 19.920000 ;
      RECT 22.160000 20.090000 22.490000 20.620000 ;
      RECT 22.160000 20.790000 22.490000 21.320000 ;
      RECT 22.160000 21.490000 22.490000 22.020000 ;
      RECT 22.160000 22.190000 22.490000 22.720000 ;
    LAYER mcon ;
      RECT  0.080000  0.580000  0.250000  0.750000 ;
      RECT  0.080000  0.940000  0.250000  1.110000 ;
      RECT  0.080000  1.300000  0.250000  1.470000 ;
      RECT  0.080000  1.660000  0.250000  1.830000 ;
      RECT  0.080000  2.020000  0.250000  2.190000 ;
      RECT  0.080000  2.380000  0.250000  2.550000 ;
      RECT  0.080000  2.740000  0.250000  2.910000 ;
      RECT  0.080000  3.100000  0.250000  3.270000 ;
      RECT  0.080000  3.460000  0.250000  3.630000 ;
      RECT  0.080000  3.820000  0.250000  3.990000 ;
      RECT  0.080000  4.180000  0.250000  4.350000 ;
      RECT  0.080000  4.540000  0.250000  4.710000 ;
      RECT  0.080000  4.900000  0.250000  5.070000 ;
      RECT  0.080000  5.260000  0.250000  5.430000 ;
      RECT  0.080000  6.260000  0.250000  6.430000 ;
      RECT  0.080000  6.620000  0.250000  6.790000 ;
      RECT  0.080000  6.980000  0.250000  7.150000 ;
      RECT  0.080000  7.340000  0.250000  7.510000 ;
      RECT  0.080000  7.700000  0.250000  7.870000 ;
      RECT  0.080000  8.060000  0.250000  8.230000 ;
      RECT  0.080000  8.420000  0.250000  8.590000 ;
      RECT  0.080000  8.780000  0.250000  8.950000 ;
      RECT  0.080000  9.140000  0.250000  9.310000 ;
      RECT  0.080000  9.500000  0.250000  9.670000 ;
      RECT  0.080000  9.860000  0.250000 10.030000 ;
      RECT  0.080000 10.220000  0.250000 10.390000 ;
      RECT  0.080000 10.580000  0.250000 10.750000 ;
      RECT  0.080000 10.940000  0.250000 11.110000 ;
      RECT  0.080000 11.940000  0.250000 12.110000 ;
      RECT  0.080000 12.300000  0.250000 12.470000 ;
      RECT  0.080000 12.660000  0.250000 12.830000 ;
      RECT  0.080000 13.020000  0.250000 13.190000 ;
      RECT  0.080000 13.380000  0.250000 13.550000 ;
      RECT  0.080000 13.740000  0.250000 13.910000 ;
      RECT  0.080000 14.100000  0.250000 14.270000 ;
      RECT  0.080000 14.460000  0.250000 14.630000 ;
      RECT  0.080000 14.820000  0.250000 14.990000 ;
      RECT  0.080000 15.180000  0.250000 15.350000 ;
      RECT  0.080000 15.540000  0.250000 15.710000 ;
      RECT  0.080000 15.900000  0.250000 16.070000 ;
      RECT  0.080000 16.260000  0.250000 16.430000 ;
      RECT  0.080000 16.620000  0.250000 16.790000 ;
      RECT  0.080000 17.620000  0.250000 17.790000 ;
      RECT  0.080000 17.980000  0.250000 18.150000 ;
      RECT  0.080000 18.340000  0.250000 18.510000 ;
      RECT  0.080000 18.700000  0.250000 18.870000 ;
      RECT  0.080000 19.060000  0.250000 19.230000 ;
      RECT  0.080000 19.420000  0.250000 19.590000 ;
      RECT  0.080000 19.780000  0.250000 19.950000 ;
      RECT  0.080000 20.140000  0.250000 20.310000 ;
      RECT  0.080000 20.500000  0.250000 20.670000 ;
      RECT  0.080000 20.860000  0.250000 21.030000 ;
      RECT  0.080000 21.220000  0.250000 21.390000 ;
      RECT  0.080000 21.580000  0.250000 21.750000 ;
      RECT  0.080000 21.940000  0.250000 22.110000 ;
      RECT  0.080000 22.300000  0.250000 22.470000 ;
      RECT  0.400000  0.080000  0.570000  0.250000 ;
      RECT  0.400000 11.440000  0.570000 11.610000 ;
      RECT  0.400000 22.800000  0.570000 22.970000 ;
      RECT  0.760000  0.080000  0.930000  0.250000 ;
      RECT  0.760000 11.440000  0.930000 11.610000 ;
      RECT  0.760000 22.800000  0.930000 22.970000 ;
      RECT  1.120000  0.080000  1.290000  0.250000 ;
      RECT  1.120000 11.440000  1.290000 11.610000 ;
      RECT  1.120000 22.800000  1.290000 22.970000 ;
      RECT  1.480000  0.080000  1.650000  0.250000 ;
      RECT  1.480000 11.440000  1.650000 11.610000 ;
      RECT  1.480000 22.800000  1.650000 22.970000 ;
      RECT  1.840000  0.080000  2.010000  0.250000 ;
      RECT  1.840000 11.440000  2.010000 11.610000 ;
      RECT  1.840000 22.800000  2.010000 22.970000 ;
      RECT  2.200000  0.080000  2.370000  0.250000 ;
      RECT  2.200000 11.440000  2.370000 11.610000 ;
      RECT  2.200000 22.800000  2.370000 22.970000 ;
      RECT  2.560000  0.080000  2.730000  0.250000 ;
      RECT  2.560000 11.440000  2.730000 11.610000 ;
      RECT  2.560000 22.800000  2.730000 22.970000 ;
      RECT  2.920000  0.080000  3.090000  0.250000 ;
      RECT  2.920000 11.440000  3.090000 11.610000 ;
      RECT  2.920000 22.800000  3.090000 22.970000 ;
      RECT  3.280000  0.080000  3.450000  0.250000 ;
      RECT  3.280000 11.440000  3.450000 11.610000 ;
      RECT  3.280000 22.800000  3.450000 22.970000 ;
      RECT  3.640000  0.080000  3.810000  0.250000 ;
      RECT  3.640000 11.440000  3.810000 11.610000 ;
      RECT  3.640000 22.800000  3.810000 22.970000 ;
      RECT  4.000000  0.080000  4.170000  0.250000 ;
      RECT  4.000000 11.440000  4.170000 11.610000 ;
      RECT  4.000000 22.800000  4.170000 22.970000 ;
      RECT  4.360000  0.080000  4.530000  0.250000 ;
      RECT  4.360000 11.440000  4.530000 11.610000 ;
      RECT  4.360000 22.800000  4.530000 22.970000 ;
      RECT  4.720000  0.080000  4.890000  0.250000 ;
      RECT  4.720000 11.440000  4.890000 11.610000 ;
      RECT  4.720000 22.800000  4.890000 22.970000 ;
      RECT  5.080000  0.080000  5.250000  0.250000 ;
      RECT  5.080000 11.440000  5.250000 11.610000 ;
      RECT  5.080000 22.800000  5.250000 22.970000 ;
      RECT  5.440000  0.080000  5.610000  0.250000 ;
      RECT  5.440000 11.440000  5.610000 11.610000 ;
      RECT  5.440000 22.800000  5.610000 22.970000 ;
      RECT  5.620000  0.590000  5.790000  0.760000 ;
      RECT  5.620000  0.950000  5.790000  1.120000 ;
      RECT  5.620000  1.310000  5.790000  1.480000 ;
      RECT  5.620000  1.670000  5.790000  1.840000 ;
      RECT  5.620000  2.030000  5.790000  2.200000 ;
      RECT  5.620000  2.390000  5.790000  2.560000 ;
      RECT  5.620000  2.750000  5.790000  2.920000 ;
      RECT  5.620000  3.110000  5.790000  3.280000 ;
      RECT  5.620000  3.470000  5.790000  3.640000 ;
      RECT  5.620000  3.830000  5.790000  4.000000 ;
      RECT  5.620000  4.190000  5.790000  4.360000 ;
      RECT  5.620000  4.550000  5.790000  4.720000 ;
      RECT  5.620000  4.910000  5.790000  5.080000 ;
      RECT  5.620000  5.270000  5.790000  5.440000 ;
      RECT  5.620000  6.250000  5.790000  6.420000 ;
      RECT  5.620000  6.610000  5.790000  6.780000 ;
      RECT  5.620000  6.970000  5.790000  7.140000 ;
      RECT  5.620000  7.330000  5.790000  7.500000 ;
      RECT  5.620000  7.690000  5.790000  7.860000 ;
      RECT  5.620000  8.050000  5.790000  8.220000 ;
      RECT  5.620000  8.410000  5.790000  8.580000 ;
      RECT  5.620000  8.770000  5.790000  8.940000 ;
      RECT  5.620000  9.130000  5.790000  9.300000 ;
      RECT  5.620000  9.490000  5.790000  9.660000 ;
      RECT  5.620000  9.850000  5.790000 10.020000 ;
      RECT  5.620000 10.210000  5.790000 10.380000 ;
      RECT  5.620000 10.570000  5.790000 10.740000 ;
      RECT  5.620000 10.930000  5.790000 11.100000 ;
      RECT  5.620000 11.950000  5.790000 12.120000 ;
      RECT  5.620000 12.310000  5.790000 12.480000 ;
      RECT  5.620000 12.670000  5.790000 12.840000 ;
      RECT  5.620000 13.030000  5.790000 13.200000 ;
      RECT  5.620000 13.390000  5.790000 13.560000 ;
      RECT  5.620000 13.750000  5.790000 13.920000 ;
      RECT  5.620000 14.110000  5.790000 14.280000 ;
      RECT  5.620000 14.470000  5.790000 14.640000 ;
      RECT  5.620000 14.830000  5.790000 15.000000 ;
      RECT  5.620000 15.190000  5.790000 15.360000 ;
      RECT  5.620000 15.550000  5.790000 15.720000 ;
      RECT  5.620000 15.910000  5.790000 16.080000 ;
      RECT  5.620000 16.270000  5.790000 16.440000 ;
      RECT  5.620000 16.630000  5.790000 16.800000 ;
      RECT  5.620000 17.610000  5.790000 17.780000 ;
      RECT  5.620000 17.970000  5.790000 18.140000 ;
      RECT  5.620000 18.330000  5.790000 18.500000 ;
      RECT  5.620000 18.690000  5.790000 18.860000 ;
      RECT  5.620000 19.050000  5.790000 19.220000 ;
      RECT  5.620000 19.410000  5.790000 19.580000 ;
      RECT  5.620000 19.770000  5.790000 19.940000 ;
      RECT  5.620000 20.130000  5.790000 20.300000 ;
      RECT  5.620000 20.490000  5.790000 20.660000 ;
      RECT  5.620000 20.850000  5.790000 21.020000 ;
      RECT  5.620000 21.210000  5.790000 21.380000 ;
      RECT  5.620000 21.570000  5.790000 21.740000 ;
      RECT  5.620000 21.930000  5.790000 22.100000 ;
      RECT  5.620000 22.290000  5.790000 22.460000 ;
      RECT  5.800000  0.080000  5.970000  0.250000 ;
      RECT  5.800000 11.440000  5.970000 11.610000 ;
      RECT  5.800000 22.800000  5.970000 22.970000 ;
      RECT  6.160000  0.080000  6.330000  0.250000 ;
      RECT  6.160000 11.440000  6.330000 11.610000 ;
      RECT  6.160000 22.800000  6.330000 22.970000 ;
      RECT  6.520000  0.080000  6.690000  0.250000 ;
      RECT  6.520000 11.440000  6.690000 11.610000 ;
      RECT  6.520000 22.800000  6.690000 22.970000 ;
      RECT  6.880000  0.080000  7.050000  0.250000 ;
      RECT  6.880000 11.440000  7.050000 11.610000 ;
      RECT  6.880000 22.800000  7.050000 22.970000 ;
      RECT  7.240000  0.080000  7.410000  0.250000 ;
      RECT  7.240000 11.440000  7.410000 11.610000 ;
      RECT  7.240000 22.800000  7.410000 22.970000 ;
      RECT  7.600000  0.080000  7.770000  0.250000 ;
      RECT  7.600000 11.440000  7.770000 11.610000 ;
      RECT  7.600000 22.800000  7.770000 22.970000 ;
      RECT  7.960000  0.080000  8.130000  0.250000 ;
      RECT  7.960000 11.440000  8.130000 11.610000 ;
      RECT  7.960000 22.800000  8.130000 22.970000 ;
      RECT  8.320000  0.080000  8.490000  0.250000 ;
      RECT  8.320000 11.440000  8.490000 11.610000 ;
      RECT  8.320000 22.800000  8.490000 22.970000 ;
      RECT  8.680000  0.080000  8.850000  0.250000 ;
      RECT  8.680000 11.440000  8.850000 11.610000 ;
      RECT  8.680000 22.800000  8.850000 22.970000 ;
      RECT  9.040000  0.080000  9.210000  0.250000 ;
      RECT  9.040000 11.440000  9.210000 11.610000 ;
      RECT  9.040000 22.800000  9.210000 22.970000 ;
      RECT  9.400000  0.080000  9.570000  0.250000 ;
      RECT  9.400000 11.440000  9.570000 11.610000 ;
      RECT  9.400000 22.800000  9.570000 22.970000 ;
      RECT  9.760000  0.080000  9.930000  0.250000 ;
      RECT  9.760000 11.440000  9.930000 11.610000 ;
      RECT  9.760000 22.800000  9.930000 22.970000 ;
      RECT 10.120000  0.080000 10.290000  0.250000 ;
      RECT 10.120000 11.440000 10.290000 11.610000 ;
      RECT 10.120000 22.800000 10.290000 22.970000 ;
      RECT 10.480000  0.080000 10.650000  0.250000 ;
      RECT 10.480000 11.440000 10.650000 11.610000 ;
      RECT 10.480000 22.800000 10.650000 22.970000 ;
      RECT 10.840000  0.080000 11.010000  0.250000 ;
      RECT 10.840000 11.440000 11.010000 11.610000 ;
      RECT 10.840000 22.800000 11.010000 22.970000 ;
      RECT 11.160000  0.580000 11.330000  0.750000 ;
      RECT 11.160000  0.940000 11.330000  1.110000 ;
      RECT 11.160000  1.300000 11.330000  1.470000 ;
      RECT 11.160000  1.660000 11.330000  1.830000 ;
      RECT 11.160000  2.020000 11.330000  2.190000 ;
      RECT 11.160000  2.380000 11.330000  2.550000 ;
      RECT 11.160000  2.740000 11.330000  2.910000 ;
      RECT 11.160000  3.100000 11.330000  3.270000 ;
      RECT 11.160000  3.460000 11.330000  3.630000 ;
      RECT 11.160000  3.820000 11.330000  3.990000 ;
      RECT 11.160000  4.180000 11.330000  4.350000 ;
      RECT 11.160000  4.540000 11.330000  4.710000 ;
      RECT 11.160000  4.900000 11.330000  5.070000 ;
      RECT 11.160000  5.260000 11.330000  5.430000 ;
      RECT 11.160000  6.260000 11.330000  6.430000 ;
      RECT 11.160000  6.620000 11.330000  6.790000 ;
      RECT 11.160000  6.980000 11.330000  7.150000 ;
      RECT 11.160000  7.340000 11.330000  7.510000 ;
      RECT 11.160000  7.700000 11.330000  7.870000 ;
      RECT 11.160000  8.060000 11.330000  8.230000 ;
      RECT 11.160000  8.420000 11.330000  8.590000 ;
      RECT 11.160000  8.780000 11.330000  8.950000 ;
      RECT 11.160000  9.140000 11.330000  9.310000 ;
      RECT 11.160000  9.500000 11.330000  9.670000 ;
      RECT 11.160000  9.860000 11.330000 10.030000 ;
      RECT 11.160000 10.220000 11.330000 10.390000 ;
      RECT 11.160000 10.580000 11.330000 10.750000 ;
      RECT 11.160000 10.940000 11.330000 11.110000 ;
      RECT 11.160000 11.940000 11.330000 12.110000 ;
      RECT 11.160000 12.300000 11.330000 12.470000 ;
      RECT 11.160000 12.660000 11.330000 12.830000 ;
      RECT 11.160000 13.020000 11.330000 13.190000 ;
      RECT 11.160000 13.380000 11.330000 13.550000 ;
      RECT 11.160000 13.740000 11.330000 13.910000 ;
      RECT 11.160000 14.100000 11.330000 14.270000 ;
      RECT 11.160000 14.460000 11.330000 14.630000 ;
      RECT 11.160000 14.820000 11.330000 14.990000 ;
      RECT 11.160000 15.180000 11.330000 15.350000 ;
      RECT 11.160000 15.540000 11.330000 15.710000 ;
      RECT 11.160000 15.900000 11.330000 16.070000 ;
      RECT 11.160000 16.260000 11.330000 16.430000 ;
      RECT 11.160000 16.620000 11.330000 16.790000 ;
      RECT 11.160000 17.620000 11.330000 17.790000 ;
      RECT 11.160000 17.980000 11.330000 18.150000 ;
      RECT 11.160000 18.340000 11.330000 18.510000 ;
      RECT 11.160000 18.700000 11.330000 18.870000 ;
      RECT 11.160000 19.060000 11.330000 19.230000 ;
      RECT 11.160000 19.420000 11.330000 19.590000 ;
      RECT 11.160000 19.780000 11.330000 19.950000 ;
      RECT 11.160000 20.140000 11.330000 20.310000 ;
      RECT 11.160000 20.500000 11.330000 20.670000 ;
      RECT 11.160000 20.860000 11.330000 21.030000 ;
      RECT 11.160000 21.220000 11.330000 21.390000 ;
      RECT 11.160000 21.580000 11.330000 21.750000 ;
      RECT 11.160000 21.940000 11.330000 22.110000 ;
      RECT 11.160000 22.300000 11.330000 22.470000 ;
      RECT 11.480000  0.080000 11.650000  0.250000 ;
      RECT 11.480000 11.440000 11.650000 11.610000 ;
      RECT 11.480000 22.800000 11.650000 22.970000 ;
      RECT 11.840000  0.080000 12.010000  0.250000 ;
      RECT 11.840000 11.440000 12.010000 11.610000 ;
      RECT 11.840000 22.800000 12.010000 22.970000 ;
      RECT 12.200000  0.080000 12.370000  0.250000 ;
      RECT 12.200000 11.440000 12.370000 11.610000 ;
      RECT 12.200000 22.800000 12.370000 22.970000 ;
      RECT 12.560000  0.080000 12.730000  0.250000 ;
      RECT 12.560000 11.440000 12.730000 11.610000 ;
      RECT 12.560000 22.800000 12.730000 22.970000 ;
      RECT 12.920000  0.080000 13.090000  0.250000 ;
      RECT 12.920000 11.440000 13.090000 11.610000 ;
      RECT 12.920000 22.800000 13.090000 22.970000 ;
      RECT 13.280000  0.080000 13.450000  0.250000 ;
      RECT 13.280000 11.440000 13.450000 11.610000 ;
      RECT 13.280000 22.800000 13.450000 22.970000 ;
      RECT 13.640000  0.080000 13.810000  0.250000 ;
      RECT 13.640000 11.440000 13.810000 11.610000 ;
      RECT 13.640000 22.800000 13.810000 22.970000 ;
      RECT 14.000000  0.080000 14.170000  0.250000 ;
      RECT 14.000000 11.440000 14.170000 11.610000 ;
      RECT 14.000000 22.800000 14.170000 22.970000 ;
      RECT 14.360000  0.080000 14.530000  0.250000 ;
      RECT 14.360000 11.440000 14.530000 11.610000 ;
      RECT 14.360000 22.800000 14.530000 22.970000 ;
      RECT 14.720000  0.080000 14.890000  0.250000 ;
      RECT 14.720000 11.440000 14.890000 11.610000 ;
      RECT 14.720000 22.800000 14.890000 22.970000 ;
      RECT 15.080000  0.080000 15.250000  0.250000 ;
      RECT 15.080000 11.440000 15.250000 11.610000 ;
      RECT 15.080000 22.800000 15.250000 22.970000 ;
      RECT 15.440000  0.080000 15.610000  0.250000 ;
      RECT 15.440000 11.440000 15.610000 11.610000 ;
      RECT 15.440000 22.800000 15.610000 22.970000 ;
      RECT 15.800000  0.080000 15.970000  0.250000 ;
      RECT 15.800000 11.440000 15.970000 11.610000 ;
      RECT 15.800000 22.800000 15.970000 22.970000 ;
      RECT 16.160000  0.080000 16.330000  0.250000 ;
      RECT 16.160000 11.440000 16.330000 11.610000 ;
      RECT 16.160000 22.800000 16.330000 22.970000 ;
      RECT 16.520000  0.080000 16.690000  0.250000 ;
      RECT 16.520000 11.440000 16.690000 11.610000 ;
      RECT 16.520000 22.800000 16.690000 22.970000 ;
      RECT 16.700000  0.590000 16.870000  0.760000 ;
      RECT 16.700000  0.950000 16.870000  1.120000 ;
      RECT 16.700000  1.310000 16.870000  1.480000 ;
      RECT 16.700000  1.670000 16.870000  1.840000 ;
      RECT 16.700000  2.030000 16.870000  2.200000 ;
      RECT 16.700000  2.390000 16.870000  2.560000 ;
      RECT 16.700000  2.750000 16.870000  2.920000 ;
      RECT 16.700000  3.110000 16.870000  3.280000 ;
      RECT 16.700000  3.470000 16.870000  3.640000 ;
      RECT 16.700000  3.830000 16.870000  4.000000 ;
      RECT 16.700000  4.190000 16.870000  4.360000 ;
      RECT 16.700000  4.550000 16.870000  4.720000 ;
      RECT 16.700000  4.910000 16.870000  5.080000 ;
      RECT 16.700000  5.270000 16.870000  5.440000 ;
      RECT 16.700000  6.250000 16.870000  6.420000 ;
      RECT 16.700000  6.610000 16.870000  6.780000 ;
      RECT 16.700000  6.970000 16.870000  7.140000 ;
      RECT 16.700000  7.330000 16.870000  7.500000 ;
      RECT 16.700000  7.690000 16.870000  7.860000 ;
      RECT 16.700000  8.050000 16.870000  8.220000 ;
      RECT 16.700000  8.410000 16.870000  8.580000 ;
      RECT 16.700000  8.770000 16.870000  8.940000 ;
      RECT 16.700000  9.130000 16.870000  9.300000 ;
      RECT 16.700000  9.490000 16.870000  9.660000 ;
      RECT 16.700000  9.850000 16.870000 10.020000 ;
      RECT 16.700000 10.210000 16.870000 10.380000 ;
      RECT 16.700000 10.570000 16.870000 10.740000 ;
      RECT 16.700000 10.930000 16.870000 11.100000 ;
      RECT 16.700000 11.950000 16.870000 12.120000 ;
      RECT 16.700000 12.310000 16.870000 12.480000 ;
      RECT 16.700000 12.670000 16.870000 12.840000 ;
      RECT 16.700000 13.030000 16.870000 13.200000 ;
      RECT 16.700000 13.390000 16.870000 13.560000 ;
      RECT 16.700000 13.750000 16.870000 13.920000 ;
      RECT 16.700000 14.110000 16.870000 14.280000 ;
      RECT 16.700000 14.470000 16.870000 14.640000 ;
      RECT 16.700000 14.830000 16.870000 15.000000 ;
      RECT 16.700000 15.190000 16.870000 15.360000 ;
      RECT 16.700000 15.550000 16.870000 15.720000 ;
      RECT 16.700000 15.910000 16.870000 16.080000 ;
      RECT 16.700000 16.270000 16.870000 16.440000 ;
      RECT 16.700000 16.630000 16.870000 16.800000 ;
      RECT 16.700000 17.610000 16.870000 17.780000 ;
      RECT 16.700000 17.970000 16.870000 18.140000 ;
      RECT 16.700000 18.330000 16.870000 18.500000 ;
      RECT 16.700000 18.690000 16.870000 18.860000 ;
      RECT 16.700000 19.050000 16.870000 19.220000 ;
      RECT 16.700000 19.410000 16.870000 19.580000 ;
      RECT 16.700000 19.770000 16.870000 19.940000 ;
      RECT 16.700000 20.130000 16.870000 20.300000 ;
      RECT 16.700000 20.490000 16.870000 20.660000 ;
      RECT 16.700000 20.850000 16.870000 21.020000 ;
      RECT 16.700000 21.210000 16.870000 21.380000 ;
      RECT 16.700000 21.570000 16.870000 21.740000 ;
      RECT 16.700000 21.930000 16.870000 22.100000 ;
      RECT 16.700000 22.290000 16.870000 22.460000 ;
      RECT 16.880000  0.080000 17.050000  0.250000 ;
      RECT 16.880000 11.440000 17.050000 11.610000 ;
      RECT 16.880000 22.800000 17.050000 22.970000 ;
      RECT 17.240000  0.080000 17.410000  0.250000 ;
      RECT 17.240000 11.440000 17.410000 11.610000 ;
      RECT 17.240000 22.800000 17.410000 22.970000 ;
      RECT 17.600000  0.080000 17.770000  0.250000 ;
      RECT 17.600000 11.440000 17.770000 11.610000 ;
      RECT 17.600000 22.800000 17.770000 22.970000 ;
      RECT 17.960000  0.080000 18.130000  0.250000 ;
      RECT 17.960000 11.440000 18.130000 11.610000 ;
      RECT 17.960000 22.800000 18.130000 22.970000 ;
      RECT 18.320000  0.080000 18.490000  0.250000 ;
      RECT 18.320000 11.440000 18.490000 11.610000 ;
      RECT 18.320000 22.800000 18.490000 22.970000 ;
      RECT 18.680000  0.080000 18.850000  0.250000 ;
      RECT 18.680000 11.440000 18.850000 11.610000 ;
      RECT 18.680000 22.800000 18.850000 22.970000 ;
      RECT 19.040000  0.080000 19.210000  0.250000 ;
      RECT 19.040000 11.440000 19.210000 11.610000 ;
      RECT 19.040000 22.800000 19.210000 22.970000 ;
      RECT 19.400000  0.080000 19.570000  0.250000 ;
      RECT 19.400000 11.440000 19.570000 11.610000 ;
      RECT 19.400000 22.800000 19.570000 22.970000 ;
      RECT 19.760000  0.080000 19.930000  0.250000 ;
      RECT 19.760000 11.440000 19.930000 11.610000 ;
      RECT 19.760000 22.800000 19.930000 22.970000 ;
      RECT 20.120000  0.080000 20.290000  0.250000 ;
      RECT 20.120000 11.440000 20.290000 11.610000 ;
      RECT 20.120000 22.800000 20.290000 22.970000 ;
      RECT 20.480000  0.080000 20.650000  0.250000 ;
      RECT 20.480000 11.440000 20.650000 11.610000 ;
      RECT 20.480000 22.800000 20.650000 22.970000 ;
      RECT 20.840000  0.080000 21.010000  0.250000 ;
      RECT 20.840000 11.440000 21.010000 11.610000 ;
      RECT 20.840000 22.800000 21.010000 22.970000 ;
      RECT 21.200000  0.080000 21.370000  0.250000 ;
      RECT 21.200000 11.440000 21.370000 11.610000 ;
      RECT 21.200000 22.800000 21.370000 22.970000 ;
      RECT 21.560000  0.080000 21.730000  0.250000 ;
      RECT 21.560000 11.440000 21.730000 11.610000 ;
      RECT 21.560000 22.800000 21.730000 22.970000 ;
      RECT 21.920000  0.080000 22.090000  0.250000 ;
      RECT 21.920000 11.440000 22.090000 11.610000 ;
      RECT 21.920000 22.800000 22.090000 22.970000 ;
      RECT 22.240000  0.580000 22.410000  0.750000 ;
      RECT 22.240000  0.940000 22.410000  1.110000 ;
      RECT 22.240000  1.300000 22.410000  1.470000 ;
      RECT 22.240000  1.660000 22.410000  1.830000 ;
      RECT 22.240000  2.020000 22.410000  2.190000 ;
      RECT 22.240000  2.380000 22.410000  2.550000 ;
      RECT 22.240000  2.740000 22.410000  2.910000 ;
      RECT 22.240000  3.100000 22.410000  3.270000 ;
      RECT 22.240000  3.460000 22.410000  3.630000 ;
      RECT 22.240000  3.820000 22.410000  3.990000 ;
      RECT 22.240000  4.180000 22.410000  4.350000 ;
      RECT 22.240000  4.540000 22.410000  4.710000 ;
      RECT 22.240000  4.900000 22.410000  5.070000 ;
      RECT 22.240000  5.260000 22.410000  5.430000 ;
      RECT 22.240000  6.260000 22.410000  6.430000 ;
      RECT 22.240000  6.620000 22.410000  6.790000 ;
      RECT 22.240000  6.980000 22.410000  7.150000 ;
      RECT 22.240000  7.340000 22.410000  7.510000 ;
      RECT 22.240000  7.700000 22.410000  7.870000 ;
      RECT 22.240000  8.060000 22.410000  8.230000 ;
      RECT 22.240000  8.420000 22.410000  8.590000 ;
      RECT 22.240000  8.780000 22.410000  8.950000 ;
      RECT 22.240000  9.140000 22.410000  9.310000 ;
      RECT 22.240000  9.500000 22.410000  9.670000 ;
      RECT 22.240000  9.860000 22.410000 10.030000 ;
      RECT 22.240000 10.220000 22.410000 10.390000 ;
      RECT 22.240000 10.580000 22.410000 10.750000 ;
      RECT 22.240000 10.940000 22.410000 11.110000 ;
      RECT 22.240000 11.940000 22.410000 12.110000 ;
      RECT 22.240000 12.300000 22.410000 12.470000 ;
      RECT 22.240000 12.660000 22.410000 12.830000 ;
      RECT 22.240000 13.020000 22.410000 13.190000 ;
      RECT 22.240000 13.380000 22.410000 13.550000 ;
      RECT 22.240000 13.740000 22.410000 13.910000 ;
      RECT 22.240000 14.100000 22.410000 14.270000 ;
      RECT 22.240000 14.460000 22.410000 14.630000 ;
      RECT 22.240000 14.820000 22.410000 14.990000 ;
      RECT 22.240000 15.180000 22.410000 15.350000 ;
      RECT 22.240000 15.540000 22.410000 15.710000 ;
      RECT 22.240000 15.900000 22.410000 16.070000 ;
      RECT 22.240000 16.260000 22.410000 16.430000 ;
      RECT 22.240000 16.620000 22.410000 16.790000 ;
      RECT 22.240000 17.620000 22.410000 17.790000 ;
      RECT 22.240000 17.980000 22.410000 18.150000 ;
      RECT 22.240000 18.340000 22.410000 18.510000 ;
      RECT 22.240000 18.700000 22.410000 18.870000 ;
      RECT 22.240000 19.060000 22.410000 19.230000 ;
      RECT 22.240000 19.420000 22.410000 19.590000 ;
      RECT 22.240000 19.780000 22.410000 19.950000 ;
      RECT 22.240000 20.140000 22.410000 20.310000 ;
      RECT 22.240000 20.500000 22.410000 20.670000 ;
      RECT 22.240000 20.860000 22.410000 21.030000 ;
      RECT 22.240000 21.220000 22.410000 21.390000 ;
      RECT 22.240000 21.580000 22.410000 21.750000 ;
      RECT 22.240000 21.940000 22.410000 22.110000 ;
      RECT 22.240000 22.300000 22.410000 22.470000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 22.490000  0.330000 ;
      RECT  0.000000  0.330000  0.330000 11.360000 ;
      RECT  0.000000 11.360000 22.490000 11.690000 ;
      RECT  0.000000 11.690000  0.330000 22.720000 ;
      RECT  0.000000 22.720000 22.490000 23.050000 ;
      RECT  0.500000  0.470000  0.640000  5.685000 ;
      RECT  0.500000  5.685000 10.910000  6.005000 ;
      RECT  0.500000  6.005000  0.640000 11.220000 ;
      RECT  0.500000 11.830000  0.640000 17.045000 ;
      RECT  0.500000 17.045000 10.910000 17.365000 ;
      RECT  0.500000 17.365000  0.640000 22.580000 ;
      RECT  0.780000  0.330000  0.920000  5.545000 ;
      RECT  0.780000  6.145000  0.920000 11.360000 ;
      RECT  0.780000 11.690000  0.920000 16.905000 ;
      RECT  0.780000 17.505000  0.920000 22.720000 ;
      RECT  1.060000  0.470000  1.200000  5.685000 ;
      RECT  1.060000  6.005000  1.200000 11.220000 ;
      RECT  1.060000 11.830000  1.200000 17.045000 ;
      RECT  1.060000 17.365000  1.200000 22.580000 ;
      RECT  1.340000  0.330000  1.480000  5.545000 ;
      RECT  1.340000  6.145000  1.480000 11.360000 ;
      RECT  1.340000 11.690000  1.480000 16.905000 ;
      RECT  1.340000 17.505000  1.480000 22.720000 ;
      RECT  1.620000  0.470000  1.760000  5.685000 ;
      RECT  1.620000  6.005000  1.760000 11.220000 ;
      RECT  1.620000 11.830000  1.760000 17.045000 ;
      RECT  1.620000 17.365000  1.760000 22.580000 ;
      RECT  1.900000  0.330000  2.040000  5.545000 ;
      RECT  1.900000  6.145000  2.040000 11.360000 ;
      RECT  1.900000 11.690000  2.040000 16.905000 ;
      RECT  1.900000 17.505000  2.040000 22.720000 ;
      RECT  2.180000  0.470000  2.320000  5.685000 ;
      RECT  2.180000  6.005000  2.320000 11.220000 ;
      RECT  2.180000 11.830000  2.320000 17.045000 ;
      RECT  2.180000 17.365000  2.320000 22.580000 ;
      RECT  2.460000  0.330000  2.600000  5.545000 ;
      RECT  2.460000  6.145000  2.600000 11.360000 ;
      RECT  2.460000 11.690000  2.600000 16.905000 ;
      RECT  2.460000 17.505000  2.600000 22.720000 ;
      RECT  2.740000  0.470000  2.880000  5.685000 ;
      RECT  2.740000  6.005000  2.880000 11.220000 ;
      RECT  2.740000 11.830000  2.880000 17.045000 ;
      RECT  2.740000 17.365000  2.880000 22.580000 ;
      RECT  3.020000  0.330000  3.160000  5.545000 ;
      RECT  3.020000  6.145000  3.160000 11.360000 ;
      RECT  3.020000 11.690000  3.160000 16.905000 ;
      RECT  3.020000 17.505000  3.160000 22.720000 ;
      RECT  3.300000  0.470000  3.440000  5.685000 ;
      RECT  3.300000  6.005000  3.440000 11.220000 ;
      RECT  3.300000 11.830000  3.440000 17.045000 ;
      RECT  3.300000 17.365000  3.440000 22.580000 ;
      RECT  3.580000  0.330000  3.720000  5.545000 ;
      RECT  3.580000  6.145000  3.720000 11.360000 ;
      RECT  3.580000 11.690000  3.720000 16.905000 ;
      RECT  3.580000 17.505000  3.720000 22.720000 ;
      RECT  3.860000  0.470000  4.000000  5.685000 ;
      RECT  3.860000  6.005000  4.000000 11.220000 ;
      RECT  3.860000 11.830000  4.000000 17.045000 ;
      RECT  3.860000 17.365000  4.000000 22.580000 ;
      RECT  4.140000  0.330000  4.280000  5.545000 ;
      RECT  4.140000  6.145000  4.280000 11.360000 ;
      RECT  4.140000 11.690000  4.280000 16.905000 ;
      RECT  4.140000 17.505000  4.280000 22.720000 ;
      RECT  4.420000  0.470000  4.560000  5.685000 ;
      RECT  4.420000  6.005000  4.560000 11.220000 ;
      RECT  4.420000 11.830000  4.560000 17.045000 ;
      RECT  4.420000 17.365000  4.560000 22.580000 ;
      RECT  4.700000  0.330000  4.840000  5.545000 ;
      RECT  4.700000  6.145000  4.840000 11.360000 ;
      RECT  4.700000 11.690000  4.840000 16.905000 ;
      RECT  4.700000 17.505000  4.840000 22.720000 ;
      RECT  4.980000  0.470000  5.120000  5.685000 ;
      RECT  4.980000  6.005000  5.120000 11.220000 ;
      RECT  4.980000 11.830000  5.120000 17.045000 ;
      RECT  4.980000 17.365000  5.120000 22.580000 ;
      RECT  5.260000  0.330000  5.400000  5.545000 ;
      RECT  5.260000  6.145000  5.400000 11.360000 ;
      RECT  5.260000 11.690000  5.400000 16.905000 ;
      RECT  5.260000 17.505000  5.400000 22.720000 ;
      RECT  5.570000  0.470000  5.840000  5.685000 ;
      RECT  5.570000  6.005000  5.840000 11.220000 ;
      RECT  5.570000 11.830000  5.840000 17.045000 ;
      RECT  5.570000 17.365000  5.840000 22.580000 ;
      RECT  6.010000  0.330000  6.150000  5.545000 ;
      RECT  6.010000  6.145000  6.150000 11.360000 ;
      RECT  6.010000 11.690000  6.150000 16.905000 ;
      RECT  6.010000 17.505000  6.150000 22.720000 ;
      RECT  6.290000  0.470000  6.430000  5.685000 ;
      RECT  6.290000  6.005000  6.430000 11.220000 ;
      RECT  6.290000 11.830000  6.430000 17.045000 ;
      RECT  6.290000 17.365000  6.430000 22.580000 ;
      RECT  6.570000  0.330000  6.710000  5.545000 ;
      RECT  6.570000  6.145000  6.710000 11.360000 ;
      RECT  6.570000 11.690000  6.710000 16.905000 ;
      RECT  6.570000 17.505000  6.710000 22.720000 ;
      RECT  6.850000  0.470000  6.990000  5.685000 ;
      RECT  6.850000  6.005000  6.990000 11.220000 ;
      RECT  6.850000 11.830000  6.990000 17.045000 ;
      RECT  6.850000 17.365000  6.990000 22.580000 ;
      RECT  7.130000  0.330000  7.270000  5.545000 ;
      RECT  7.130000  6.145000  7.270000 11.360000 ;
      RECT  7.130000 11.690000  7.270000 16.905000 ;
      RECT  7.130000 17.505000  7.270000 22.720000 ;
      RECT  7.410000  0.470000  7.550000  5.685000 ;
      RECT  7.410000  6.005000  7.550000 11.220000 ;
      RECT  7.410000 11.830000  7.550000 17.045000 ;
      RECT  7.410000 17.365000  7.550000 22.580000 ;
      RECT  7.690000  0.330000  7.830000  5.545000 ;
      RECT  7.690000  6.145000  7.830000 11.360000 ;
      RECT  7.690000 11.690000  7.830000 16.905000 ;
      RECT  7.690000 17.505000  7.830000 22.720000 ;
      RECT  7.970000  0.470000  8.110000  5.685000 ;
      RECT  7.970000  6.005000  8.110000 11.220000 ;
      RECT  7.970000 11.830000  8.110000 17.045000 ;
      RECT  7.970000 17.365000  8.110000 22.580000 ;
      RECT  8.250000  0.330000  8.390000  5.545000 ;
      RECT  8.250000  6.145000  8.390000 11.360000 ;
      RECT  8.250000 11.690000  8.390000 16.905000 ;
      RECT  8.250000 17.505000  8.390000 22.720000 ;
      RECT  8.530000  0.470000  8.670000  5.685000 ;
      RECT  8.530000  6.005000  8.670000 11.220000 ;
      RECT  8.530000 11.830000  8.670000 17.045000 ;
      RECT  8.530000 17.365000  8.670000 22.580000 ;
      RECT  8.810000  0.330000  8.950000  5.545000 ;
      RECT  8.810000  6.145000  8.950000 11.360000 ;
      RECT  8.810000 11.690000  8.950000 16.905000 ;
      RECT  8.810000 17.505000  8.950000 22.720000 ;
      RECT  9.090000  0.470000  9.230000  5.685000 ;
      RECT  9.090000  6.005000  9.230000 11.220000 ;
      RECT  9.090000 11.830000  9.230000 17.045000 ;
      RECT  9.090000 17.365000  9.230000 22.580000 ;
      RECT  9.370000  0.330000  9.510000  5.545000 ;
      RECT  9.370000  6.145000  9.510000 11.360000 ;
      RECT  9.370000 11.690000  9.510000 16.905000 ;
      RECT  9.370000 17.505000  9.510000 22.720000 ;
      RECT  9.650000  0.470000  9.790000  5.685000 ;
      RECT  9.650000  6.005000  9.790000 11.220000 ;
      RECT  9.650000 11.830000  9.790000 17.045000 ;
      RECT  9.650000 17.365000  9.790000 22.580000 ;
      RECT  9.930000  0.330000 10.070000  5.545000 ;
      RECT  9.930000  6.145000 10.070000 11.360000 ;
      RECT  9.930000 11.690000 10.070000 16.905000 ;
      RECT  9.930000 17.505000 10.070000 22.720000 ;
      RECT 10.210000  0.470000 10.350000  5.685000 ;
      RECT 10.210000  6.005000 10.350000 11.220000 ;
      RECT 10.210000 11.830000 10.350000 17.045000 ;
      RECT 10.210000 17.365000 10.350000 22.580000 ;
      RECT 10.490000  0.330000 10.630000  5.545000 ;
      RECT 10.490000  6.145000 10.630000 11.360000 ;
      RECT 10.490000 11.690000 10.630000 16.905000 ;
      RECT 10.490000 17.505000 10.630000 22.720000 ;
      RECT 10.770000  0.470000 10.910000  5.685000 ;
      RECT 10.770000  6.005000 10.910000 11.220000 ;
      RECT 10.770000 11.830000 10.910000 17.045000 ;
      RECT 10.770000 17.365000 10.910000 22.580000 ;
      RECT 11.080000  0.330000 11.410000 11.360000 ;
      RECT 11.080000 11.690000 11.410000 22.720000 ;
      RECT 11.580000  0.470000 11.720000  5.685000 ;
      RECT 11.580000  5.685000 21.990000  6.005000 ;
      RECT 11.580000  6.005000 11.720000 11.220000 ;
      RECT 11.580000 11.830000 11.720000 17.045000 ;
      RECT 11.580000 17.045000 21.990000 17.365000 ;
      RECT 11.580000 17.365000 11.720000 22.580000 ;
      RECT 11.860000  0.330000 12.000000  5.545000 ;
      RECT 11.860000  6.145000 12.000000 11.360000 ;
      RECT 11.860000 11.690000 12.000000 16.905000 ;
      RECT 11.860000 17.505000 12.000000 22.720000 ;
      RECT 12.140000  0.470000 12.280000  5.685000 ;
      RECT 12.140000  6.005000 12.280000 11.220000 ;
      RECT 12.140000 11.830000 12.280000 17.045000 ;
      RECT 12.140000 17.365000 12.280000 22.580000 ;
      RECT 12.420000  0.330000 12.560000  5.545000 ;
      RECT 12.420000  6.145000 12.560000 11.360000 ;
      RECT 12.420000 11.690000 12.560000 16.905000 ;
      RECT 12.420000 17.505000 12.560000 22.720000 ;
      RECT 12.700000  0.470000 12.840000  5.685000 ;
      RECT 12.700000  6.005000 12.840000 11.220000 ;
      RECT 12.700000 11.830000 12.840000 17.045000 ;
      RECT 12.700000 17.365000 12.840000 22.580000 ;
      RECT 12.980000  0.330000 13.120000  5.545000 ;
      RECT 12.980000  6.145000 13.120000 11.360000 ;
      RECT 12.980000 11.690000 13.120000 16.905000 ;
      RECT 12.980000 17.505000 13.120000 22.720000 ;
      RECT 13.260000  0.470000 13.400000  5.685000 ;
      RECT 13.260000  6.005000 13.400000 11.220000 ;
      RECT 13.260000 11.830000 13.400000 17.045000 ;
      RECT 13.260000 17.365000 13.400000 22.580000 ;
      RECT 13.540000  0.330000 13.680000  5.545000 ;
      RECT 13.540000  6.145000 13.680000 11.360000 ;
      RECT 13.540000 11.690000 13.680000 16.905000 ;
      RECT 13.540000 17.505000 13.680000 22.720000 ;
      RECT 13.820000  0.470000 13.960000  5.685000 ;
      RECT 13.820000  6.005000 13.960000 11.220000 ;
      RECT 13.820000 11.830000 13.960000 17.045000 ;
      RECT 13.820000 17.365000 13.960000 22.580000 ;
      RECT 14.100000  0.330000 14.240000  5.545000 ;
      RECT 14.100000  6.145000 14.240000 11.360000 ;
      RECT 14.100000 11.690000 14.240000 16.905000 ;
      RECT 14.100000 17.505000 14.240000 22.720000 ;
      RECT 14.380000  0.470000 14.520000  5.685000 ;
      RECT 14.380000  6.005000 14.520000 11.220000 ;
      RECT 14.380000 11.830000 14.520000 17.045000 ;
      RECT 14.380000 17.365000 14.520000 22.580000 ;
      RECT 14.660000  0.330000 14.800000  5.545000 ;
      RECT 14.660000  6.145000 14.800000 11.360000 ;
      RECT 14.660000 11.690000 14.800000 16.905000 ;
      RECT 14.660000 17.505000 14.800000 22.720000 ;
      RECT 14.940000  0.470000 15.080000  5.685000 ;
      RECT 14.940000  6.005000 15.080000 11.220000 ;
      RECT 14.940000 11.830000 15.080000 17.045000 ;
      RECT 14.940000 17.365000 15.080000 22.580000 ;
      RECT 15.220000  0.330000 15.360000  5.545000 ;
      RECT 15.220000  6.145000 15.360000 11.360000 ;
      RECT 15.220000 11.690000 15.360000 16.905000 ;
      RECT 15.220000 17.505000 15.360000 22.720000 ;
      RECT 15.500000  0.470000 15.640000  5.685000 ;
      RECT 15.500000  6.005000 15.640000 11.220000 ;
      RECT 15.500000 11.830000 15.640000 17.045000 ;
      RECT 15.500000 17.365000 15.640000 22.580000 ;
      RECT 15.780000  0.330000 15.920000  5.545000 ;
      RECT 15.780000  6.145000 15.920000 11.360000 ;
      RECT 15.780000 11.690000 15.920000 16.905000 ;
      RECT 15.780000 17.505000 15.920000 22.720000 ;
      RECT 16.060000  0.470000 16.200000  5.685000 ;
      RECT 16.060000  6.005000 16.200000 11.220000 ;
      RECT 16.060000 11.830000 16.200000 17.045000 ;
      RECT 16.060000 17.365000 16.200000 22.580000 ;
      RECT 16.340000  0.330000 16.480000  5.545000 ;
      RECT 16.340000  6.145000 16.480000 11.360000 ;
      RECT 16.340000 11.690000 16.480000 16.905000 ;
      RECT 16.340000 17.505000 16.480000 22.720000 ;
      RECT 16.650000  0.470000 16.920000  5.685000 ;
      RECT 16.650000  6.005000 16.920000 11.220000 ;
      RECT 16.650000 11.830000 16.920000 17.045000 ;
      RECT 16.650000 17.365000 16.920000 22.580000 ;
      RECT 17.090000  0.330000 17.230000  5.545000 ;
      RECT 17.090000  6.145000 17.230000 11.360000 ;
      RECT 17.090000 11.690000 17.230000 16.905000 ;
      RECT 17.090000 17.505000 17.230000 22.720000 ;
      RECT 17.370000  0.470000 17.510000  5.685000 ;
      RECT 17.370000  6.005000 17.510000 11.220000 ;
      RECT 17.370000 11.830000 17.510000 17.045000 ;
      RECT 17.370000 17.365000 17.510000 22.580000 ;
      RECT 17.650000  0.330000 17.790000  5.545000 ;
      RECT 17.650000  6.145000 17.790000 11.360000 ;
      RECT 17.650000 11.690000 17.790000 16.905000 ;
      RECT 17.650000 17.505000 17.790000 22.720000 ;
      RECT 17.930000  0.470000 18.070000  5.685000 ;
      RECT 17.930000  6.005000 18.070000 11.220000 ;
      RECT 17.930000 11.830000 18.070000 17.045000 ;
      RECT 17.930000 17.365000 18.070000 22.580000 ;
      RECT 18.210000  0.330000 18.350000  5.545000 ;
      RECT 18.210000  6.145000 18.350000 11.360000 ;
      RECT 18.210000 11.690000 18.350000 16.905000 ;
      RECT 18.210000 17.505000 18.350000 22.720000 ;
      RECT 18.490000  0.470000 18.630000  5.685000 ;
      RECT 18.490000  6.005000 18.630000 11.220000 ;
      RECT 18.490000 11.830000 18.630000 17.045000 ;
      RECT 18.490000 17.365000 18.630000 22.580000 ;
      RECT 18.770000  0.330000 18.910000  5.545000 ;
      RECT 18.770000  6.145000 18.910000 11.360000 ;
      RECT 18.770000 11.690000 18.910000 16.905000 ;
      RECT 18.770000 17.505000 18.910000 22.720000 ;
      RECT 19.050000  0.470000 19.190000  5.685000 ;
      RECT 19.050000  6.005000 19.190000 11.220000 ;
      RECT 19.050000 11.830000 19.190000 17.045000 ;
      RECT 19.050000 17.365000 19.190000 22.580000 ;
      RECT 19.330000  0.330000 19.470000  5.545000 ;
      RECT 19.330000  6.145000 19.470000 11.360000 ;
      RECT 19.330000 11.690000 19.470000 16.905000 ;
      RECT 19.330000 17.505000 19.470000 22.720000 ;
      RECT 19.610000  0.470000 19.750000  5.685000 ;
      RECT 19.610000  6.005000 19.750000 11.220000 ;
      RECT 19.610000 11.830000 19.750000 17.045000 ;
      RECT 19.610000 17.365000 19.750000 22.580000 ;
      RECT 19.890000  0.330000 20.030000  5.545000 ;
      RECT 19.890000  6.145000 20.030000 11.360000 ;
      RECT 19.890000 11.690000 20.030000 16.905000 ;
      RECT 19.890000 17.505000 20.030000 22.720000 ;
      RECT 20.170000  0.470000 20.310000  5.685000 ;
      RECT 20.170000  6.005000 20.310000 11.220000 ;
      RECT 20.170000 11.830000 20.310000 17.045000 ;
      RECT 20.170000 17.365000 20.310000 22.580000 ;
      RECT 20.450000  0.330000 20.590000  5.545000 ;
      RECT 20.450000  6.145000 20.590000 11.360000 ;
      RECT 20.450000 11.690000 20.590000 16.905000 ;
      RECT 20.450000 17.505000 20.590000 22.720000 ;
      RECT 20.730000  0.470000 20.870000  5.685000 ;
      RECT 20.730000  6.005000 20.870000 11.220000 ;
      RECT 20.730000 11.830000 20.870000 17.045000 ;
      RECT 20.730000 17.365000 20.870000 22.580000 ;
      RECT 21.010000  0.330000 21.150000  5.545000 ;
      RECT 21.010000  6.145000 21.150000 11.360000 ;
      RECT 21.010000 11.690000 21.150000 16.905000 ;
      RECT 21.010000 17.505000 21.150000 22.720000 ;
      RECT 21.290000  0.470000 21.430000  5.685000 ;
      RECT 21.290000  6.005000 21.430000 11.220000 ;
      RECT 21.290000 11.830000 21.430000 17.045000 ;
      RECT 21.290000 17.365000 21.430000 22.580000 ;
      RECT 21.570000  0.330000 21.710000  5.545000 ;
      RECT 21.570000  6.145000 21.710000 11.360000 ;
      RECT 21.570000 11.690000 21.710000 16.905000 ;
      RECT 21.570000 17.505000 21.710000 22.720000 ;
      RECT 21.850000  0.470000 21.990000  5.685000 ;
      RECT 21.850000  6.005000 21.990000 11.220000 ;
      RECT 21.850000 11.830000 21.990000 17.045000 ;
      RECT 21.850000 17.365000 21.990000 22.580000 ;
      RECT 22.160000  0.330000 22.490000 11.360000 ;
      RECT 22.160000 11.690000 22.490000 22.720000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  5.430000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.750000 ;
      RECT  0.000000  0.750000  5.425000  0.890000 ;
      RECT  0.000000  0.890000  0.330000  1.310000 ;
      RECT  0.000000  1.310000  5.425000  1.450000 ;
      RECT  0.000000  1.450000  0.330000  1.870000 ;
      RECT  0.000000  1.870000  5.425000  2.010000 ;
      RECT  0.000000  2.010000  0.330000  2.430000 ;
      RECT  0.000000  2.430000  5.425000  2.570000 ;
      RECT  0.000000  2.570000  0.330000  2.990000 ;
      RECT  0.000000  2.990000  5.425000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.550000 ;
      RECT  0.000000  3.550000  5.425000  3.690000 ;
      RECT  0.000000  3.690000  0.330000  4.110000 ;
      RECT  0.000000  4.110000  5.425000  4.250000 ;
      RECT  0.000000  4.250000  0.330000  4.670000 ;
      RECT  0.000000  4.670000  5.425000  4.810000 ;
      RECT  0.000000  4.810000  0.330000  5.230000 ;
      RECT  0.000000  5.230000  5.425000  5.565000 ;
      RECT  0.000000  5.565000  0.330000  5.570000 ;
      RECT  0.000000  5.710000 22.490000  5.980000 ;
      RECT  0.000000  6.120000  0.330000  6.125000 ;
      RECT  0.000000  6.125000  5.425000  6.460000 ;
      RECT  0.000000  6.460000  0.330000  6.880000 ;
      RECT  0.000000  6.880000  5.425000  7.020000 ;
      RECT  0.000000  7.020000  0.330000  7.440000 ;
      RECT  0.000000  7.440000  5.425000  7.580000 ;
      RECT  0.000000  7.580000  0.330000  8.000000 ;
      RECT  0.000000  8.000000  5.425000  8.140000 ;
      RECT  0.000000  8.140000  0.330000  8.560000 ;
      RECT  0.000000  8.560000  5.425000  8.700000 ;
      RECT  0.000000  8.700000  0.330000  9.120000 ;
      RECT  0.000000  9.120000  5.425000  9.260000 ;
      RECT  0.000000  9.260000  0.330000  9.680000 ;
      RECT  0.000000  9.680000  5.425000  9.820000 ;
      RECT  0.000000  9.820000  0.330000 10.240000 ;
      RECT  0.000000 10.240000  5.425000 10.380000 ;
      RECT  0.000000 10.380000  0.330000 10.800000 ;
      RECT  0.000000 10.800000  5.425000 10.940000 ;
      RECT  0.000000 10.940000  0.330000 11.360000 ;
      RECT  0.000000 11.360000  5.430000 11.690000 ;
      RECT  0.000000 11.690000  0.330000 12.110000 ;
      RECT  0.000000 12.110000  5.425000 12.250000 ;
      RECT  0.000000 12.250000  0.330000 12.670000 ;
      RECT  0.000000 12.670000  5.425000 12.810000 ;
      RECT  0.000000 12.810000  0.330000 13.230000 ;
      RECT  0.000000 13.230000  5.425000 13.370000 ;
      RECT  0.000000 13.370000  0.330000 13.790000 ;
      RECT  0.000000 13.790000  5.425000 13.930000 ;
      RECT  0.000000 13.930000  0.330000 14.350000 ;
      RECT  0.000000 14.350000  5.425000 14.490000 ;
      RECT  0.000000 14.490000  0.330000 14.910000 ;
      RECT  0.000000 14.910000  5.425000 15.050000 ;
      RECT  0.000000 15.050000  0.330000 15.470000 ;
      RECT  0.000000 15.470000  5.425000 15.610000 ;
      RECT  0.000000 15.610000  0.330000 16.030000 ;
      RECT  0.000000 16.030000  5.425000 16.170000 ;
      RECT  0.000000 16.170000  0.330000 16.590000 ;
      RECT  0.000000 16.590000  5.425000 16.925000 ;
      RECT  0.000000 16.925000  0.330000 16.930000 ;
      RECT  0.000000 17.070000 22.490000 17.340000 ;
      RECT  0.000000 17.480000  0.330000 17.485000 ;
      RECT  0.000000 17.485000  5.425000 17.820000 ;
      RECT  0.000000 17.820000  0.330000 18.240000 ;
      RECT  0.000000 18.240000  5.425000 18.380000 ;
      RECT  0.000000 18.380000  0.330000 18.800000 ;
      RECT  0.000000 18.800000  5.425000 18.940000 ;
      RECT  0.000000 18.940000  0.330000 19.360000 ;
      RECT  0.000000 19.360000  5.425000 19.500000 ;
      RECT  0.000000 19.500000  0.330000 19.920000 ;
      RECT  0.000000 19.920000  5.425000 20.060000 ;
      RECT  0.000000 20.060000  0.330000 20.480000 ;
      RECT  0.000000 20.480000  5.425000 20.620000 ;
      RECT  0.000000 20.620000  0.330000 21.040000 ;
      RECT  0.000000 21.040000  5.425000 21.180000 ;
      RECT  0.000000 21.180000  0.330000 21.600000 ;
      RECT  0.000000 21.600000  5.425000 21.740000 ;
      RECT  0.000000 21.740000  0.330000 22.160000 ;
      RECT  0.000000 22.160000  5.425000 22.300000 ;
      RECT  0.000000 22.300000  0.330000 22.720000 ;
      RECT  0.000000 22.720000  5.430000 23.050000 ;
      RECT  0.370000  5.705000 11.040000  5.710000 ;
      RECT  0.370000  5.980000 11.040000  5.985000 ;
      RECT  0.370000 17.065000 11.040000 17.070000 ;
      RECT  0.370000 17.340000 11.040000 17.345000 ;
      RECT  0.470000  0.470000 10.940000  0.610000 ;
      RECT  0.470000  1.030000 10.940000  1.170000 ;
      RECT  0.470000  1.590000 10.940000  1.730000 ;
      RECT  0.470000  2.150000 10.940000  2.290000 ;
      RECT  0.470000  2.710000 10.940000  2.850000 ;
      RECT  0.470000  3.270000 10.940000  3.410000 ;
      RECT  0.470000  3.830000 10.940000  3.970000 ;
      RECT  0.470000  4.390000 10.940000  4.530000 ;
      RECT  0.470000  4.950000 10.940000  5.090000 ;
      RECT  0.470000  6.600000 10.940000  6.740000 ;
      RECT  0.470000  7.160000 10.940000  7.300000 ;
      RECT  0.470000  7.720000 10.940000  7.860000 ;
      RECT  0.470000  8.280000 10.940000  8.420000 ;
      RECT  0.470000  8.840000 10.940000  8.980000 ;
      RECT  0.470000  9.400000 10.940000  9.540000 ;
      RECT  0.470000  9.960000 10.940000 10.100000 ;
      RECT  0.470000 10.520000 10.940000 10.660000 ;
      RECT  0.470000 11.080000 10.940000 11.220000 ;
      RECT  0.470000 11.830000 10.940000 11.970000 ;
      RECT  0.470000 12.390000 10.940000 12.530000 ;
      RECT  0.470000 12.950000 10.940000 13.090000 ;
      RECT  0.470000 13.510000 10.940000 13.650000 ;
      RECT  0.470000 14.070000 10.940000 14.210000 ;
      RECT  0.470000 14.630000 10.940000 14.770000 ;
      RECT  0.470000 15.190000 10.940000 15.330000 ;
      RECT  0.470000 15.750000 10.940000 15.890000 ;
      RECT  0.470000 16.310000 10.940000 16.450000 ;
      RECT  0.470000 17.960000 10.940000 18.100000 ;
      RECT  0.470000 18.520000 10.940000 18.660000 ;
      RECT  0.470000 19.080000 10.940000 19.220000 ;
      RECT  0.470000 19.640000 10.940000 19.780000 ;
      RECT  0.470000 20.200000 10.940000 20.340000 ;
      RECT  0.470000 20.760000 10.940000 20.900000 ;
      RECT  0.470000 21.320000 10.940000 21.460000 ;
      RECT  0.470000 21.880000 10.940000 22.020000 ;
      RECT  0.470000 22.440000 10.940000 22.580000 ;
      RECT  5.565000  0.610000  5.845000  1.030000 ;
      RECT  5.565000  1.170000  5.845000  1.590000 ;
      RECT  5.565000  1.730000  5.845000  2.150000 ;
      RECT  5.565000  2.290000  5.845000  2.710000 ;
      RECT  5.565000  2.850000  5.845000  3.270000 ;
      RECT  5.565000  3.410000  5.845000  3.830000 ;
      RECT  5.565000  3.970000  5.845000  4.390000 ;
      RECT  5.565000  4.530000  5.845000  4.950000 ;
      RECT  5.565000  5.090000  5.845000  5.705000 ;
      RECT  5.565000  5.985000  5.845000  6.600000 ;
      RECT  5.565000  6.740000  5.845000  7.160000 ;
      RECT  5.565000  7.300000  5.845000  7.720000 ;
      RECT  5.565000  7.860000  5.845000  8.280000 ;
      RECT  5.565000  8.420000  5.845000  8.840000 ;
      RECT  5.565000  8.980000  5.845000  9.400000 ;
      RECT  5.565000  9.540000  5.845000  9.960000 ;
      RECT  5.565000 10.100000  5.845000 10.520000 ;
      RECT  5.565000 10.660000  5.845000 11.080000 ;
      RECT  5.565000 11.970000  5.845000 12.390000 ;
      RECT  5.565000 12.530000  5.845000 12.950000 ;
      RECT  5.565000 13.090000  5.845000 13.510000 ;
      RECT  5.565000 13.650000  5.845000 14.070000 ;
      RECT  5.565000 14.210000  5.845000 14.630000 ;
      RECT  5.565000 14.770000  5.845000 15.190000 ;
      RECT  5.565000 15.330000  5.845000 15.750000 ;
      RECT  5.565000 15.890000  5.845000 16.310000 ;
      RECT  5.565000 16.450000  5.845000 17.065000 ;
      RECT  5.565000 17.345000  5.845000 17.960000 ;
      RECT  5.565000 18.100000  5.845000 18.520000 ;
      RECT  5.565000 18.660000  5.845000 19.080000 ;
      RECT  5.565000 19.220000  5.845000 19.640000 ;
      RECT  5.565000 19.780000  5.845000 20.200000 ;
      RECT  5.565000 20.340000  5.845000 20.760000 ;
      RECT  5.565000 20.900000  5.845000 21.320000 ;
      RECT  5.565000 21.460000  5.845000 21.880000 ;
      RECT  5.565000 22.020000  5.845000 22.440000 ;
      RECT  5.570000  0.000000  5.840000  0.470000 ;
      RECT  5.570000 11.220000  5.840000 11.830000 ;
      RECT  5.570000 22.580000  5.840000 23.050000 ;
      RECT  5.980000  0.000000 16.510000  0.330000 ;
      RECT  5.980000 11.360000 16.510000 11.690000 ;
      RECT  5.980000 22.720000 16.510000 23.050000 ;
      RECT  5.985000  0.750000 16.505000  0.890000 ;
      RECT  5.985000  1.310000 16.505000  1.450000 ;
      RECT  5.985000  1.870000 16.505000  2.010000 ;
      RECT  5.985000  2.430000 16.505000  2.570000 ;
      RECT  5.985000  2.990000 16.505000  3.130000 ;
      RECT  5.985000  3.550000 16.505000  3.690000 ;
      RECT  5.985000  4.110000 16.505000  4.250000 ;
      RECT  5.985000  4.670000 16.505000  4.810000 ;
      RECT  5.985000  5.230000 16.505000  5.565000 ;
      RECT  5.985000  6.125000 16.505000  6.460000 ;
      RECT  5.985000  6.880000 16.505000  7.020000 ;
      RECT  5.985000  7.440000 16.505000  7.580000 ;
      RECT  5.985000  8.000000 16.505000  8.140000 ;
      RECT  5.985000  8.560000 16.505000  8.700000 ;
      RECT  5.985000  9.120000 16.505000  9.260000 ;
      RECT  5.985000  9.680000 16.505000  9.820000 ;
      RECT  5.985000 10.240000 16.505000 10.380000 ;
      RECT  5.985000 10.800000 16.505000 10.940000 ;
      RECT  5.985000 12.110000 16.505000 12.250000 ;
      RECT  5.985000 12.670000 16.505000 12.810000 ;
      RECT  5.985000 13.230000 16.505000 13.370000 ;
      RECT  5.985000 13.790000 16.505000 13.930000 ;
      RECT  5.985000 14.350000 16.505000 14.490000 ;
      RECT  5.985000 14.910000 16.505000 15.050000 ;
      RECT  5.985000 15.470000 16.505000 15.610000 ;
      RECT  5.985000 16.030000 16.505000 16.170000 ;
      RECT  5.985000 16.590000 16.505000 16.925000 ;
      RECT  5.985000 17.485000 16.505000 17.820000 ;
      RECT  5.985000 18.240000 16.505000 18.380000 ;
      RECT  5.985000 18.800000 16.505000 18.940000 ;
      RECT  5.985000 19.360000 16.505000 19.500000 ;
      RECT  5.985000 19.920000 16.505000 20.060000 ;
      RECT  5.985000 20.480000 16.505000 20.620000 ;
      RECT  5.985000 21.040000 16.505000 21.180000 ;
      RECT  5.985000 21.600000 16.505000 21.740000 ;
      RECT  5.985000 22.160000 16.505000 22.300000 ;
      RECT 11.080000  0.330000 11.410000  0.750000 ;
      RECT 11.080000  0.890000 11.410000  1.310000 ;
      RECT 11.080000  1.450000 11.410000  1.870000 ;
      RECT 11.080000  2.010000 11.410000  2.430000 ;
      RECT 11.080000  2.570000 11.410000  2.990000 ;
      RECT 11.080000  3.130000 11.410000  3.550000 ;
      RECT 11.080000  3.690000 11.410000  4.110000 ;
      RECT 11.080000  4.250000 11.410000  4.670000 ;
      RECT 11.080000  4.810000 11.410000  5.230000 ;
      RECT 11.080000  5.565000 11.410000  5.570000 ;
      RECT 11.080000  6.120000 11.410000  6.125000 ;
      RECT 11.080000  6.460000 11.410000  6.880000 ;
      RECT 11.080000  7.020000 11.410000  7.440000 ;
      RECT 11.080000  7.580000 11.410000  8.000000 ;
      RECT 11.080000  8.140000 11.410000  8.560000 ;
      RECT 11.080000  8.700000 11.410000  9.120000 ;
      RECT 11.080000  9.260000 11.410000  9.680000 ;
      RECT 11.080000  9.820000 11.410000 10.240000 ;
      RECT 11.080000 10.380000 11.410000 10.800000 ;
      RECT 11.080000 10.940000 11.410000 11.360000 ;
      RECT 11.080000 11.690000 11.410000 12.110000 ;
      RECT 11.080000 12.250000 11.410000 12.670000 ;
      RECT 11.080000 12.810000 11.410000 13.230000 ;
      RECT 11.080000 13.370000 11.410000 13.790000 ;
      RECT 11.080000 13.930000 11.410000 14.350000 ;
      RECT 11.080000 14.490000 11.410000 14.910000 ;
      RECT 11.080000 15.050000 11.410000 15.470000 ;
      RECT 11.080000 15.610000 11.410000 16.030000 ;
      RECT 11.080000 16.170000 11.410000 16.590000 ;
      RECT 11.080000 16.925000 11.410000 16.930000 ;
      RECT 11.080000 17.480000 11.410000 17.485000 ;
      RECT 11.080000 17.820000 11.410000 18.240000 ;
      RECT 11.080000 18.380000 11.410000 18.800000 ;
      RECT 11.080000 18.940000 11.410000 19.360000 ;
      RECT 11.080000 19.500000 11.410000 19.920000 ;
      RECT 11.080000 20.060000 11.410000 20.480000 ;
      RECT 11.080000 20.620000 11.410000 21.040000 ;
      RECT 11.080000 21.180000 11.410000 21.600000 ;
      RECT 11.080000 21.740000 11.410000 22.160000 ;
      RECT 11.080000 22.300000 11.410000 22.720000 ;
      RECT 11.450000  5.705000 22.120000  5.710000 ;
      RECT 11.450000  5.980000 22.120000  5.985000 ;
      RECT 11.450000 17.065000 22.120000 17.070000 ;
      RECT 11.450000 17.340000 22.120000 17.345000 ;
      RECT 11.550000  0.470000 22.020000  0.610000 ;
      RECT 11.550000  1.030000 22.020000  1.170000 ;
      RECT 11.550000  1.590000 22.020000  1.730000 ;
      RECT 11.550000  2.150000 22.020000  2.290000 ;
      RECT 11.550000  2.710000 22.020000  2.850000 ;
      RECT 11.550000  3.270000 22.020000  3.410000 ;
      RECT 11.550000  3.830000 22.020000  3.970000 ;
      RECT 11.550000  4.390000 22.020000  4.530000 ;
      RECT 11.550000  4.950000 22.020000  5.090000 ;
      RECT 11.550000  6.600000 22.020000  6.740000 ;
      RECT 11.550000  7.160000 22.020000  7.300000 ;
      RECT 11.550000  7.720000 22.020000  7.860000 ;
      RECT 11.550000  8.280000 22.020000  8.420000 ;
      RECT 11.550000  8.840000 22.020000  8.980000 ;
      RECT 11.550000  9.400000 22.020000  9.540000 ;
      RECT 11.550000  9.960000 22.020000 10.100000 ;
      RECT 11.550000 10.520000 22.020000 10.660000 ;
      RECT 11.550000 11.080000 22.020000 11.220000 ;
      RECT 11.550000 11.830000 22.020000 11.970000 ;
      RECT 11.550000 12.390000 22.020000 12.530000 ;
      RECT 11.550000 12.950000 22.020000 13.090000 ;
      RECT 11.550000 13.510000 22.020000 13.650000 ;
      RECT 11.550000 14.070000 22.020000 14.210000 ;
      RECT 11.550000 14.630000 22.020000 14.770000 ;
      RECT 11.550000 15.190000 22.020000 15.330000 ;
      RECT 11.550000 15.750000 22.020000 15.890000 ;
      RECT 11.550000 16.310000 22.020000 16.450000 ;
      RECT 11.550000 17.960000 22.020000 18.100000 ;
      RECT 11.550000 18.520000 22.020000 18.660000 ;
      RECT 11.550000 19.080000 22.020000 19.220000 ;
      RECT 11.550000 19.640000 22.020000 19.780000 ;
      RECT 11.550000 20.200000 22.020000 20.340000 ;
      RECT 11.550000 20.760000 22.020000 20.900000 ;
      RECT 11.550000 21.320000 22.020000 21.460000 ;
      RECT 11.550000 21.880000 22.020000 22.020000 ;
      RECT 11.550000 22.440000 22.020000 22.580000 ;
      RECT 16.645000  0.610000 16.925000  1.030000 ;
      RECT 16.645000  1.170000 16.925000  1.590000 ;
      RECT 16.645000  1.730000 16.925000  2.150000 ;
      RECT 16.645000  2.290000 16.925000  2.710000 ;
      RECT 16.645000  2.850000 16.925000  3.270000 ;
      RECT 16.645000  3.410000 16.925000  3.830000 ;
      RECT 16.645000  3.970000 16.925000  4.390000 ;
      RECT 16.645000  4.530000 16.925000  4.950000 ;
      RECT 16.645000  5.090000 16.925000  5.705000 ;
      RECT 16.645000  5.985000 16.925000  6.600000 ;
      RECT 16.645000  6.740000 16.925000  7.160000 ;
      RECT 16.645000  7.300000 16.925000  7.720000 ;
      RECT 16.645000  7.860000 16.925000  8.280000 ;
      RECT 16.645000  8.420000 16.925000  8.840000 ;
      RECT 16.645000  8.980000 16.925000  9.400000 ;
      RECT 16.645000  9.540000 16.925000  9.960000 ;
      RECT 16.645000 10.100000 16.925000 10.520000 ;
      RECT 16.645000 10.660000 16.925000 11.080000 ;
      RECT 16.645000 11.970000 16.925000 12.390000 ;
      RECT 16.645000 12.530000 16.925000 12.950000 ;
      RECT 16.645000 13.090000 16.925000 13.510000 ;
      RECT 16.645000 13.650000 16.925000 14.070000 ;
      RECT 16.645000 14.210000 16.925000 14.630000 ;
      RECT 16.645000 14.770000 16.925000 15.190000 ;
      RECT 16.645000 15.330000 16.925000 15.750000 ;
      RECT 16.645000 15.890000 16.925000 16.310000 ;
      RECT 16.645000 16.450000 16.925000 17.065000 ;
      RECT 16.645000 17.345000 16.925000 17.960000 ;
      RECT 16.645000 18.100000 16.925000 18.520000 ;
      RECT 16.645000 18.660000 16.925000 19.080000 ;
      RECT 16.645000 19.220000 16.925000 19.640000 ;
      RECT 16.645000 19.780000 16.925000 20.200000 ;
      RECT 16.645000 20.340000 16.925000 20.760000 ;
      RECT 16.645000 20.900000 16.925000 21.320000 ;
      RECT 16.645000 21.460000 16.925000 21.880000 ;
      RECT 16.645000 22.020000 16.925000 22.440000 ;
      RECT 16.650000  0.000000 16.920000  0.470000 ;
      RECT 16.650000 11.220000 16.920000 11.830000 ;
      RECT 16.650000 22.580000 16.920000 23.050000 ;
      RECT 17.060000  0.000000 22.490000  0.330000 ;
      RECT 17.060000 11.360000 22.490000 11.690000 ;
      RECT 17.060000 22.720000 22.490000 23.050000 ;
      RECT 17.065000  0.750000 22.490000  0.890000 ;
      RECT 17.065000  1.310000 22.490000  1.450000 ;
      RECT 17.065000  1.870000 22.490000  2.010000 ;
      RECT 17.065000  2.430000 22.490000  2.570000 ;
      RECT 17.065000  2.990000 22.490000  3.130000 ;
      RECT 17.065000  3.550000 22.490000  3.690000 ;
      RECT 17.065000  4.110000 22.490000  4.250000 ;
      RECT 17.065000  4.670000 22.490000  4.810000 ;
      RECT 17.065000  5.230000 22.490000  5.565000 ;
      RECT 17.065000  6.125000 22.490000  6.460000 ;
      RECT 17.065000  6.880000 22.490000  7.020000 ;
      RECT 17.065000  7.440000 22.490000  7.580000 ;
      RECT 17.065000  8.000000 22.490000  8.140000 ;
      RECT 17.065000  8.560000 22.490000  8.700000 ;
      RECT 17.065000  9.120000 22.490000  9.260000 ;
      RECT 17.065000  9.680000 22.490000  9.820000 ;
      RECT 17.065000 10.240000 22.490000 10.380000 ;
      RECT 17.065000 10.800000 22.490000 10.940000 ;
      RECT 17.065000 12.110000 22.490000 12.250000 ;
      RECT 17.065000 12.670000 22.490000 12.810000 ;
      RECT 17.065000 13.230000 22.490000 13.370000 ;
      RECT 17.065000 13.790000 22.490000 13.930000 ;
      RECT 17.065000 14.350000 22.490000 14.490000 ;
      RECT 17.065000 14.910000 22.490000 15.050000 ;
      RECT 17.065000 15.470000 22.490000 15.610000 ;
      RECT 17.065000 16.030000 22.490000 16.170000 ;
      RECT 17.065000 16.590000 22.490000 16.925000 ;
      RECT 17.065000 17.485000 22.490000 17.820000 ;
      RECT 17.065000 18.240000 22.490000 18.380000 ;
      RECT 17.065000 18.800000 22.490000 18.940000 ;
      RECT 17.065000 19.360000 22.490000 19.500000 ;
      RECT 17.065000 19.920000 22.490000 20.060000 ;
      RECT 17.065000 20.480000 22.490000 20.620000 ;
      RECT 17.065000 21.040000 22.490000 21.180000 ;
      RECT 17.065000 21.600000 22.490000 21.740000 ;
      RECT 17.065000 22.160000 22.490000 22.300000 ;
      RECT 22.160000  0.330000 22.490000  0.750000 ;
      RECT 22.160000  0.890000 22.490000  1.310000 ;
      RECT 22.160000  1.450000 22.490000  1.870000 ;
      RECT 22.160000  2.010000 22.490000  2.430000 ;
      RECT 22.160000  2.570000 22.490000  2.990000 ;
      RECT 22.160000  3.130000 22.490000  3.550000 ;
      RECT 22.160000  3.690000 22.490000  4.110000 ;
      RECT 22.160000  4.250000 22.490000  4.670000 ;
      RECT 22.160000  4.810000 22.490000  5.230000 ;
      RECT 22.160000  5.565000 22.490000  5.570000 ;
      RECT 22.160000  6.120000 22.490000  6.125000 ;
      RECT 22.160000  6.460000 22.490000  6.880000 ;
      RECT 22.160000  7.020000 22.490000  7.440000 ;
      RECT 22.160000  7.580000 22.490000  8.000000 ;
      RECT 22.160000  8.140000 22.490000  8.560000 ;
      RECT 22.160000  8.700000 22.490000  9.120000 ;
      RECT 22.160000  9.260000 22.490000  9.680000 ;
      RECT 22.160000  9.820000 22.490000 10.240000 ;
      RECT 22.160000 10.380000 22.490000 10.800000 ;
      RECT 22.160000 10.940000 22.490000 11.360000 ;
      RECT 22.160000 11.690000 22.490000 12.110000 ;
      RECT 22.160000 12.250000 22.490000 12.670000 ;
      RECT 22.160000 12.810000 22.490000 13.230000 ;
      RECT 22.160000 13.370000 22.490000 13.790000 ;
      RECT 22.160000 13.930000 22.490000 14.350000 ;
      RECT 22.160000 14.490000 22.490000 14.910000 ;
      RECT 22.160000 15.050000 22.490000 15.470000 ;
      RECT 22.160000 15.610000 22.490000 16.030000 ;
      RECT 22.160000 16.170000 22.490000 16.590000 ;
      RECT 22.160000 16.925000 22.490000 16.930000 ;
      RECT 22.160000 17.480000 22.490000 17.485000 ;
      RECT 22.160000 17.820000 22.490000 18.240000 ;
      RECT 22.160000 18.380000 22.490000 18.800000 ;
      RECT 22.160000 18.940000 22.490000 19.360000 ;
      RECT 22.160000 19.500000 22.490000 19.920000 ;
      RECT 22.160000 20.060000 22.490000 20.480000 ;
      RECT 22.160000 20.620000 22.490000 21.040000 ;
      RECT 22.160000 21.180000 22.490000 21.600000 ;
      RECT 22.160000 21.740000 22.490000 22.160000 ;
      RECT 22.160000 22.300000 22.490000 22.720000 ;
    LAYER pwell ;
      RECT  5.890000  7.080000  5.995000  7.325000 ;
      RECT  5.890000 18.440000  5.995000 18.685000 ;
      RECT 16.970000  7.080000 17.075000  7.325000 ;
      RECT 16.970000 18.440000 17.075000 18.685000 ;
    LAYER via ;
      RECT  0.035000  0.280000  0.295000  0.540000 ;
      RECT  0.035000  0.600000  0.295000  0.860000 ;
      RECT  0.035000  0.920000  0.295000  1.180000 ;
      RECT  0.035000  1.240000  0.295000  1.500000 ;
      RECT  0.035000  1.560000  0.295000  1.820000 ;
      RECT  0.035000  1.880000  0.295000  2.140000 ;
      RECT  0.035000  2.200000  0.295000  2.460000 ;
      RECT  0.035000  2.520000  0.295000  2.780000 ;
      RECT  0.035000  2.840000  0.295000  3.100000 ;
      RECT  0.035000  3.160000  0.295000  3.420000 ;
      RECT  0.035000  3.480000  0.295000  3.740000 ;
      RECT  0.035000  3.800000  0.295000  4.060000 ;
      RECT  0.035000  4.120000  0.295000  4.380000 ;
      RECT  0.035000  4.440000  0.295000  4.700000 ;
      RECT  0.035000  4.760000  0.295000  5.020000 ;
      RECT  0.035000  5.080000  0.295000  5.340000 ;
      RECT  0.035000  6.350000  0.295000  6.610000 ;
      RECT  0.035000  6.670000  0.295000  6.930000 ;
      RECT  0.035000  6.990000  0.295000  7.250000 ;
      RECT  0.035000  7.310000  0.295000  7.570000 ;
      RECT  0.035000  7.630000  0.295000  7.890000 ;
      RECT  0.035000  7.950000  0.295000  8.210000 ;
      RECT  0.035000  8.270000  0.295000  8.530000 ;
      RECT  0.035000  8.590000  0.295000  8.850000 ;
      RECT  0.035000  8.910000  0.295000  9.170000 ;
      RECT  0.035000  9.230000  0.295000  9.490000 ;
      RECT  0.035000  9.550000  0.295000  9.810000 ;
      RECT  0.035000  9.870000  0.295000 10.130000 ;
      RECT  0.035000 10.190000  0.295000 10.450000 ;
      RECT  0.035000 10.510000  0.295000 10.770000 ;
      RECT  0.035000 10.830000  0.295000 11.090000 ;
      RECT  0.035000 11.150000  0.295000 11.410000 ;
      RECT  0.035000 11.640000  0.295000 11.900000 ;
      RECT  0.035000 11.960000  0.295000 12.220000 ;
      RECT  0.035000 12.280000  0.295000 12.540000 ;
      RECT  0.035000 12.600000  0.295000 12.860000 ;
      RECT  0.035000 12.920000  0.295000 13.180000 ;
      RECT  0.035000 13.240000  0.295000 13.500000 ;
      RECT  0.035000 13.560000  0.295000 13.820000 ;
      RECT  0.035000 13.880000  0.295000 14.140000 ;
      RECT  0.035000 14.200000  0.295000 14.460000 ;
      RECT  0.035000 14.520000  0.295000 14.780000 ;
      RECT  0.035000 14.840000  0.295000 15.100000 ;
      RECT  0.035000 15.160000  0.295000 15.420000 ;
      RECT  0.035000 15.480000  0.295000 15.740000 ;
      RECT  0.035000 15.800000  0.295000 16.060000 ;
      RECT  0.035000 16.120000  0.295000 16.380000 ;
      RECT  0.035000 16.440000  0.295000 16.700000 ;
      RECT  0.035000 17.710000  0.295000 17.970000 ;
      RECT  0.035000 18.030000  0.295000 18.290000 ;
      RECT  0.035000 18.350000  0.295000 18.610000 ;
      RECT  0.035000 18.670000  0.295000 18.930000 ;
      RECT  0.035000 18.990000  0.295000 19.250000 ;
      RECT  0.035000 19.310000  0.295000 19.570000 ;
      RECT  0.035000 19.630000  0.295000 19.890000 ;
      RECT  0.035000 19.950000  0.295000 20.210000 ;
      RECT  0.035000 20.270000  0.295000 20.530000 ;
      RECT  0.035000 20.590000  0.295000 20.850000 ;
      RECT  0.035000 20.910000  0.295000 21.170000 ;
      RECT  0.035000 21.230000  0.295000 21.490000 ;
      RECT  0.035000 21.550000  0.295000 21.810000 ;
      RECT  0.035000 21.870000  0.295000 22.130000 ;
      RECT  0.035000 22.190000  0.295000 22.450000 ;
      RECT  0.035000 22.510000  0.295000 22.770000 ;
      RECT  0.440000  0.035000  0.700000  0.295000 ;
      RECT  0.440000 11.395000  0.700000 11.655000 ;
      RECT  0.440000 22.755000  0.700000 23.015000 ;
      RECT  0.760000  0.035000  1.020000  0.295000 ;
      RECT  0.760000  5.715000  1.020000  5.975000 ;
      RECT  0.760000 11.395000  1.020000 11.655000 ;
      RECT  0.760000 17.075000  1.020000 17.335000 ;
      RECT  0.760000 22.755000  1.020000 23.015000 ;
      RECT  1.080000  0.035000  1.340000  0.295000 ;
      RECT  1.080000  5.715000  1.340000  5.975000 ;
      RECT  1.080000 11.395000  1.340000 11.655000 ;
      RECT  1.080000 17.075000  1.340000 17.335000 ;
      RECT  1.080000 22.755000  1.340000 23.015000 ;
      RECT  1.400000  0.035000  1.660000  0.295000 ;
      RECT  1.400000  5.715000  1.660000  5.975000 ;
      RECT  1.400000 11.395000  1.660000 11.655000 ;
      RECT  1.400000 17.075000  1.660000 17.335000 ;
      RECT  1.400000 22.755000  1.660000 23.015000 ;
      RECT  1.720000  0.035000  1.980000  0.295000 ;
      RECT  1.720000  5.715000  1.980000  5.975000 ;
      RECT  1.720000 11.395000  1.980000 11.655000 ;
      RECT  1.720000 17.075000  1.980000 17.335000 ;
      RECT  1.720000 22.755000  1.980000 23.015000 ;
      RECT  2.040000  0.035000  2.300000  0.295000 ;
      RECT  2.040000  5.715000  2.300000  5.975000 ;
      RECT  2.040000 11.395000  2.300000 11.655000 ;
      RECT  2.040000 17.075000  2.300000 17.335000 ;
      RECT  2.040000 22.755000  2.300000 23.015000 ;
      RECT  2.360000  0.035000  2.620000  0.295000 ;
      RECT  2.360000  5.715000  2.620000  5.975000 ;
      RECT  2.360000 11.395000  2.620000 11.655000 ;
      RECT  2.360000 17.075000  2.620000 17.335000 ;
      RECT  2.360000 22.755000  2.620000 23.015000 ;
      RECT  2.680000  0.035000  2.940000  0.295000 ;
      RECT  2.680000  5.715000  2.940000  5.975000 ;
      RECT  2.680000 11.395000  2.940000 11.655000 ;
      RECT  2.680000 17.075000  2.940000 17.335000 ;
      RECT  2.680000 22.755000  2.940000 23.015000 ;
      RECT  3.000000  0.035000  3.260000  0.295000 ;
      RECT  3.000000  5.715000  3.260000  5.975000 ;
      RECT  3.000000 11.395000  3.260000 11.655000 ;
      RECT  3.000000 17.075000  3.260000 17.335000 ;
      RECT  3.000000 22.755000  3.260000 23.015000 ;
      RECT  3.320000  0.035000  3.580000  0.295000 ;
      RECT  3.320000  5.715000  3.580000  5.975000 ;
      RECT  3.320000 11.395000  3.580000 11.655000 ;
      RECT  3.320000 17.075000  3.580000 17.335000 ;
      RECT  3.320000 22.755000  3.580000 23.015000 ;
      RECT  3.640000  0.035000  3.900000  0.295000 ;
      RECT  3.640000  5.715000  3.900000  5.975000 ;
      RECT  3.640000 11.395000  3.900000 11.655000 ;
      RECT  3.640000 17.075000  3.900000 17.335000 ;
      RECT  3.640000 22.755000  3.900000 23.015000 ;
      RECT  3.960000  0.035000  4.220000  0.295000 ;
      RECT  3.960000  5.715000  4.220000  5.975000 ;
      RECT  3.960000 11.395000  4.220000 11.655000 ;
      RECT  3.960000 17.075000  4.220000 17.335000 ;
      RECT  3.960000 22.755000  4.220000 23.015000 ;
      RECT  4.280000  0.035000  4.540000  0.295000 ;
      RECT  4.280000  5.715000  4.540000  5.975000 ;
      RECT  4.280000 11.395000  4.540000 11.655000 ;
      RECT  4.280000 17.075000  4.540000 17.335000 ;
      RECT  4.280000 22.755000  4.540000 23.015000 ;
      RECT  4.600000  0.035000  4.860000  0.295000 ;
      RECT  4.600000  5.715000  4.860000  5.975000 ;
      RECT  4.600000 11.395000  4.860000 11.655000 ;
      RECT  4.600000 17.075000  4.860000 17.335000 ;
      RECT  4.600000 22.755000  4.860000 23.015000 ;
      RECT  4.920000  0.035000  5.180000  0.295000 ;
      RECT  4.920000  5.715000  5.180000  5.975000 ;
      RECT  4.920000 11.395000  5.180000 11.655000 ;
      RECT  4.920000 17.075000  5.180000 17.335000 ;
      RECT  4.920000 22.755000  5.180000 23.015000 ;
      RECT  5.240000  5.715000  5.500000  5.975000 ;
      RECT  5.240000 17.075000  5.500000 17.335000 ;
      RECT  5.575000  0.505000  5.835000  0.765000 ;
      RECT  5.575000  0.825000  5.835000  1.085000 ;
      RECT  5.575000  1.145000  5.835000  1.405000 ;
      RECT  5.575000  1.465000  5.835000  1.725000 ;
      RECT  5.575000  1.785000  5.835000  2.045000 ;
      RECT  5.575000  2.105000  5.835000  2.365000 ;
      RECT  5.575000  2.425000  5.835000  2.685000 ;
      RECT  5.575000  2.745000  5.835000  3.005000 ;
      RECT  5.575000  3.065000  5.835000  3.325000 ;
      RECT  5.575000  3.385000  5.835000  3.645000 ;
      RECT  5.575000  3.705000  5.835000  3.965000 ;
      RECT  5.575000  4.025000  5.835000  4.285000 ;
      RECT  5.575000  4.345000  5.835000  4.605000 ;
      RECT  5.575000  4.665000  5.835000  4.925000 ;
      RECT  5.575000  4.985000  5.835000  5.245000 ;
      RECT  5.575000  5.305000  5.835000  5.565000 ;
      RECT  5.575000  6.125000  5.835000  6.385000 ;
      RECT  5.575000  6.445000  5.835000  6.705000 ;
      RECT  5.575000  6.765000  5.835000  7.025000 ;
      RECT  5.575000  7.085000  5.835000  7.345000 ;
      RECT  5.575000  7.405000  5.835000  7.665000 ;
      RECT  5.575000  7.725000  5.835000  7.985000 ;
      RECT  5.575000  8.045000  5.835000  8.305000 ;
      RECT  5.575000  8.365000  5.835000  8.625000 ;
      RECT  5.575000  8.685000  5.835000  8.945000 ;
      RECT  5.575000  9.005000  5.835000  9.265000 ;
      RECT  5.575000  9.325000  5.835000  9.585000 ;
      RECT  5.575000  9.645000  5.835000  9.905000 ;
      RECT  5.575000  9.965000  5.835000 10.225000 ;
      RECT  5.575000 10.285000  5.835000 10.545000 ;
      RECT  5.575000 10.605000  5.835000 10.865000 ;
      RECT  5.575000 10.925000  5.835000 11.185000 ;
      RECT  5.575000 11.865000  5.835000 12.125000 ;
      RECT  5.575000 12.185000  5.835000 12.445000 ;
      RECT  5.575000 12.505000  5.835000 12.765000 ;
      RECT  5.575000 12.825000  5.835000 13.085000 ;
      RECT  5.575000 13.145000  5.835000 13.405000 ;
      RECT  5.575000 13.465000  5.835000 13.725000 ;
      RECT  5.575000 13.785000  5.835000 14.045000 ;
      RECT  5.575000 14.105000  5.835000 14.365000 ;
      RECT  5.575000 14.425000  5.835000 14.685000 ;
      RECT  5.575000 14.745000  5.835000 15.005000 ;
      RECT  5.575000 15.065000  5.835000 15.325000 ;
      RECT  5.575000 15.385000  5.835000 15.645000 ;
      RECT  5.575000 15.705000  5.835000 15.965000 ;
      RECT  5.575000 16.025000  5.835000 16.285000 ;
      RECT  5.575000 16.345000  5.835000 16.605000 ;
      RECT  5.575000 16.665000  5.835000 16.925000 ;
      RECT  5.575000 17.485000  5.835000 17.745000 ;
      RECT  5.575000 17.805000  5.835000 18.065000 ;
      RECT  5.575000 18.125000  5.835000 18.385000 ;
      RECT  5.575000 18.445000  5.835000 18.705000 ;
      RECT  5.575000 18.765000  5.835000 19.025000 ;
      RECT  5.575000 19.085000  5.835000 19.345000 ;
      RECT  5.575000 19.405000  5.835000 19.665000 ;
      RECT  5.575000 19.725000  5.835000 19.985000 ;
      RECT  5.575000 20.045000  5.835000 20.305000 ;
      RECT  5.575000 20.365000  5.835000 20.625000 ;
      RECT  5.575000 20.685000  5.835000 20.945000 ;
      RECT  5.575000 21.005000  5.835000 21.265000 ;
      RECT  5.575000 21.325000  5.835000 21.585000 ;
      RECT  5.575000 21.645000  5.835000 21.905000 ;
      RECT  5.575000 21.965000  5.835000 22.225000 ;
      RECT  5.575000 22.285000  5.835000 22.545000 ;
      RECT  5.910000  5.715000  6.170000  5.975000 ;
      RECT  5.910000 17.075000  6.170000 17.335000 ;
      RECT  6.230000  0.035000  6.490000  0.295000 ;
      RECT  6.230000  5.715000  6.490000  5.975000 ;
      RECT  6.230000 11.395000  6.490000 11.655000 ;
      RECT  6.230000 17.075000  6.490000 17.335000 ;
      RECT  6.230000 22.755000  6.490000 23.015000 ;
      RECT  6.550000  0.035000  6.810000  0.295000 ;
      RECT  6.550000  5.715000  6.810000  5.975000 ;
      RECT  6.550000 11.395000  6.810000 11.655000 ;
      RECT  6.550000 17.075000  6.810000 17.335000 ;
      RECT  6.550000 22.755000  6.810000 23.015000 ;
      RECT  6.870000  0.035000  7.130000  0.295000 ;
      RECT  6.870000  5.715000  7.130000  5.975000 ;
      RECT  6.870000 11.395000  7.130000 11.655000 ;
      RECT  6.870000 17.075000  7.130000 17.335000 ;
      RECT  6.870000 22.755000  7.130000 23.015000 ;
      RECT  7.190000  0.035000  7.450000  0.295000 ;
      RECT  7.190000  5.715000  7.450000  5.975000 ;
      RECT  7.190000 11.395000  7.450000 11.655000 ;
      RECT  7.190000 17.075000  7.450000 17.335000 ;
      RECT  7.190000 22.755000  7.450000 23.015000 ;
      RECT  7.510000  0.035000  7.770000  0.295000 ;
      RECT  7.510000  5.715000  7.770000  5.975000 ;
      RECT  7.510000 11.395000  7.770000 11.655000 ;
      RECT  7.510000 17.075000  7.770000 17.335000 ;
      RECT  7.510000 22.755000  7.770000 23.015000 ;
      RECT  7.830000  0.035000  8.090000  0.295000 ;
      RECT  7.830000  5.715000  8.090000  5.975000 ;
      RECT  7.830000 11.395000  8.090000 11.655000 ;
      RECT  7.830000 17.075000  8.090000 17.335000 ;
      RECT  7.830000 22.755000  8.090000 23.015000 ;
      RECT  8.150000  0.035000  8.410000  0.295000 ;
      RECT  8.150000  5.715000  8.410000  5.975000 ;
      RECT  8.150000 11.395000  8.410000 11.655000 ;
      RECT  8.150000 17.075000  8.410000 17.335000 ;
      RECT  8.150000 22.755000  8.410000 23.015000 ;
      RECT  8.470000  0.035000  8.730000  0.295000 ;
      RECT  8.470000  5.715000  8.730000  5.975000 ;
      RECT  8.470000 11.395000  8.730000 11.655000 ;
      RECT  8.470000 17.075000  8.730000 17.335000 ;
      RECT  8.470000 22.755000  8.730000 23.015000 ;
      RECT  8.790000  0.035000  9.050000  0.295000 ;
      RECT  8.790000  5.715000  9.050000  5.975000 ;
      RECT  8.790000 11.395000  9.050000 11.655000 ;
      RECT  8.790000 17.075000  9.050000 17.335000 ;
      RECT  8.790000 22.755000  9.050000 23.015000 ;
      RECT  9.110000  0.035000  9.370000  0.295000 ;
      RECT  9.110000  5.715000  9.370000  5.975000 ;
      RECT  9.110000 11.395000  9.370000 11.655000 ;
      RECT  9.110000 17.075000  9.370000 17.335000 ;
      RECT  9.110000 22.755000  9.370000 23.015000 ;
      RECT  9.430000  0.035000  9.690000  0.295000 ;
      RECT  9.430000  5.715000  9.690000  5.975000 ;
      RECT  9.430000 11.395000  9.690000 11.655000 ;
      RECT  9.430000 17.075000  9.690000 17.335000 ;
      RECT  9.430000 22.755000  9.690000 23.015000 ;
      RECT  9.750000  0.035000 10.010000  0.295000 ;
      RECT  9.750000  5.715000 10.010000  5.975000 ;
      RECT  9.750000 11.395000 10.010000 11.655000 ;
      RECT  9.750000 17.075000 10.010000 17.335000 ;
      RECT  9.750000 22.755000 10.010000 23.015000 ;
      RECT 10.070000  0.035000 10.330000  0.295000 ;
      RECT 10.070000  5.715000 10.330000  5.975000 ;
      RECT 10.070000 11.395000 10.330000 11.655000 ;
      RECT 10.070000 17.075000 10.330000 17.335000 ;
      RECT 10.070000 22.755000 10.330000 23.015000 ;
      RECT 10.390000  0.035000 10.650000  0.295000 ;
      RECT 10.390000  5.715000 10.650000  5.975000 ;
      RECT 10.390000 11.395000 10.650000 11.655000 ;
      RECT 10.390000 17.075000 10.650000 17.335000 ;
      RECT 10.390000 22.755000 10.650000 23.015000 ;
      RECT 10.710000  0.035000 10.970000  0.295000 ;
      RECT 10.710000 11.395000 10.970000 11.655000 ;
      RECT 10.710000 22.755000 10.970000 23.015000 ;
      RECT 11.115000  0.280000 11.375000  0.540000 ;
      RECT 11.115000  0.600000 11.375000  0.860000 ;
      RECT 11.115000  0.920000 11.375000  1.180000 ;
      RECT 11.115000  1.240000 11.375000  1.500000 ;
      RECT 11.115000  1.560000 11.375000  1.820000 ;
      RECT 11.115000  1.880000 11.375000  2.140000 ;
      RECT 11.115000  2.200000 11.375000  2.460000 ;
      RECT 11.115000  2.520000 11.375000  2.780000 ;
      RECT 11.115000  2.840000 11.375000  3.100000 ;
      RECT 11.115000  3.160000 11.375000  3.420000 ;
      RECT 11.115000  3.480000 11.375000  3.740000 ;
      RECT 11.115000  3.800000 11.375000  4.060000 ;
      RECT 11.115000  4.120000 11.375000  4.380000 ;
      RECT 11.115000  4.440000 11.375000  4.700000 ;
      RECT 11.115000  4.760000 11.375000  5.020000 ;
      RECT 11.115000  5.080000 11.375000  5.340000 ;
      RECT 11.115000  6.350000 11.375000  6.610000 ;
      RECT 11.115000  6.670000 11.375000  6.930000 ;
      RECT 11.115000  6.990000 11.375000  7.250000 ;
      RECT 11.115000  7.310000 11.375000  7.570000 ;
      RECT 11.115000  7.630000 11.375000  7.890000 ;
      RECT 11.115000  7.950000 11.375000  8.210000 ;
      RECT 11.115000  8.270000 11.375000  8.530000 ;
      RECT 11.115000  8.590000 11.375000  8.850000 ;
      RECT 11.115000  8.910000 11.375000  9.170000 ;
      RECT 11.115000  9.230000 11.375000  9.490000 ;
      RECT 11.115000  9.550000 11.375000  9.810000 ;
      RECT 11.115000  9.870000 11.375000 10.130000 ;
      RECT 11.115000 10.190000 11.375000 10.450000 ;
      RECT 11.115000 10.510000 11.375000 10.770000 ;
      RECT 11.115000 10.830000 11.375000 11.090000 ;
      RECT 11.115000 11.150000 11.375000 11.410000 ;
      RECT 11.115000 11.640000 11.375000 11.900000 ;
      RECT 11.115000 11.960000 11.375000 12.220000 ;
      RECT 11.115000 12.280000 11.375000 12.540000 ;
      RECT 11.115000 12.600000 11.375000 12.860000 ;
      RECT 11.115000 12.920000 11.375000 13.180000 ;
      RECT 11.115000 13.240000 11.375000 13.500000 ;
      RECT 11.115000 13.560000 11.375000 13.820000 ;
      RECT 11.115000 13.880000 11.375000 14.140000 ;
      RECT 11.115000 14.200000 11.375000 14.460000 ;
      RECT 11.115000 14.520000 11.375000 14.780000 ;
      RECT 11.115000 14.840000 11.375000 15.100000 ;
      RECT 11.115000 15.160000 11.375000 15.420000 ;
      RECT 11.115000 15.480000 11.375000 15.740000 ;
      RECT 11.115000 15.800000 11.375000 16.060000 ;
      RECT 11.115000 16.120000 11.375000 16.380000 ;
      RECT 11.115000 16.440000 11.375000 16.700000 ;
      RECT 11.115000 17.710000 11.375000 17.970000 ;
      RECT 11.115000 18.030000 11.375000 18.290000 ;
      RECT 11.115000 18.350000 11.375000 18.610000 ;
      RECT 11.115000 18.670000 11.375000 18.930000 ;
      RECT 11.115000 18.990000 11.375000 19.250000 ;
      RECT 11.115000 19.310000 11.375000 19.570000 ;
      RECT 11.115000 19.630000 11.375000 19.890000 ;
      RECT 11.115000 19.950000 11.375000 20.210000 ;
      RECT 11.115000 20.270000 11.375000 20.530000 ;
      RECT 11.115000 20.590000 11.375000 20.850000 ;
      RECT 11.115000 20.910000 11.375000 21.170000 ;
      RECT 11.115000 21.230000 11.375000 21.490000 ;
      RECT 11.115000 21.550000 11.375000 21.810000 ;
      RECT 11.115000 21.870000 11.375000 22.130000 ;
      RECT 11.115000 22.190000 11.375000 22.450000 ;
      RECT 11.115000 22.510000 11.375000 22.770000 ;
      RECT 11.520000  0.035000 11.780000  0.295000 ;
      RECT 11.520000 11.395000 11.780000 11.655000 ;
      RECT 11.520000 22.755000 11.780000 23.015000 ;
      RECT 11.840000  0.035000 12.100000  0.295000 ;
      RECT 11.840000  5.715000 12.100000  5.975000 ;
      RECT 11.840000 11.395000 12.100000 11.655000 ;
      RECT 11.840000 17.075000 12.100000 17.335000 ;
      RECT 11.840000 22.755000 12.100000 23.015000 ;
      RECT 12.160000  0.035000 12.420000  0.295000 ;
      RECT 12.160000  5.715000 12.420000  5.975000 ;
      RECT 12.160000 11.395000 12.420000 11.655000 ;
      RECT 12.160000 17.075000 12.420000 17.335000 ;
      RECT 12.160000 22.755000 12.420000 23.015000 ;
      RECT 12.480000  0.035000 12.740000  0.295000 ;
      RECT 12.480000  5.715000 12.740000  5.975000 ;
      RECT 12.480000 11.395000 12.740000 11.655000 ;
      RECT 12.480000 17.075000 12.740000 17.335000 ;
      RECT 12.480000 22.755000 12.740000 23.015000 ;
      RECT 12.800000  0.035000 13.060000  0.295000 ;
      RECT 12.800000  5.715000 13.060000  5.975000 ;
      RECT 12.800000 11.395000 13.060000 11.655000 ;
      RECT 12.800000 17.075000 13.060000 17.335000 ;
      RECT 12.800000 22.755000 13.060000 23.015000 ;
      RECT 13.120000  0.035000 13.380000  0.295000 ;
      RECT 13.120000  5.715000 13.380000  5.975000 ;
      RECT 13.120000 11.395000 13.380000 11.655000 ;
      RECT 13.120000 17.075000 13.380000 17.335000 ;
      RECT 13.120000 22.755000 13.380000 23.015000 ;
      RECT 13.440000  0.035000 13.700000  0.295000 ;
      RECT 13.440000  5.715000 13.700000  5.975000 ;
      RECT 13.440000 11.395000 13.700000 11.655000 ;
      RECT 13.440000 17.075000 13.700000 17.335000 ;
      RECT 13.440000 22.755000 13.700000 23.015000 ;
      RECT 13.760000  0.035000 14.020000  0.295000 ;
      RECT 13.760000  5.715000 14.020000  5.975000 ;
      RECT 13.760000 11.395000 14.020000 11.655000 ;
      RECT 13.760000 17.075000 14.020000 17.335000 ;
      RECT 13.760000 22.755000 14.020000 23.015000 ;
      RECT 14.080000  0.035000 14.340000  0.295000 ;
      RECT 14.080000  5.715000 14.340000  5.975000 ;
      RECT 14.080000 11.395000 14.340000 11.655000 ;
      RECT 14.080000 17.075000 14.340000 17.335000 ;
      RECT 14.080000 22.755000 14.340000 23.015000 ;
      RECT 14.400000  0.035000 14.660000  0.295000 ;
      RECT 14.400000  5.715000 14.660000  5.975000 ;
      RECT 14.400000 11.395000 14.660000 11.655000 ;
      RECT 14.400000 17.075000 14.660000 17.335000 ;
      RECT 14.400000 22.755000 14.660000 23.015000 ;
      RECT 14.720000  0.035000 14.980000  0.295000 ;
      RECT 14.720000  5.715000 14.980000  5.975000 ;
      RECT 14.720000 11.395000 14.980000 11.655000 ;
      RECT 14.720000 17.075000 14.980000 17.335000 ;
      RECT 14.720000 22.755000 14.980000 23.015000 ;
      RECT 15.040000  0.035000 15.300000  0.295000 ;
      RECT 15.040000  5.715000 15.300000  5.975000 ;
      RECT 15.040000 11.395000 15.300000 11.655000 ;
      RECT 15.040000 17.075000 15.300000 17.335000 ;
      RECT 15.040000 22.755000 15.300000 23.015000 ;
      RECT 15.360000  0.035000 15.620000  0.295000 ;
      RECT 15.360000  5.715000 15.620000  5.975000 ;
      RECT 15.360000 11.395000 15.620000 11.655000 ;
      RECT 15.360000 17.075000 15.620000 17.335000 ;
      RECT 15.360000 22.755000 15.620000 23.015000 ;
      RECT 15.680000  0.035000 15.940000  0.295000 ;
      RECT 15.680000  5.715000 15.940000  5.975000 ;
      RECT 15.680000 11.395000 15.940000 11.655000 ;
      RECT 15.680000 17.075000 15.940000 17.335000 ;
      RECT 15.680000 22.755000 15.940000 23.015000 ;
      RECT 16.000000  0.035000 16.260000  0.295000 ;
      RECT 16.000000  5.715000 16.260000  5.975000 ;
      RECT 16.000000 11.395000 16.260000 11.655000 ;
      RECT 16.000000 17.075000 16.260000 17.335000 ;
      RECT 16.000000 22.755000 16.260000 23.015000 ;
      RECT 16.320000  5.715000 16.580000  5.975000 ;
      RECT 16.320000 17.075000 16.580000 17.335000 ;
      RECT 16.655000  0.505000 16.915000  0.765000 ;
      RECT 16.655000  0.825000 16.915000  1.085000 ;
      RECT 16.655000  1.145000 16.915000  1.405000 ;
      RECT 16.655000  1.465000 16.915000  1.725000 ;
      RECT 16.655000  1.785000 16.915000  2.045000 ;
      RECT 16.655000  2.105000 16.915000  2.365000 ;
      RECT 16.655000  2.425000 16.915000  2.685000 ;
      RECT 16.655000  2.745000 16.915000  3.005000 ;
      RECT 16.655000  3.065000 16.915000  3.325000 ;
      RECT 16.655000  3.385000 16.915000  3.645000 ;
      RECT 16.655000  3.705000 16.915000  3.965000 ;
      RECT 16.655000  4.025000 16.915000  4.285000 ;
      RECT 16.655000  4.345000 16.915000  4.605000 ;
      RECT 16.655000  4.665000 16.915000  4.925000 ;
      RECT 16.655000  4.985000 16.915000  5.245000 ;
      RECT 16.655000  5.305000 16.915000  5.565000 ;
      RECT 16.655000  6.125000 16.915000  6.385000 ;
      RECT 16.655000  6.445000 16.915000  6.705000 ;
      RECT 16.655000  6.765000 16.915000  7.025000 ;
      RECT 16.655000  7.085000 16.915000  7.345000 ;
      RECT 16.655000  7.405000 16.915000  7.665000 ;
      RECT 16.655000  7.725000 16.915000  7.985000 ;
      RECT 16.655000  8.045000 16.915000  8.305000 ;
      RECT 16.655000  8.365000 16.915000  8.625000 ;
      RECT 16.655000  8.685000 16.915000  8.945000 ;
      RECT 16.655000  9.005000 16.915000  9.265000 ;
      RECT 16.655000  9.325000 16.915000  9.585000 ;
      RECT 16.655000  9.645000 16.915000  9.905000 ;
      RECT 16.655000  9.965000 16.915000 10.225000 ;
      RECT 16.655000 10.285000 16.915000 10.545000 ;
      RECT 16.655000 10.605000 16.915000 10.865000 ;
      RECT 16.655000 10.925000 16.915000 11.185000 ;
      RECT 16.655000 11.865000 16.915000 12.125000 ;
      RECT 16.655000 12.185000 16.915000 12.445000 ;
      RECT 16.655000 12.505000 16.915000 12.765000 ;
      RECT 16.655000 12.825000 16.915000 13.085000 ;
      RECT 16.655000 13.145000 16.915000 13.405000 ;
      RECT 16.655000 13.465000 16.915000 13.725000 ;
      RECT 16.655000 13.785000 16.915000 14.045000 ;
      RECT 16.655000 14.105000 16.915000 14.365000 ;
      RECT 16.655000 14.425000 16.915000 14.685000 ;
      RECT 16.655000 14.745000 16.915000 15.005000 ;
      RECT 16.655000 15.065000 16.915000 15.325000 ;
      RECT 16.655000 15.385000 16.915000 15.645000 ;
      RECT 16.655000 15.705000 16.915000 15.965000 ;
      RECT 16.655000 16.025000 16.915000 16.285000 ;
      RECT 16.655000 16.345000 16.915000 16.605000 ;
      RECT 16.655000 16.665000 16.915000 16.925000 ;
      RECT 16.655000 17.485000 16.915000 17.745000 ;
      RECT 16.655000 17.805000 16.915000 18.065000 ;
      RECT 16.655000 18.125000 16.915000 18.385000 ;
      RECT 16.655000 18.445000 16.915000 18.705000 ;
      RECT 16.655000 18.765000 16.915000 19.025000 ;
      RECT 16.655000 19.085000 16.915000 19.345000 ;
      RECT 16.655000 19.405000 16.915000 19.665000 ;
      RECT 16.655000 19.725000 16.915000 19.985000 ;
      RECT 16.655000 20.045000 16.915000 20.305000 ;
      RECT 16.655000 20.365000 16.915000 20.625000 ;
      RECT 16.655000 20.685000 16.915000 20.945000 ;
      RECT 16.655000 21.005000 16.915000 21.265000 ;
      RECT 16.655000 21.325000 16.915000 21.585000 ;
      RECT 16.655000 21.645000 16.915000 21.905000 ;
      RECT 16.655000 21.965000 16.915000 22.225000 ;
      RECT 16.655000 22.285000 16.915000 22.545000 ;
      RECT 16.990000  5.715000 17.250000  5.975000 ;
      RECT 16.990000 17.075000 17.250000 17.335000 ;
      RECT 17.310000  0.035000 17.570000  0.295000 ;
      RECT 17.310000  5.715000 17.570000  5.975000 ;
      RECT 17.310000 11.395000 17.570000 11.655000 ;
      RECT 17.310000 17.075000 17.570000 17.335000 ;
      RECT 17.310000 22.755000 17.570000 23.015000 ;
      RECT 17.630000  0.035000 17.890000  0.295000 ;
      RECT 17.630000  5.715000 17.890000  5.975000 ;
      RECT 17.630000 11.395000 17.890000 11.655000 ;
      RECT 17.630000 17.075000 17.890000 17.335000 ;
      RECT 17.630000 22.755000 17.890000 23.015000 ;
      RECT 17.950000  0.035000 18.210000  0.295000 ;
      RECT 17.950000  5.715000 18.210000  5.975000 ;
      RECT 17.950000 11.395000 18.210000 11.655000 ;
      RECT 17.950000 17.075000 18.210000 17.335000 ;
      RECT 17.950000 22.755000 18.210000 23.015000 ;
      RECT 18.270000  0.035000 18.530000  0.295000 ;
      RECT 18.270000  5.715000 18.530000  5.975000 ;
      RECT 18.270000 11.395000 18.530000 11.655000 ;
      RECT 18.270000 17.075000 18.530000 17.335000 ;
      RECT 18.270000 22.755000 18.530000 23.015000 ;
      RECT 18.590000  0.035000 18.850000  0.295000 ;
      RECT 18.590000  5.715000 18.850000  5.975000 ;
      RECT 18.590000 11.395000 18.850000 11.655000 ;
      RECT 18.590000 17.075000 18.850000 17.335000 ;
      RECT 18.590000 22.755000 18.850000 23.015000 ;
      RECT 18.910000  0.035000 19.170000  0.295000 ;
      RECT 18.910000  5.715000 19.170000  5.975000 ;
      RECT 18.910000 11.395000 19.170000 11.655000 ;
      RECT 18.910000 17.075000 19.170000 17.335000 ;
      RECT 18.910000 22.755000 19.170000 23.015000 ;
      RECT 19.230000  0.035000 19.490000  0.295000 ;
      RECT 19.230000  5.715000 19.490000  5.975000 ;
      RECT 19.230000 11.395000 19.490000 11.655000 ;
      RECT 19.230000 17.075000 19.490000 17.335000 ;
      RECT 19.230000 22.755000 19.490000 23.015000 ;
      RECT 19.550000  0.035000 19.810000  0.295000 ;
      RECT 19.550000  5.715000 19.810000  5.975000 ;
      RECT 19.550000 11.395000 19.810000 11.655000 ;
      RECT 19.550000 17.075000 19.810000 17.335000 ;
      RECT 19.550000 22.755000 19.810000 23.015000 ;
      RECT 19.870000  0.035000 20.130000  0.295000 ;
      RECT 19.870000  5.715000 20.130000  5.975000 ;
      RECT 19.870000 11.395000 20.130000 11.655000 ;
      RECT 19.870000 17.075000 20.130000 17.335000 ;
      RECT 19.870000 22.755000 20.130000 23.015000 ;
      RECT 20.190000  0.035000 20.450000  0.295000 ;
      RECT 20.190000  5.715000 20.450000  5.975000 ;
      RECT 20.190000 11.395000 20.450000 11.655000 ;
      RECT 20.190000 17.075000 20.450000 17.335000 ;
      RECT 20.190000 22.755000 20.450000 23.015000 ;
      RECT 20.510000  0.035000 20.770000  0.295000 ;
      RECT 20.510000  5.715000 20.770000  5.975000 ;
      RECT 20.510000 11.395000 20.770000 11.655000 ;
      RECT 20.510000 17.075000 20.770000 17.335000 ;
      RECT 20.510000 22.755000 20.770000 23.015000 ;
      RECT 20.830000  0.035000 21.090000  0.295000 ;
      RECT 20.830000  5.715000 21.090000  5.975000 ;
      RECT 20.830000 11.395000 21.090000 11.655000 ;
      RECT 20.830000 17.075000 21.090000 17.335000 ;
      RECT 20.830000 22.755000 21.090000 23.015000 ;
      RECT 21.150000  0.035000 21.410000  0.295000 ;
      RECT 21.150000  5.715000 21.410000  5.975000 ;
      RECT 21.150000 11.395000 21.410000 11.655000 ;
      RECT 21.150000 17.075000 21.410000 17.335000 ;
      RECT 21.150000 22.755000 21.410000 23.015000 ;
      RECT 21.470000  0.035000 21.730000  0.295000 ;
      RECT 21.470000  5.715000 21.730000  5.975000 ;
      RECT 21.470000 11.395000 21.730000 11.655000 ;
      RECT 21.470000 17.075000 21.730000 17.335000 ;
      RECT 21.470000 22.755000 21.730000 23.015000 ;
      RECT 21.790000  0.035000 22.050000  0.295000 ;
      RECT 21.790000 11.395000 22.050000 11.655000 ;
      RECT 21.790000 22.755000 22.050000 23.015000 ;
      RECT 22.195000  0.280000 22.455000  0.540000 ;
      RECT 22.195000  0.600000 22.455000  0.860000 ;
      RECT 22.195000  0.920000 22.455000  1.180000 ;
      RECT 22.195000  1.240000 22.455000  1.500000 ;
      RECT 22.195000  1.560000 22.455000  1.820000 ;
      RECT 22.195000  1.880000 22.455000  2.140000 ;
      RECT 22.195000  2.200000 22.455000  2.460000 ;
      RECT 22.195000  2.520000 22.455000  2.780000 ;
      RECT 22.195000  2.840000 22.455000  3.100000 ;
      RECT 22.195000  3.160000 22.455000  3.420000 ;
      RECT 22.195000  3.480000 22.455000  3.740000 ;
      RECT 22.195000  3.800000 22.455000  4.060000 ;
      RECT 22.195000  4.120000 22.455000  4.380000 ;
      RECT 22.195000  4.440000 22.455000  4.700000 ;
      RECT 22.195000  4.760000 22.455000  5.020000 ;
      RECT 22.195000  5.080000 22.455000  5.340000 ;
      RECT 22.195000  6.350000 22.455000  6.610000 ;
      RECT 22.195000  6.670000 22.455000  6.930000 ;
      RECT 22.195000  6.990000 22.455000  7.250000 ;
      RECT 22.195000  7.310000 22.455000  7.570000 ;
      RECT 22.195000  7.630000 22.455000  7.890000 ;
      RECT 22.195000  7.950000 22.455000  8.210000 ;
      RECT 22.195000  8.270000 22.455000  8.530000 ;
      RECT 22.195000  8.590000 22.455000  8.850000 ;
      RECT 22.195000  8.910000 22.455000  9.170000 ;
      RECT 22.195000  9.230000 22.455000  9.490000 ;
      RECT 22.195000  9.550000 22.455000  9.810000 ;
      RECT 22.195000  9.870000 22.455000 10.130000 ;
      RECT 22.195000 10.190000 22.455000 10.450000 ;
      RECT 22.195000 10.510000 22.455000 10.770000 ;
      RECT 22.195000 10.830000 22.455000 11.090000 ;
      RECT 22.195000 11.150000 22.455000 11.410000 ;
      RECT 22.195000 11.640000 22.455000 11.900000 ;
      RECT 22.195000 11.960000 22.455000 12.220000 ;
      RECT 22.195000 12.280000 22.455000 12.540000 ;
      RECT 22.195000 12.600000 22.455000 12.860000 ;
      RECT 22.195000 12.920000 22.455000 13.180000 ;
      RECT 22.195000 13.240000 22.455000 13.500000 ;
      RECT 22.195000 13.560000 22.455000 13.820000 ;
      RECT 22.195000 13.880000 22.455000 14.140000 ;
      RECT 22.195000 14.200000 22.455000 14.460000 ;
      RECT 22.195000 14.520000 22.455000 14.780000 ;
      RECT 22.195000 14.840000 22.455000 15.100000 ;
      RECT 22.195000 15.160000 22.455000 15.420000 ;
      RECT 22.195000 15.480000 22.455000 15.740000 ;
      RECT 22.195000 15.800000 22.455000 16.060000 ;
      RECT 22.195000 16.120000 22.455000 16.380000 ;
      RECT 22.195000 16.440000 22.455000 16.700000 ;
      RECT 22.195000 17.710000 22.455000 17.970000 ;
      RECT 22.195000 18.030000 22.455000 18.290000 ;
      RECT 22.195000 18.350000 22.455000 18.610000 ;
      RECT 22.195000 18.670000 22.455000 18.930000 ;
      RECT 22.195000 18.990000 22.455000 19.250000 ;
      RECT 22.195000 19.310000 22.455000 19.570000 ;
      RECT 22.195000 19.630000 22.455000 19.890000 ;
      RECT 22.195000 19.950000 22.455000 20.210000 ;
      RECT 22.195000 20.270000 22.455000 20.530000 ;
      RECT 22.195000 20.590000 22.455000 20.850000 ;
      RECT 22.195000 20.910000 22.455000 21.170000 ;
      RECT 22.195000 21.230000 22.455000 21.490000 ;
      RECT 22.195000 21.550000 22.455000 21.810000 ;
      RECT 22.195000 21.870000 22.455000 22.130000 ;
      RECT 22.195000 22.190000 22.455000 22.450000 ;
      RECT 22.195000 22.510000 22.455000 22.770000 ;
    LAYER via2 ;
      RECT  0.025000  0.445000  0.305000  0.725000 ;
      RECT  0.025000  0.845000  0.305000  1.125000 ;
      RECT  0.025000  1.245000  0.305000  1.525000 ;
      RECT  0.025000  1.645000  0.305000  1.925000 ;
      RECT  0.025000  2.045000  0.305000  2.325000 ;
      RECT  0.025000  2.445000  0.305000  2.725000 ;
      RECT  0.025000  2.845000  0.305000  3.125000 ;
      RECT  0.025000  3.245000  0.305000  3.525000 ;
      RECT  0.025000  3.645000  0.305000  3.925000 ;
      RECT  0.025000  4.045000  0.305000  4.325000 ;
      RECT  0.025000  4.445000  0.305000  4.725000 ;
      RECT  0.025000  4.845000  0.305000  5.125000 ;
      RECT  0.025000  5.245000  0.305000  5.525000 ;
      RECT  0.025000  6.165000  0.305000  6.445000 ;
      RECT  0.025000  6.565000  0.305000  6.845000 ;
      RECT  0.025000  6.965000  0.305000  7.245000 ;
      RECT  0.025000  7.365000  0.305000  7.645000 ;
      RECT  0.025000  7.765000  0.305000  8.045000 ;
      RECT  0.025000  8.165000  0.305000  8.445000 ;
      RECT  0.025000  8.565000  0.305000  8.845000 ;
      RECT  0.025000  8.965000  0.305000  9.245000 ;
      RECT  0.025000  9.365000  0.305000  9.645000 ;
      RECT  0.025000  9.765000  0.305000 10.045000 ;
      RECT  0.025000 10.165000  0.305000 10.445000 ;
      RECT  0.025000 10.565000  0.305000 10.845000 ;
      RECT  0.025000 10.965000  0.305000 11.245000 ;
      RECT  0.025000 11.805000  0.305000 12.085000 ;
      RECT  0.025000 12.205000  0.305000 12.485000 ;
      RECT  0.025000 12.605000  0.305000 12.885000 ;
      RECT  0.025000 13.005000  0.305000 13.285000 ;
      RECT  0.025000 13.405000  0.305000 13.685000 ;
      RECT  0.025000 13.805000  0.305000 14.085000 ;
      RECT  0.025000 14.205000  0.305000 14.485000 ;
      RECT  0.025000 14.605000  0.305000 14.885000 ;
      RECT  0.025000 15.005000  0.305000 15.285000 ;
      RECT  0.025000 15.405000  0.305000 15.685000 ;
      RECT  0.025000 15.805000  0.305000 16.085000 ;
      RECT  0.025000 16.205000  0.305000 16.485000 ;
      RECT  0.025000 16.605000  0.305000 16.885000 ;
      RECT  0.025000 17.525000  0.305000 17.805000 ;
      RECT  0.025000 17.925000  0.305000 18.205000 ;
      RECT  0.025000 18.325000  0.305000 18.605000 ;
      RECT  0.025000 18.725000  0.305000 19.005000 ;
      RECT  0.025000 19.125000  0.305000 19.405000 ;
      RECT  0.025000 19.525000  0.305000 19.805000 ;
      RECT  0.025000 19.925000  0.305000 20.205000 ;
      RECT  0.025000 20.325000  0.305000 20.605000 ;
      RECT  0.025000 20.725000  0.305000 21.005000 ;
      RECT  0.025000 21.125000  0.305000 21.405000 ;
      RECT  0.025000 21.525000  0.305000 21.805000 ;
      RECT  0.025000 21.925000  0.305000 22.205000 ;
      RECT  0.025000 22.325000  0.305000 22.605000 ;
      RECT  0.305000  0.025000  0.585000  0.305000 ;
      RECT  0.305000 11.385000  0.585000 11.665000 ;
      RECT  0.305000 22.745000  0.585000 23.025000 ;
      RECT  0.705000  0.025000  0.985000  0.305000 ;
      RECT  0.705000 11.385000  0.985000 11.665000 ;
      RECT  0.705000 22.745000  0.985000 23.025000 ;
      RECT  0.765000  5.705000  1.045000  5.985000 ;
      RECT  0.765000 17.065000  1.045000 17.345000 ;
      RECT  1.105000  0.025000  1.385000  0.305000 ;
      RECT  1.105000 11.385000  1.385000 11.665000 ;
      RECT  1.105000 22.745000  1.385000 23.025000 ;
      RECT  1.165000  5.705000  1.445000  5.985000 ;
      RECT  1.165000 17.065000  1.445000 17.345000 ;
      RECT  1.505000  0.025000  1.785000  0.305000 ;
      RECT  1.505000 11.385000  1.785000 11.665000 ;
      RECT  1.505000 22.745000  1.785000 23.025000 ;
      RECT  1.565000  5.705000  1.845000  5.985000 ;
      RECT  1.565000 17.065000  1.845000 17.345000 ;
      RECT  1.905000  0.025000  2.185000  0.305000 ;
      RECT  1.905000 11.385000  2.185000 11.665000 ;
      RECT  1.905000 22.745000  2.185000 23.025000 ;
      RECT  1.965000  5.705000  2.245000  5.985000 ;
      RECT  1.965000 17.065000  2.245000 17.345000 ;
      RECT  2.305000  0.025000  2.585000  0.305000 ;
      RECT  2.305000 11.385000  2.585000 11.665000 ;
      RECT  2.305000 22.745000  2.585000 23.025000 ;
      RECT  2.365000  5.705000  2.645000  5.985000 ;
      RECT  2.365000 17.065000  2.645000 17.345000 ;
      RECT  2.705000  0.025000  2.985000  0.305000 ;
      RECT  2.705000 11.385000  2.985000 11.665000 ;
      RECT  2.705000 22.745000  2.985000 23.025000 ;
      RECT  2.765000  5.705000  3.045000  5.985000 ;
      RECT  2.765000 17.065000  3.045000 17.345000 ;
      RECT  3.105000  0.025000  3.385000  0.305000 ;
      RECT  3.105000 11.385000  3.385000 11.665000 ;
      RECT  3.105000 22.745000  3.385000 23.025000 ;
      RECT  3.165000  5.705000  3.445000  5.985000 ;
      RECT  3.165000 17.065000  3.445000 17.345000 ;
      RECT  3.505000  0.025000  3.785000  0.305000 ;
      RECT  3.505000 11.385000  3.785000 11.665000 ;
      RECT  3.505000 22.745000  3.785000 23.025000 ;
      RECT  3.565000  5.705000  3.845000  5.985000 ;
      RECT  3.565000 17.065000  3.845000 17.345000 ;
      RECT  3.905000  0.025000  4.185000  0.305000 ;
      RECT  3.905000 11.385000  4.185000 11.665000 ;
      RECT  3.905000 22.745000  4.185000 23.025000 ;
      RECT  3.965000  5.705000  4.245000  5.985000 ;
      RECT  3.965000 17.065000  4.245000 17.345000 ;
      RECT  4.305000  0.025000  4.585000  0.305000 ;
      RECT  4.305000 11.385000  4.585000 11.665000 ;
      RECT  4.305000 22.745000  4.585000 23.025000 ;
      RECT  4.365000  5.705000  4.645000  5.985000 ;
      RECT  4.365000 17.065000  4.645000 17.345000 ;
      RECT  4.705000  0.025000  4.985000  0.305000 ;
      RECT  4.705000 11.385000  4.985000 11.665000 ;
      RECT  4.705000 22.745000  4.985000 23.025000 ;
      RECT  4.765000  5.705000  5.045000  5.985000 ;
      RECT  4.765000 17.065000  5.045000 17.345000 ;
      RECT  5.105000  0.025000  5.385000  0.305000 ;
      RECT  5.105000 11.385000  5.385000 11.665000 ;
      RECT  5.105000 22.745000  5.385000 23.025000 ;
      RECT  5.165000  5.705000  5.445000  5.985000 ;
      RECT  5.165000 17.065000  5.445000 17.345000 ;
      RECT  5.565000  0.905000  5.845000  1.185000 ;
      RECT  5.565000  1.305000  5.845000  1.585000 ;
      RECT  5.565000  1.705000  5.845000  1.985000 ;
      RECT  5.565000  2.105000  5.845000  2.385000 ;
      RECT  5.565000  2.505000  5.845000  2.785000 ;
      RECT  5.565000  2.905000  5.845000  3.185000 ;
      RECT  5.565000  3.305000  5.845000  3.585000 ;
      RECT  5.565000  3.705000  5.845000  3.985000 ;
      RECT  5.565000  4.105000  5.845000  4.385000 ;
      RECT  5.565000  4.505000  5.845000  4.785000 ;
      RECT  5.565000  4.905000  5.845000  5.185000 ;
      RECT  5.565000  5.305000  5.845000  5.585000 ;
      RECT  5.565000  5.705000  5.845000  5.985000 ;
      RECT  5.565000  6.105000  5.845000  6.385000 ;
      RECT  5.565000  6.505000  5.845000  6.785000 ;
      RECT  5.565000  6.905000  5.845000  7.185000 ;
      RECT  5.565000  7.305000  5.845000  7.585000 ;
      RECT  5.565000  7.705000  5.845000  7.985000 ;
      RECT  5.565000  8.105000  5.845000  8.385000 ;
      RECT  5.565000  8.505000  5.845000  8.785000 ;
      RECT  5.565000  8.905000  5.845000  9.185000 ;
      RECT  5.565000  9.305000  5.845000  9.585000 ;
      RECT  5.565000  9.705000  5.845000  9.985000 ;
      RECT  5.565000 10.105000  5.845000 10.385000 ;
      RECT  5.565000 10.505000  5.845000 10.785000 ;
      RECT  5.565000 12.265000  5.845000 12.545000 ;
      RECT  5.565000 12.665000  5.845000 12.945000 ;
      RECT  5.565000 13.065000  5.845000 13.345000 ;
      RECT  5.565000 13.465000  5.845000 13.745000 ;
      RECT  5.565000 13.865000  5.845000 14.145000 ;
      RECT  5.565000 14.265000  5.845000 14.545000 ;
      RECT  5.565000 14.665000  5.845000 14.945000 ;
      RECT  5.565000 15.065000  5.845000 15.345000 ;
      RECT  5.565000 15.465000  5.845000 15.745000 ;
      RECT  5.565000 15.865000  5.845000 16.145000 ;
      RECT  5.565000 16.265000  5.845000 16.545000 ;
      RECT  5.565000 16.665000  5.845000 16.945000 ;
      RECT  5.565000 17.065000  5.845000 17.345000 ;
      RECT  5.565000 17.465000  5.845000 17.745000 ;
      RECT  5.565000 17.865000  5.845000 18.145000 ;
      RECT  5.565000 18.265000  5.845000 18.545000 ;
      RECT  5.565000 18.665000  5.845000 18.945000 ;
      RECT  5.565000 19.065000  5.845000 19.345000 ;
      RECT  5.565000 19.465000  5.845000 19.745000 ;
      RECT  5.565000 19.865000  5.845000 20.145000 ;
      RECT  5.565000 20.265000  5.845000 20.545000 ;
      RECT  5.565000 20.665000  5.845000 20.945000 ;
      RECT  5.565000 21.065000  5.845000 21.345000 ;
      RECT  5.565000 21.465000  5.845000 21.745000 ;
      RECT  5.565000 21.865000  5.845000 22.145000 ;
      RECT  5.965000  5.705000  6.245000  5.985000 ;
      RECT  5.965000 17.065000  6.245000 17.345000 ;
      RECT  6.025000  0.025000  6.305000  0.305000 ;
      RECT  6.025000 11.385000  6.305000 11.665000 ;
      RECT  6.025000 22.745000  6.305000 23.025000 ;
      RECT  6.365000  5.705000  6.645000  5.985000 ;
      RECT  6.365000 17.065000  6.645000 17.345000 ;
      RECT  6.425000  0.025000  6.705000  0.305000 ;
      RECT  6.425000 11.385000  6.705000 11.665000 ;
      RECT  6.425000 22.745000  6.705000 23.025000 ;
      RECT  6.765000  5.705000  7.045000  5.985000 ;
      RECT  6.765000 17.065000  7.045000 17.345000 ;
      RECT  6.825000  0.025000  7.105000  0.305000 ;
      RECT  6.825000 11.385000  7.105000 11.665000 ;
      RECT  6.825000 22.745000  7.105000 23.025000 ;
      RECT  7.165000  5.705000  7.445000  5.985000 ;
      RECT  7.165000 17.065000  7.445000 17.345000 ;
      RECT  7.225000  0.025000  7.505000  0.305000 ;
      RECT  7.225000 11.385000  7.505000 11.665000 ;
      RECT  7.225000 22.745000  7.505000 23.025000 ;
      RECT  7.565000  5.705000  7.845000  5.985000 ;
      RECT  7.565000 17.065000  7.845000 17.345000 ;
      RECT  7.625000  0.025000  7.905000  0.305000 ;
      RECT  7.625000 11.385000  7.905000 11.665000 ;
      RECT  7.625000 22.745000  7.905000 23.025000 ;
      RECT  7.965000  5.705000  8.245000  5.985000 ;
      RECT  7.965000 17.065000  8.245000 17.345000 ;
      RECT  8.025000  0.025000  8.305000  0.305000 ;
      RECT  8.025000 11.385000  8.305000 11.665000 ;
      RECT  8.025000 22.745000  8.305000 23.025000 ;
      RECT  8.365000  5.705000  8.645000  5.985000 ;
      RECT  8.365000 17.065000  8.645000 17.345000 ;
      RECT  8.425000  0.025000  8.705000  0.305000 ;
      RECT  8.425000 11.385000  8.705000 11.665000 ;
      RECT  8.425000 22.745000  8.705000 23.025000 ;
      RECT  8.765000  5.705000  9.045000  5.985000 ;
      RECT  8.765000 17.065000  9.045000 17.345000 ;
      RECT  8.825000  0.025000  9.105000  0.305000 ;
      RECT  8.825000 11.385000  9.105000 11.665000 ;
      RECT  8.825000 22.745000  9.105000 23.025000 ;
      RECT  9.165000  5.705000  9.445000  5.985000 ;
      RECT  9.165000 17.065000  9.445000 17.345000 ;
      RECT  9.225000  0.025000  9.505000  0.305000 ;
      RECT  9.225000 11.385000  9.505000 11.665000 ;
      RECT  9.225000 22.745000  9.505000 23.025000 ;
      RECT  9.565000  5.705000  9.845000  5.985000 ;
      RECT  9.565000 17.065000  9.845000 17.345000 ;
      RECT  9.625000  0.025000  9.905000  0.305000 ;
      RECT  9.625000 11.385000  9.905000 11.665000 ;
      RECT  9.625000 22.745000  9.905000 23.025000 ;
      RECT  9.965000  5.705000 10.245000  5.985000 ;
      RECT  9.965000 17.065000 10.245000 17.345000 ;
      RECT 10.025000  0.025000 10.305000  0.305000 ;
      RECT 10.025000 11.385000 10.305000 11.665000 ;
      RECT 10.025000 22.745000 10.305000 23.025000 ;
      RECT 10.365000  5.705000 10.645000  5.985000 ;
      RECT 10.365000 17.065000 10.645000 17.345000 ;
      RECT 10.425000  0.025000 10.705000  0.305000 ;
      RECT 10.425000 11.385000 10.705000 11.665000 ;
      RECT 10.425000 22.745000 10.705000 23.025000 ;
      RECT 10.825000  0.025000 11.105000  0.305000 ;
      RECT 10.825000 11.385000 11.105000 11.665000 ;
      RECT 10.825000 22.745000 11.105000 23.025000 ;
      RECT 11.105000  0.445000 11.385000  0.725000 ;
      RECT 11.105000  0.845000 11.385000  1.125000 ;
      RECT 11.105000  1.245000 11.385000  1.525000 ;
      RECT 11.105000  1.645000 11.385000  1.925000 ;
      RECT 11.105000  2.045000 11.385000  2.325000 ;
      RECT 11.105000  2.445000 11.385000  2.725000 ;
      RECT 11.105000  2.845000 11.385000  3.125000 ;
      RECT 11.105000  3.245000 11.385000  3.525000 ;
      RECT 11.105000  3.645000 11.385000  3.925000 ;
      RECT 11.105000  4.045000 11.385000  4.325000 ;
      RECT 11.105000  4.445000 11.385000  4.725000 ;
      RECT 11.105000  4.845000 11.385000  5.125000 ;
      RECT 11.105000  5.245000 11.385000  5.525000 ;
      RECT 11.105000  6.165000 11.385000  6.445000 ;
      RECT 11.105000  6.565000 11.385000  6.845000 ;
      RECT 11.105000  6.965000 11.385000  7.245000 ;
      RECT 11.105000  7.365000 11.385000  7.645000 ;
      RECT 11.105000  7.765000 11.385000  8.045000 ;
      RECT 11.105000  8.165000 11.385000  8.445000 ;
      RECT 11.105000  8.565000 11.385000  8.845000 ;
      RECT 11.105000  8.965000 11.385000  9.245000 ;
      RECT 11.105000  9.365000 11.385000  9.645000 ;
      RECT 11.105000  9.765000 11.385000 10.045000 ;
      RECT 11.105000 10.165000 11.385000 10.445000 ;
      RECT 11.105000 10.565000 11.385000 10.845000 ;
      RECT 11.105000 10.965000 11.385000 11.245000 ;
      RECT 11.105000 11.805000 11.385000 12.085000 ;
      RECT 11.105000 12.205000 11.385000 12.485000 ;
      RECT 11.105000 12.605000 11.385000 12.885000 ;
      RECT 11.105000 13.005000 11.385000 13.285000 ;
      RECT 11.105000 13.405000 11.385000 13.685000 ;
      RECT 11.105000 13.805000 11.385000 14.085000 ;
      RECT 11.105000 14.205000 11.385000 14.485000 ;
      RECT 11.105000 14.605000 11.385000 14.885000 ;
      RECT 11.105000 15.005000 11.385000 15.285000 ;
      RECT 11.105000 15.405000 11.385000 15.685000 ;
      RECT 11.105000 15.805000 11.385000 16.085000 ;
      RECT 11.105000 16.205000 11.385000 16.485000 ;
      RECT 11.105000 16.605000 11.385000 16.885000 ;
      RECT 11.105000 17.525000 11.385000 17.805000 ;
      RECT 11.105000 17.925000 11.385000 18.205000 ;
      RECT 11.105000 18.325000 11.385000 18.605000 ;
      RECT 11.105000 18.725000 11.385000 19.005000 ;
      RECT 11.105000 19.125000 11.385000 19.405000 ;
      RECT 11.105000 19.525000 11.385000 19.805000 ;
      RECT 11.105000 19.925000 11.385000 20.205000 ;
      RECT 11.105000 20.325000 11.385000 20.605000 ;
      RECT 11.105000 20.725000 11.385000 21.005000 ;
      RECT 11.105000 21.125000 11.385000 21.405000 ;
      RECT 11.105000 21.525000 11.385000 21.805000 ;
      RECT 11.105000 21.925000 11.385000 22.205000 ;
      RECT 11.105000 22.325000 11.385000 22.605000 ;
      RECT 11.385000  0.025000 11.665000  0.305000 ;
      RECT 11.385000 11.385000 11.665000 11.665000 ;
      RECT 11.385000 22.745000 11.665000 23.025000 ;
      RECT 11.785000  0.025000 12.065000  0.305000 ;
      RECT 11.785000 11.385000 12.065000 11.665000 ;
      RECT 11.785000 22.745000 12.065000 23.025000 ;
      RECT 11.845000  5.705000 12.125000  5.985000 ;
      RECT 11.845000 17.065000 12.125000 17.345000 ;
      RECT 12.185000  0.025000 12.465000  0.305000 ;
      RECT 12.185000 11.385000 12.465000 11.665000 ;
      RECT 12.185000 22.745000 12.465000 23.025000 ;
      RECT 12.245000  5.705000 12.525000  5.985000 ;
      RECT 12.245000 17.065000 12.525000 17.345000 ;
      RECT 12.585000  0.025000 12.865000  0.305000 ;
      RECT 12.585000 11.385000 12.865000 11.665000 ;
      RECT 12.585000 22.745000 12.865000 23.025000 ;
      RECT 12.645000  5.705000 12.925000  5.985000 ;
      RECT 12.645000 17.065000 12.925000 17.345000 ;
      RECT 12.985000  0.025000 13.265000  0.305000 ;
      RECT 12.985000 11.385000 13.265000 11.665000 ;
      RECT 12.985000 22.745000 13.265000 23.025000 ;
      RECT 13.045000  5.705000 13.325000  5.985000 ;
      RECT 13.045000 17.065000 13.325000 17.345000 ;
      RECT 13.385000  0.025000 13.665000  0.305000 ;
      RECT 13.385000 11.385000 13.665000 11.665000 ;
      RECT 13.385000 22.745000 13.665000 23.025000 ;
      RECT 13.445000  5.705000 13.725000  5.985000 ;
      RECT 13.445000 17.065000 13.725000 17.345000 ;
      RECT 13.785000  0.025000 14.065000  0.305000 ;
      RECT 13.785000 11.385000 14.065000 11.665000 ;
      RECT 13.785000 22.745000 14.065000 23.025000 ;
      RECT 13.845000  5.705000 14.125000  5.985000 ;
      RECT 13.845000 17.065000 14.125000 17.345000 ;
      RECT 14.185000  0.025000 14.465000  0.305000 ;
      RECT 14.185000 11.385000 14.465000 11.665000 ;
      RECT 14.185000 22.745000 14.465000 23.025000 ;
      RECT 14.245000  5.705000 14.525000  5.985000 ;
      RECT 14.245000 17.065000 14.525000 17.345000 ;
      RECT 14.585000  0.025000 14.865000  0.305000 ;
      RECT 14.585000 11.385000 14.865000 11.665000 ;
      RECT 14.585000 22.745000 14.865000 23.025000 ;
      RECT 14.645000  5.705000 14.925000  5.985000 ;
      RECT 14.645000 17.065000 14.925000 17.345000 ;
      RECT 14.985000  0.025000 15.265000  0.305000 ;
      RECT 14.985000 11.385000 15.265000 11.665000 ;
      RECT 14.985000 22.745000 15.265000 23.025000 ;
      RECT 15.045000  5.705000 15.325000  5.985000 ;
      RECT 15.045000 17.065000 15.325000 17.345000 ;
      RECT 15.385000  0.025000 15.665000  0.305000 ;
      RECT 15.385000 11.385000 15.665000 11.665000 ;
      RECT 15.385000 22.745000 15.665000 23.025000 ;
      RECT 15.445000  5.705000 15.725000  5.985000 ;
      RECT 15.445000 17.065000 15.725000 17.345000 ;
      RECT 15.785000  0.025000 16.065000  0.305000 ;
      RECT 15.785000 11.385000 16.065000 11.665000 ;
      RECT 15.785000 22.745000 16.065000 23.025000 ;
      RECT 15.845000  5.705000 16.125000  5.985000 ;
      RECT 15.845000 17.065000 16.125000 17.345000 ;
      RECT 16.185000  0.025000 16.465000  0.305000 ;
      RECT 16.185000 11.385000 16.465000 11.665000 ;
      RECT 16.185000 22.745000 16.465000 23.025000 ;
      RECT 16.245000  5.705000 16.525000  5.985000 ;
      RECT 16.245000 17.065000 16.525000 17.345000 ;
      RECT 16.645000  0.905000 16.925000  1.185000 ;
      RECT 16.645000  1.305000 16.925000  1.585000 ;
      RECT 16.645000  1.705000 16.925000  1.985000 ;
      RECT 16.645000  2.105000 16.925000  2.385000 ;
      RECT 16.645000  2.505000 16.925000  2.785000 ;
      RECT 16.645000  2.905000 16.925000  3.185000 ;
      RECT 16.645000  3.305000 16.925000  3.585000 ;
      RECT 16.645000  3.705000 16.925000  3.985000 ;
      RECT 16.645000  4.105000 16.925000  4.385000 ;
      RECT 16.645000  4.505000 16.925000  4.785000 ;
      RECT 16.645000  4.905000 16.925000  5.185000 ;
      RECT 16.645000  5.305000 16.925000  5.585000 ;
      RECT 16.645000  5.705000 16.925000  5.985000 ;
      RECT 16.645000  6.105000 16.925000  6.385000 ;
      RECT 16.645000  6.505000 16.925000  6.785000 ;
      RECT 16.645000  6.905000 16.925000  7.185000 ;
      RECT 16.645000  7.305000 16.925000  7.585000 ;
      RECT 16.645000  7.705000 16.925000  7.985000 ;
      RECT 16.645000  8.105000 16.925000  8.385000 ;
      RECT 16.645000  8.505000 16.925000  8.785000 ;
      RECT 16.645000  8.905000 16.925000  9.185000 ;
      RECT 16.645000  9.305000 16.925000  9.585000 ;
      RECT 16.645000  9.705000 16.925000  9.985000 ;
      RECT 16.645000 10.105000 16.925000 10.385000 ;
      RECT 16.645000 10.505000 16.925000 10.785000 ;
      RECT 16.645000 12.265000 16.925000 12.545000 ;
      RECT 16.645000 12.665000 16.925000 12.945000 ;
      RECT 16.645000 13.065000 16.925000 13.345000 ;
      RECT 16.645000 13.465000 16.925000 13.745000 ;
      RECT 16.645000 13.865000 16.925000 14.145000 ;
      RECT 16.645000 14.265000 16.925000 14.545000 ;
      RECT 16.645000 14.665000 16.925000 14.945000 ;
      RECT 16.645000 15.065000 16.925000 15.345000 ;
      RECT 16.645000 15.465000 16.925000 15.745000 ;
      RECT 16.645000 15.865000 16.925000 16.145000 ;
      RECT 16.645000 16.265000 16.925000 16.545000 ;
      RECT 16.645000 16.665000 16.925000 16.945000 ;
      RECT 16.645000 17.065000 16.925000 17.345000 ;
      RECT 16.645000 17.465000 16.925000 17.745000 ;
      RECT 16.645000 17.865000 16.925000 18.145000 ;
      RECT 16.645000 18.265000 16.925000 18.545000 ;
      RECT 16.645000 18.665000 16.925000 18.945000 ;
      RECT 16.645000 19.065000 16.925000 19.345000 ;
      RECT 16.645000 19.465000 16.925000 19.745000 ;
      RECT 16.645000 19.865000 16.925000 20.145000 ;
      RECT 16.645000 20.265000 16.925000 20.545000 ;
      RECT 16.645000 20.665000 16.925000 20.945000 ;
      RECT 16.645000 21.065000 16.925000 21.345000 ;
      RECT 16.645000 21.465000 16.925000 21.745000 ;
      RECT 16.645000 21.865000 16.925000 22.145000 ;
      RECT 17.045000  5.705000 17.325000  5.985000 ;
      RECT 17.045000 17.065000 17.325000 17.345000 ;
      RECT 17.105000  0.025000 17.385000  0.305000 ;
      RECT 17.105000 11.385000 17.385000 11.665000 ;
      RECT 17.105000 22.745000 17.385000 23.025000 ;
      RECT 17.445000  5.705000 17.725000  5.985000 ;
      RECT 17.445000 17.065000 17.725000 17.345000 ;
      RECT 17.505000  0.025000 17.785000  0.305000 ;
      RECT 17.505000 11.385000 17.785000 11.665000 ;
      RECT 17.505000 22.745000 17.785000 23.025000 ;
      RECT 17.845000  5.705000 18.125000  5.985000 ;
      RECT 17.845000 17.065000 18.125000 17.345000 ;
      RECT 17.905000  0.025000 18.185000  0.305000 ;
      RECT 17.905000 11.385000 18.185000 11.665000 ;
      RECT 17.905000 22.745000 18.185000 23.025000 ;
      RECT 18.245000  5.705000 18.525000  5.985000 ;
      RECT 18.245000 17.065000 18.525000 17.345000 ;
      RECT 18.305000  0.025000 18.585000  0.305000 ;
      RECT 18.305000 11.385000 18.585000 11.665000 ;
      RECT 18.305000 22.745000 18.585000 23.025000 ;
      RECT 18.645000  5.705000 18.925000  5.985000 ;
      RECT 18.645000 17.065000 18.925000 17.345000 ;
      RECT 18.705000  0.025000 18.985000  0.305000 ;
      RECT 18.705000 11.385000 18.985000 11.665000 ;
      RECT 18.705000 22.745000 18.985000 23.025000 ;
      RECT 19.045000  5.705000 19.325000  5.985000 ;
      RECT 19.045000 17.065000 19.325000 17.345000 ;
      RECT 19.105000  0.025000 19.385000  0.305000 ;
      RECT 19.105000 11.385000 19.385000 11.665000 ;
      RECT 19.105000 22.745000 19.385000 23.025000 ;
      RECT 19.445000  5.705000 19.725000  5.985000 ;
      RECT 19.445000 17.065000 19.725000 17.345000 ;
      RECT 19.505000  0.025000 19.785000  0.305000 ;
      RECT 19.505000 11.385000 19.785000 11.665000 ;
      RECT 19.505000 22.745000 19.785000 23.025000 ;
      RECT 19.845000  5.705000 20.125000  5.985000 ;
      RECT 19.845000 17.065000 20.125000 17.345000 ;
      RECT 19.905000  0.025000 20.185000  0.305000 ;
      RECT 19.905000 11.385000 20.185000 11.665000 ;
      RECT 19.905000 22.745000 20.185000 23.025000 ;
      RECT 20.245000  5.705000 20.525000  5.985000 ;
      RECT 20.245000 17.065000 20.525000 17.345000 ;
      RECT 20.305000  0.025000 20.585000  0.305000 ;
      RECT 20.305000 11.385000 20.585000 11.665000 ;
      RECT 20.305000 22.745000 20.585000 23.025000 ;
      RECT 20.645000  5.705000 20.925000  5.985000 ;
      RECT 20.645000 17.065000 20.925000 17.345000 ;
      RECT 20.705000  0.025000 20.985000  0.305000 ;
      RECT 20.705000 11.385000 20.985000 11.665000 ;
      RECT 20.705000 22.745000 20.985000 23.025000 ;
      RECT 21.045000  5.705000 21.325000  5.985000 ;
      RECT 21.045000 17.065000 21.325000 17.345000 ;
      RECT 21.105000  0.025000 21.385000  0.305000 ;
      RECT 21.105000 11.385000 21.385000 11.665000 ;
      RECT 21.105000 22.745000 21.385000 23.025000 ;
      RECT 21.445000  5.705000 21.725000  5.985000 ;
      RECT 21.445000 17.065000 21.725000 17.345000 ;
      RECT 21.505000  0.025000 21.785000  0.305000 ;
      RECT 21.505000 11.385000 21.785000 11.665000 ;
      RECT 21.505000 22.745000 21.785000 23.025000 ;
      RECT 21.905000  0.025000 22.185000  0.305000 ;
      RECT 21.905000 11.385000 22.185000 11.665000 ;
      RECT 21.905000 22.745000 22.185000 23.025000 ;
      RECT 22.185000  0.445000 22.465000  0.725000 ;
      RECT 22.185000  0.845000 22.465000  1.125000 ;
      RECT 22.185000  1.245000 22.465000  1.525000 ;
      RECT 22.185000  1.645000 22.465000  1.925000 ;
      RECT 22.185000  2.045000 22.465000  2.325000 ;
      RECT 22.185000  2.445000 22.465000  2.725000 ;
      RECT 22.185000  2.845000 22.465000  3.125000 ;
      RECT 22.185000  3.245000 22.465000  3.525000 ;
      RECT 22.185000  3.645000 22.465000  3.925000 ;
      RECT 22.185000  4.045000 22.465000  4.325000 ;
      RECT 22.185000  4.445000 22.465000  4.725000 ;
      RECT 22.185000  4.845000 22.465000  5.125000 ;
      RECT 22.185000  5.245000 22.465000  5.525000 ;
      RECT 22.185000  6.165000 22.465000  6.445000 ;
      RECT 22.185000  6.565000 22.465000  6.845000 ;
      RECT 22.185000  6.965000 22.465000  7.245000 ;
      RECT 22.185000  7.365000 22.465000  7.645000 ;
      RECT 22.185000  7.765000 22.465000  8.045000 ;
      RECT 22.185000  8.165000 22.465000  8.445000 ;
      RECT 22.185000  8.565000 22.465000  8.845000 ;
      RECT 22.185000  8.965000 22.465000  9.245000 ;
      RECT 22.185000  9.365000 22.465000  9.645000 ;
      RECT 22.185000  9.765000 22.465000 10.045000 ;
      RECT 22.185000 10.165000 22.465000 10.445000 ;
      RECT 22.185000 10.565000 22.465000 10.845000 ;
      RECT 22.185000 10.965000 22.465000 11.245000 ;
      RECT 22.185000 11.805000 22.465000 12.085000 ;
      RECT 22.185000 12.205000 22.465000 12.485000 ;
      RECT 22.185000 12.605000 22.465000 12.885000 ;
      RECT 22.185000 13.005000 22.465000 13.285000 ;
      RECT 22.185000 13.405000 22.465000 13.685000 ;
      RECT 22.185000 13.805000 22.465000 14.085000 ;
      RECT 22.185000 14.205000 22.465000 14.485000 ;
      RECT 22.185000 14.605000 22.465000 14.885000 ;
      RECT 22.185000 15.005000 22.465000 15.285000 ;
      RECT 22.185000 15.405000 22.465000 15.685000 ;
      RECT 22.185000 15.805000 22.465000 16.085000 ;
      RECT 22.185000 16.205000 22.465000 16.485000 ;
      RECT 22.185000 16.605000 22.465000 16.885000 ;
      RECT 22.185000 17.525000 22.465000 17.805000 ;
      RECT 22.185000 17.925000 22.465000 18.205000 ;
      RECT 22.185000 18.325000 22.465000 18.605000 ;
      RECT 22.185000 18.725000 22.465000 19.005000 ;
      RECT 22.185000 19.125000 22.465000 19.405000 ;
      RECT 22.185000 19.525000 22.465000 19.805000 ;
      RECT 22.185000 19.925000 22.465000 20.205000 ;
      RECT 22.185000 20.325000 22.465000 20.605000 ;
      RECT 22.185000 20.725000 22.465000 21.005000 ;
      RECT 22.185000 21.125000 22.465000 21.405000 ;
      RECT 22.185000 21.525000 22.465000 21.805000 ;
      RECT 22.185000 21.925000 22.465000 22.205000 ;
      RECT 22.185000 22.325000 22.465000 22.605000 ;
  END
END sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top
END LIBRARY
