* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox_slope=0.80e-2
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox2_slope=0.86e-2  $ for L>=4 and W<=0.75
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox3_slope=0.55e-2  $ for L>=4 and W>=3.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox4_slope=2.55e-2  $ for L<=0.6 and W<=3.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox_offset=0.000
.param sky130_fd_pr__rf_nfet_g5v0d10v5__nfactor_slope=0.000
.param sky130_fd_pr__rf_nfet_g5v0d10v5__voff_slope=0.00375
.param sky130_fd_pr__rf_nfet_g5v0d10v5__voff2_slope=0.00850 $ for L>=4 and W=0.42
.param sky130_fd_pr__rf_nfet_g5v0d10v5__lint_slope=3.0e-09
.param sky130_fd_pr__rf_nfet_g5v0d10v5__lint1_slope=0.0e-09
.param sky130_fd_pr__rf_nfet_g5v0d10v5__wint_slope=0.0e-11  $ Not used
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope= .80e-2
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1= 2.05e-2 $ All W with L=0.5um
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope2= 1.00e-2 $ W=3 L=1 um All W with L=0.8um & L=0.6um
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope3= 0.67e-2 $ All W with L=4.0um
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_vth0_slope=0.000  $ All devices
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope=0.13  $ All devices
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope=0.12  $ All devices
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_lint_slope=0.0  $ All devices
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_wint_slope=0.0  $ All devices
