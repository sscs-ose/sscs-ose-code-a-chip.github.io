MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 49.15 BY 27.64 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 9.75 2.78 10.03 7.3 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.98 8.26 19.52 8.54 ;
      LAYER M3 ;
        RECT 27.38 8.24 27.66 20.32 ;
      LAYER M2 ;
        RECT 19.35 8.26 21.07 8.54 ;
      LAYER M3 ;
        RECT 20.93 8.4 21.21 8.82 ;
      LAYER M4 ;
        RECT 21.07 8.42 27.52 9.22 ;
      LAYER M3 ;
        RECT 27.38 8.635 27.66 9.005 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 28.64 2.8 39.3 3.08 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 29.5 2.38 40.16 2.66 ;
    END
  END VINP
  OBS 
  LAYER M2 ;
        RECT 5.42 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 0.69 8.68 19.95 8.96 ;
  LAYER M2 ;
        RECT 28.21 6.16 40.59 6.44 ;
  LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
  LAYER M3 ;
        RECT 15.77 6.72 16.05 8.82 ;
  LAYER M2 ;
        RECT 15.75 8.68 16.07 8.96 ;
  LAYER M2 ;
        RECT 19.62 8.68 19.94 8.96 ;
  LAYER M3 ;
        RECT 19.64 6.3 19.92 8.82 ;
  LAYER M2 ;
        RECT 19.78 6.16 28.38 6.44 ;
  LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
  LAYER M3 ;
        RECT 15.77 6.56 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.75 8.68 16.07 8.96 ;
  LAYER M3 ;
        RECT 15.77 8.66 16.05 8.98 ;
  LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
  LAYER M3 ;
        RECT 15.77 6.56 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.75 8.68 16.07 8.96 ;
  LAYER M3 ;
        RECT 15.77 8.66 16.05 8.98 ;
  LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
  LAYER M3 ;
        RECT 15.77 6.56 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.75 8.68 16.07 8.96 ;
  LAYER M3 ;
        RECT 15.77 8.66 16.05 8.98 ;
  LAYER M2 ;
        RECT 19.62 6.16 19.94 6.44 ;
  LAYER M3 ;
        RECT 19.64 6.14 19.92 6.46 ;
  LAYER M2 ;
        RECT 19.62 8.68 19.94 8.96 ;
  LAYER M3 ;
        RECT 19.64 8.66 19.92 8.98 ;
  LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
  LAYER M3 ;
        RECT 15.77 6.56 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.75 8.68 16.07 8.96 ;
  LAYER M3 ;
        RECT 15.77 8.66 16.05 8.98 ;
  LAYER M2 ;
        RECT 19.62 6.16 19.94 6.44 ;
  LAYER M3 ;
        RECT 19.64 6.14 19.92 6.46 ;
  LAYER M2 ;
        RECT 19.62 8.68 19.94 8.96 ;
  LAYER M3 ;
        RECT 19.64 8.66 19.92 8.98 ;
  LAYER M2 ;
        RECT 28.64 7 39.3 7.28 ;
  LAYER M3 ;
        RECT 27.81 7.82 28.09 24.1 ;
  LAYER M2 ;
        RECT 27.95 7 28.81 7.28 ;
  LAYER M3 ;
        RECT 27.81 7.14 28.09 7.98 ;
  LAYER M2 ;
        RECT 27.79 7 28.11 7.28 ;
  LAYER M3 ;
        RECT 27.81 6.98 28.09 7.3 ;
  LAYER M2 ;
        RECT 27.79 7 28.11 7.28 ;
  LAYER M3 ;
        RECT 27.81 6.98 28.09 7.3 ;
  LAYER M2 ;
        RECT 29.5 6.58 40.16 6.86 ;
  LAYER M3 ;
        RECT 40.71 7.82 40.99 24.1 ;
  LAYER M2 ;
        RECT 39.83 6.58 40.15 6.86 ;
  LAYER M3 ;
        RECT 39.85 6.72 40.13 7.14 ;
  LAYER M2 ;
        RECT 39.99 7 40.85 7.28 ;
  LAYER M3 ;
        RECT 40.71 7.14 40.99 7.98 ;
  LAYER M2 ;
        RECT 39.83 6.58 40.15 6.86 ;
  LAYER M3 ;
        RECT 39.85 6.56 40.13 6.88 ;
  LAYER M2 ;
        RECT 39.83 7 40.15 7.28 ;
  LAYER M3 ;
        RECT 39.85 6.98 40.13 7.3 ;
  LAYER M2 ;
        RECT 40.69 7 41.01 7.28 ;
  LAYER M3 ;
        RECT 40.71 6.98 40.99 7.3 ;
  LAYER M2 ;
        RECT 39.83 6.58 40.15 6.86 ;
  LAYER M3 ;
        RECT 39.85 6.56 40.13 6.88 ;
  LAYER M2 ;
        RECT 39.83 7 40.15 7.28 ;
  LAYER M3 ;
        RECT 39.85 6.98 40.13 7.3 ;
  LAYER M2 ;
        RECT 40.69 7 41.01 7.28 ;
  LAYER M3 ;
        RECT 40.71 6.98 40.99 7.3 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 12.34 ;
  LAYER M3 ;
        RECT 41.14 8.24 41.42 20.32 ;
  LAYER M3 ;
        RECT 9.75 11.575 10.03 11.945 ;
  LAYER M2 ;
        RECT 9.89 11.62 41.28 11.9 ;
  LAYER M3 ;
        RECT 41.14 11.575 41.42 11.945 ;
  LAYER M2 ;
        RECT 9.73 11.62 10.05 11.9 ;
  LAYER M3 ;
        RECT 9.75 11.6 10.03 11.92 ;
  LAYER M2 ;
        RECT 41.12 11.62 41.44 11.9 ;
  LAYER M3 ;
        RECT 41.14 11.6 41.42 11.92 ;
  LAYER M2 ;
        RECT 9.73 11.62 10.05 11.9 ;
  LAYER M3 ;
        RECT 9.75 11.6 10.03 11.92 ;
  LAYER M2 ;
        RECT 41.12 11.62 41.44 11.9 ;
  LAYER M3 ;
        RECT 41.14 11.6 41.42 11.92 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 16.08 3.08 ;
  LAYER M2 ;
        RECT 4.56 0.7 16.08 0.98 ;
  LAYER M2 ;
        RECT 4.13 6.16 16.51 6.44 ;
  LAYER M3 ;
        RECT 9.75 2.78 10.03 7.3 ;
  LAYER M2 ;
        RECT 5.42 6.58 16.08 6.86 ;
  LAYER M3 ;
        RECT 10.61 0.68 10.89 6.46 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 11.425 ;
  LAYER M1 ;
        RECT 32.985 11.675 33.235 12.685 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 17.305 ;
  LAYER M1 ;
        RECT 32.985 17.555 33.235 18.565 ;
  LAYER M1 ;
        RECT 32.985 19.655 33.235 23.185 ;
  LAYER M1 ;
        RECT 32.985 23.435 33.235 24.445 ;
  LAYER M1 ;
        RECT 32.985 25.535 33.235 26.545 ;
  LAYER M1 ;
        RECT 33.415 7.895 33.665 11.425 ;
  LAYER M1 ;
        RECT 33.415 13.775 33.665 17.305 ;
  LAYER M1 ;
        RECT 33.415 19.655 33.665 23.185 ;
  LAYER M1 ;
        RECT 32.555 7.895 32.805 11.425 ;
  LAYER M1 ;
        RECT 32.555 13.775 32.805 17.305 ;
  LAYER M1 ;
        RECT 32.555 19.655 32.805 23.185 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 11.425 ;
  LAYER M1 ;
        RECT 32.125 11.675 32.375 12.685 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 17.305 ;
  LAYER M1 ;
        RECT 32.125 17.555 32.375 18.565 ;
  LAYER M1 ;
        RECT 32.125 19.655 32.375 23.185 ;
  LAYER M1 ;
        RECT 32.125 23.435 32.375 24.445 ;
  LAYER M1 ;
        RECT 32.125 25.535 32.375 26.545 ;
  LAYER M1 ;
        RECT 31.695 7.895 31.945 11.425 ;
  LAYER M1 ;
        RECT 31.695 13.775 31.945 17.305 ;
  LAYER M1 ;
        RECT 31.695 19.655 31.945 23.185 ;
  LAYER M1 ;
        RECT 31.265 7.895 31.515 11.425 ;
  LAYER M1 ;
        RECT 31.265 11.675 31.515 12.685 ;
  LAYER M1 ;
        RECT 31.265 13.775 31.515 17.305 ;
  LAYER M1 ;
        RECT 31.265 17.555 31.515 18.565 ;
  LAYER M1 ;
        RECT 31.265 19.655 31.515 23.185 ;
  LAYER M1 ;
        RECT 31.265 23.435 31.515 24.445 ;
  LAYER M1 ;
        RECT 31.265 25.535 31.515 26.545 ;
  LAYER M1 ;
        RECT 30.835 7.895 31.085 11.425 ;
  LAYER M1 ;
        RECT 30.835 13.775 31.085 17.305 ;
  LAYER M1 ;
        RECT 30.835 19.655 31.085 23.185 ;
  LAYER M1 ;
        RECT 30.405 7.895 30.655 11.425 ;
  LAYER M1 ;
        RECT 30.405 11.675 30.655 12.685 ;
  LAYER M1 ;
        RECT 30.405 13.775 30.655 17.305 ;
  LAYER M1 ;
        RECT 30.405 17.555 30.655 18.565 ;
  LAYER M1 ;
        RECT 30.405 19.655 30.655 23.185 ;
  LAYER M1 ;
        RECT 30.405 23.435 30.655 24.445 ;
  LAYER M1 ;
        RECT 30.405 25.535 30.655 26.545 ;
  LAYER M1 ;
        RECT 29.975 7.895 30.225 11.425 ;
  LAYER M1 ;
        RECT 29.975 13.775 30.225 17.305 ;
  LAYER M1 ;
        RECT 29.975 19.655 30.225 23.185 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 11.425 ;
  LAYER M1 ;
        RECT 29.545 11.675 29.795 12.685 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 17.305 ;
  LAYER M1 ;
        RECT 29.545 17.555 29.795 18.565 ;
  LAYER M1 ;
        RECT 29.545 19.655 29.795 23.185 ;
  LAYER M1 ;
        RECT 29.545 23.435 29.795 24.445 ;
  LAYER M1 ;
        RECT 29.545 25.535 29.795 26.545 ;
  LAYER M1 ;
        RECT 29.115 7.895 29.365 11.425 ;
  LAYER M1 ;
        RECT 29.115 13.775 29.365 17.305 ;
  LAYER M1 ;
        RECT 29.115 19.655 29.365 23.185 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 11.425 ;
  LAYER M1 ;
        RECT 28.685 11.675 28.935 12.685 ;
  LAYER M1 ;
        RECT 28.685 13.775 28.935 17.305 ;
  LAYER M1 ;
        RECT 28.685 17.555 28.935 18.565 ;
  LAYER M1 ;
        RECT 28.685 19.655 28.935 23.185 ;
  LAYER M1 ;
        RECT 28.685 23.435 28.935 24.445 ;
  LAYER M1 ;
        RECT 28.685 25.535 28.935 26.545 ;
  LAYER M1 ;
        RECT 28.255 7.895 28.505 11.425 ;
  LAYER M1 ;
        RECT 28.255 13.775 28.505 17.305 ;
  LAYER M1 ;
        RECT 28.255 19.655 28.505 23.185 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 11.425 ;
  LAYER M1 ;
        RECT 27.825 11.675 28.075 12.685 ;
  LAYER M1 ;
        RECT 27.825 13.775 28.075 17.305 ;
  LAYER M1 ;
        RECT 27.825 17.555 28.075 18.565 ;
  LAYER M1 ;
        RECT 27.825 19.655 28.075 23.185 ;
  LAYER M1 ;
        RECT 27.825 23.435 28.075 24.445 ;
  LAYER M1 ;
        RECT 27.825 25.535 28.075 26.545 ;
  LAYER M1 ;
        RECT 27.395 7.895 27.645 11.425 ;
  LAYER M1 ;
        RECT 27.395 13.775 27.645 17.305 ;
  LAYER M1 ;
        RECT 27.395 19.655 27.645 23.185 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 11.425 ;
  LAYER M1 ;
        RECT 26.965 11.675 27.215 12.685 ;
  LAYER M1 ;
        RECT 26.965 13.775 27.215 17.305 ;
  LAYER M1 ;
        RECT 26.965 17.555 27.215 18.565 ;
  LAYER M1 ;
        RECT 26.965 19.655 27.215 23.185 ;
  LAYER M1 ;
        RECT 26.965 23.435 27.215 24.445 ;
  LAYER M1 ;
        RECT 26.965 25.535 27.215 26.545 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M1 ;
        RECT 26.535 13.775 26.785 17.305 ;
  LAYER M1 ;
        RECT 26.535 19.655 26.785 23.185 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 11.425 ;
  LAYER M1 ;
        RECT 26.105 11.675 26.355 12.685 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 17.305 ;
  LAYER M1 ;
        RECT 26.105 17.555 26.355 18.565 ;
  LAYER M1 ;
        RECT 26.105 19.655 26.355 23.185 ;
  LAYER M1 ;
        RECT 26.105 23.435 26.355 24.445 ;
  LAYER M1 ;
        RECT 26.105 25.535 26.355 26.545 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 25.675 13.775 25.925 17.305 ;
  LAYER M1 ;
        RECT 25.675 19.655 25.925 23.185 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 11.425 ;
  LAYER M1 ;
        RECT 25.245 11.675 25.495 12.685 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 17.305 ;
  LAYER M1 ;
        RECT 25.245 17.555 25.495 18.565 ;
  LAYER M1 ;
        RECT 25.245 19.655 25.495 23.185 ;
  LAYER M1 ;
        RECT 25.245 23.435 25.495 24.445 ;
  LAYER M1 ;
        RECT 25.245 25.535 25.495 26.545 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M1 ;
        RECT 24.815 13.775 25.065 17.305 ;
  LAYER M1 ;
        RECT 24.815 19.655 25.065 23.185 ;
  LAYER M1 ;
        RECT 24.385 7.895 24.635 11.425 ;
  LAYER M1 ;
        RECT 24.385 11.675 24.635 12.685 ;
  LAYER M1 ;
        RECT 24.385 13.775 24.635 17.305 ;
  LAYER M1 ;
        RECT 24.385 17.555 24.635 18.565 ;
  LAYER M1 ;
        RECT 24.385 19.655 24.635 23.185 ;
  LAYER M1 ;
        RECT 24.385 23.435 24.635 24.445 ;
  LAYER M1 ;
        RECT 24.385 25.535 24.635 26.545 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M1 ;
        RECT 23.955 13.775 24.205 17.305 ;
  LAYER M1 ;
        RECT 23.955 19.655 24.205 23.185 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 11.425 ;
  LAYER M1 ;
        RECT 23.525 11.675 23.775 12.685 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 17.305 ;
  LAYER M1 ;
        RECT 23.525 17.555 23.775 18.565 ;
  LAYER M1 ;
        RECT 23.525 19.655 23.775 23.185 ;
  LAYER M1 ;
        RECT 23.525 23.435 23.775 24.445 ;
  LAYER M1 ;
        RECT 23.525 25.535 23.775 26.545 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 23.095 13.775 23.345 17.305 ;
  LAYER M1 ;
        RECT 23.095 19.655 23.345 23.185 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 22.665 11.675 22.915 12.685 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 17.305 ;
  LAYER M1 ;
        RECT 22.665 17.555 22.915 18.565 ;
  LAYER M1 ;
        RECT 22.665 19.655 22.915 23.185 ;
  LAYER M1 ;
        RECT 22.665 23.435 22.915 24.445 ;
  LAYER M1 ;
        RECT 22.665 25.535 22.915 26.545 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 22.235 19.655 22.485 23.185 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 17.305 ;
  LAYER M1 ;
        RECT 21.805 17.555 22.055 18.565 ;
  LAYER M1 ;
        RECT 21.805 19.655 22.055 23.185 ;
  LAYER M1 ;
        RECT 21.805 23.435 22.055 24.445 ;
  LAYER M1 ;
        RECT 21.805 25.535 22.055 26.545 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M1 ;
        RECT 21.375 13.775 21.625 17.305 ;
  LAYER M1 ;
        RECT 21.375 19.655 21.625 23.185 ;
  LAYER M2 ;
        RECT 22.62 7.84 33.28 8.12 ;
  LAYER M2 ;
        RECT 21.76 12.04 33.28 12.32 ;
  LAYER M2 ;
        RECT 21.76 8.26 32.42 8.54 ;
  LAYER M2 ;
        RECT 21.33 8.68 33.71 8.96 ;
  LAYER M2 ;
        RECT 21.76 13.72 32.42 14 ;
  LAYER M2 ;
        RECT 21.76 17.92 33.28 18.2 ;
  LAYER M2 ;
        RECT 22.62 14.14 33.28 14.42 ;
  LAYER M2 ;
        RECT 21.33 14.56 33.71 14.84 ;
  LAYER M2 ;
        RECT 22.62 19.6 33.28 19.88 ;
  LAYER M2 ;
        RECT 21.76 23.8 33.28 24.08 ;
  LAYER M2 ;
        RECT 21.76 20.02 32.42 20.3 ;
  LAYER M2 ;
        RECT 21.76 25.9 33.28 26.18 ;
  LAYER M2 ;
        RECT 21.33 20.44 33.71 20.72 ;
  LAYER M3 ;
        RECT 27.81 7.82 28.09 24.1 ;
  LAYER M3 ;
        RECT 27.38 8.24 27.66 20.32 ;
  LAYER M3 ;
        RECT 26.95 8.66 27.23 26.2 ;
  LAYER M1 ;
        RECT 35.565 7.895 35.815 11.425 ;
  LAYER M1 ;
        RECT 35.565 11.675 35.815 12.685 ;
  LAYER M1 ;
        RECT 35.565 13.775 35.815 17.305 ;
  LAYER M1 ;
        RECT 35.565 17.555 35.815 18.565 ;
  LAYER M1 ;
        RECT 35.565 19.655 35.815 23.185 ;
  LAYER M1 ;
        RECT 35.565 23.435 35.815 24.445 ;
  LAYER M1 ;
        RECT 35.565 25.535 35.815 26.545 ;
  LAYER M1 ;
        RECT 35.135 7.895 35.385 11.425 ;
  LAYER M1 ;
        RECT 35.135 13.775 35.385 17.305 ;
  LAYER M1 ;
        RECT 35.135 19.655 35.385 23.185 ;
  LAYER M1 ;
        RECT 35.995 7.895 36.245 11.425 ;
  LAYER M1 ;
        RECT 35.995 13.775 36.245 17.305 ;
  LAYER M1 ;
        RECT 35.995 19.655 36.245 23.185 ;
  LAYER M1 ;
        RECT 36.425 7.895 36.675 11.425 ;
  LAYER M1 ;
        RECT 36.425 11.675 36.675 12.685 ;
  LAYER M1 ;
        RECT 36.425 13.775 36.675 17.305 ;
  LAYER M1 ;
        RECT 36.425 17.555 36.675 18.565 ;
  LAYER M1 ;
        RECT 36.425 19.655 36.675 23.185 ;
  LAYER M1 ;
        RECT 36.425 23.435 36.675 24.445 ;
  LAYER M1 ;
        RECT 36.425 25.535 36.675 26.545 ;
  LAYER M1 ;
        RECT 36.855 7.895 37.105 11.425 ;
  LAYER M1 ;
        RECT 36.855 13.775 37.105 17.305 ;
  LAYER M1 ;
        RECT 36.855 19.655 37.105 23.185 ;
  LAYER M1 ;
        RECT 37.285 7.895 37.535 11.425 ;
  LAYER M1 ;
        RECT 37.285 11.675 37.535 12.685 ;
  LAYER M1 ;
        RECT 37.285 13.775 37.535 17.305 ;
  LAYER M1 ;
        RECT 37.285 17.555 37.535 18.565 ;
  LAYER M1 ;
        RECT 37.285 19.655 37.535 23.185 ;
  LAYER M1 ;
        RECT 37.285 23.435 37.535 24.445 ;
  LAYER M1 ;
        RECT 37.285 25.535 37.535 26.545 ;
  LAYER M1 ;
        RECT 37.715 7.895 37.965 11.425 ;
  LAYER M1 ;
        RECT 37.715 13.775 37.965 17.305 ;
  LAYER M1 ;
        RECT 37.715 19.655 37.965 23.185 ;
  LAYER M1 ;
        RECT 38.145 7.895 38.395 11.425 ;
  LAYER M1 ;
        RECT 38.145 11.675 38.395 12.685 ;
  LAYER M1 ;
        RECT 38.145 13.775 38.395 17.305 ;
  LAYER M1 ;
        RECT 38.145 17.555 38.395 18.565 ;
  LAYER M1 ;
        RECT 38.145 19.655 38.395 23.185 ;
  LAYER M1 ;
        RECT 38.145 23.435 38.395 24.445 ;
  LAYER M1 ;
        RECT 38.145 25.535 38.395 26.545 ;
  LAYER M1 ;
        RECT 38.575 7.895 38.825 11.425 ;
  LAYER M1 ;
        RECT 38.575 13.775 38.825 17.305 ;
  LAYER M1 ;
        RECT 38.575 19.655 38.825 23.185 ;
  LAYER M1 ;
        RECT 39.005 7.895 39.255 11.425 ;
  LAYER M1 ;
        RECT 39.005 11.675 39.255 12.685 ;
  LAYER M1 ;
        RECT 39.005 13.775 39.255 17.305 ;
  LAYER M1 ;
        RECT 39.005 17.555 39.255 18.565 ;
  LAYER M1 ;
        RECT 39.005 19.655 39.255 23.185 ;
  LAYER M1 ;
        RECT 39.005 23.435 39.255 24.445 ;
  LAYER M1 ;
        RECT 39.005 25.535 39.255 26.545 ;
  LAYER M1 ;
        RECT 39.435 7.895 39.685 11.425 ;
  LAYER M1 ;
        RECT 39.435 13.775 39.685 17.305 ;
  LAYER M1 ;
        RECT 39.435 19.655 39.685 23.185 ;
  LAYER M1 ;
        RECT 39.865 7.895 40.115 11.425 ;
  LAYER M1 ;
        RECT 39.865 11.675 40.115 12.685 ;
  LAYER M1 ;
        RECT 39.865 13.775 40.115 17.305 ;
  LAYER M1 ;
        RECT 39.865 17.555 40.115 18.565 ;
  LAYER M1 ;
        RECT 39.865 19.655 40.115 23.185 ;
  LAYER M1 ;
        RECT 39.865 23.435 40.115 24.445 ;
  LAYER M1 ;
        RECT 39.865 25.535 40.115 26.545 ;
  LAYER M1 ;
        RECT 40.295 7.895 40.545 11.425 ;
  LAYER M1 ;
        RECT 40.295 13.775 40.545 17.305 ;
  LAYER M1 ;
        RECT 40.295 19.655 40.545 23.185 ;
  LAYER M1 ;
        RECT 40.725 7.895 40.975 11.425 ;
  LAYER M1 ;
        RECT 40.725 11.675 40.975 12.685 ;
  LAYER M1 ;
        RECT 40.725 13.775 40.975 17.305 ;
  LAYER M1 ;
        RECT 40.725 17.555 40.975 18.565 ;
  LAYER M1 ;
        RECT 40.725 19.655 40.975 23.185 ;
  LAYER M1 ;
        RECT 40.725 23.435 40.975 24.445 ;
  LAYER M1 ;
        RECT 40.725 25.535 40.975 26.545 ;
  LAYER M1 ;
        RECT 41.155 7.895 41.405 11.425 ;
  LAYER M1 ;
        RECT 41.155 13.775 41.405 17.305 ;
  LAYER M1 ;
        RECT 41.155 19.655 41.405 23.185 ;
  LAYER M1 ;
        RECT 41.585 7.895 41.835 11.425 ;
  LAYER M1 ;
        RECT 41.585 11.675 41.835 12.685 ;
  LAYER M1 ;
        RECT 41.585 13.775 41.835 17.305 ;
  LAYER M1 ;
        RECT 41.585 17.555 41.835 18.565 ;
  LAYER M1 ;
        RECT 41.585 19.655 41.835 23.185 ;
  LAYER M1 ;
        RECT 41.585 23.435 41.835 24.445 ;
  LAYER M1 ;
        RECT 41.585 25.535 41.835 26.545 ;
  LAYER M1 ;
        RECT 42.015 7.895 42.265 11.425 ;
  LAYER M1 ;
        RECT 42.015 13.775 42.265 17.305 ;
  LAYER M1 ;
        RECT 42.015 19.655 42.265 23.185 ;
  LAYER M1 ;
        RECT 42.445 7.895 42.695 11.425 ;
  LAYER M1 ;
        RECT 42.445 11.675 42.695 12.685 ;
  LAYER M1 ;
        RECT 42.445 13.775 42.695 17.305 ;
  LAYER M1 ;
        RECT 42.445 17.555 42.695 18.565 ;
  LAYER M1 ;
        RECT 42.445 19.655 42.695 23.185 ;
  LAYER M1 ;
        RECT 42.445 23.435 42.695 24.445 ;
  LAYER M1 ;
        RECT 42.445 25.535 42.695 26.545 ;
  LAYER M1 ;
        RECT 42.875 7.895 43.125 11.425 ;
  LAYER M1 ;
        RECT 42.875 13.775 43.125 17.305 ;
  LAYER M1 ;
        RECT 42.875 19.655 43.125 23.185 ;
  LAYER M1 ;
        RECT 43.305 7.895 43.555 11.425 ;
  LAYER M1 ;
        RECT 43.305 11.675 43.555 12.685 ;
  LAYER M1 ;
        RECT 43.305 13.775 43.555 17.305 ;
  LAYER M1 ;
        RECT 43.305 17.555 43.555 18.565 ;
  LAYER M1 ;
        RECT 43.305 19.655 43.555 23.185 ;
  LAYER M1 ;
        RECT 43.305 23.435 43.555 24.445 ;
  LAYER M1 ;
        RECT 43.305 25.535 43.555 26.545 ;
  LAYER M1 ;
        RECT 43.735 7.895 43.985 11.425 ;
  LAYER M1 ;
        RECT 43.735 13.775 43.985 17.305 ;
  LAYER M1 ;
        RECT 43.735 19.655 43.985 23.185 ;
  LAYER M1 ;
        RECT 44.165 7.895 44.415 11.425 ;
  LAYER M1 ;
        RECT 44.165 11.675 44.415 12.685 ;
  LAYER M1 ;
        RECT 44.165 13.775 44.415 17.305 ;
  LAYER M1 ;
        RECT 44.165 17.555 44.415 18.565 ;
  LAYER M1 ;
        RECT 44.165 19.655 44.415 23.185 ;
  LAYER M1 ;
        RECT 44.165 23.435 44.415 24.445 ;
  LAYER M1 ;
        RECT 44.165 25.535 44.415 26.545 ;
  LAYER M1 ;
        RECT 44.595 7.895 44.845 11.425 ;
  LAYER M1 ;
        RECT 44.595 13.775 44.845 17.305 ;
  LAYER M1 ;
        RECT 44.595 19.655 44.845 23.185 ;
  LAYER M1 ;
        RECT 45.025 7.895 45.275 11.425 ;
  LAYER M1 ;
        RECT 45.025 11.675 45.275 12.685 ;
  LAYER M1 ;
        RECT 45.025 13.775 45.275 17.305 ;
  LAYER M1 ;
        RECT 45.025 17.555 45.275 18.565 ;
  LAYER M1 ;
        RECT 45.025 19.655 45.275 23.185 ;
  LAYER M1 ;
        RECT 45.025 23.435 45.275 24.445 ;
  LAYER M1 ;
        RECT 45.025 25.535 45.275 26.545 ;
  LAYER M1 ;
        RECT 45.455 7.895 45.705 11.425 ;
  LAYER M1 ;
        RECT 45.455 13.775 45.705 17.305 ;
  LAYER M1 ;
        RECT 45.455 19.655 45.705 23.185 ;
  LAYER M1 ;
        RECT 45.885 7.895 46.135 11.425 ;
  LAYER M1 ;
        RECT 45.885 11.675 46.135 12.685 ;
  LAYER M1 ;
        RECT 45.885 13.775 46.135 17.305 ;
  LAYER M1 ;
        RECT 45.885 17.555 46.135 18.565 ;
  LAYER M1 ;
        RECT 45.885 19.655 46.135 23.185 ;
  LAYER M1 ;
        RECT 45.885 23.435 46.135 24.445 ;
  LAYER M1 ;
        RECT 45.885 25.535 46.135 26.545 ;
  LAYER M1 ;
        RECT 46.315 7.895 46.565 11.425 ;
  LAYER M1 ;
        RECT 46.315 13.775 46.565 17.305 ;
  LAYER M1 ;
        RECT 46.315 19.655 46.565 23.185 ;
  LAYER M1 ;
        RECT 46.745 7.895 46.995 11.425 ;
  LAYER M1 ;
        RECT 46.745 11.675 46.995 12.685 ;
  LAYER M1 ;
        RECT 46.745 13.775 46.995 17.305 ;
  LAYER M1 ;
        RECT 46.745 17.555 46.995 18.565 ;
  LAYER M1 ;
        RECT 46.745 19.655 46.995 23.185 ;
  LAYER M1 ;
        RECT 46.745 23.435 46.995 24.445 ;
  LAYER M1 ;
        RECT 46.745 25.535 46.995 26.545 ;
  LAYER M1 ;
        RECT 47.175 7.895 47.425 11.425 ;
  LAYER M1 ;
        RECT 47.175 13.775 47.425 17.305 ;
  LAYER M1 ;
        RECT 47.175 19.655 47.425 23.185 ;
  LAYER M2 ;
        RECT 35.52 7.84 46.18 8.12 ;
  LAYER M2 ;
        RECT 35.52 12.04 47.04 12.32 ;
  LAYER M2 ;
        RECT 36.38 8.26 47.04 8.54 ;
  LAYER M2 ;
        RECT 35.09 8.68 47.47 8.96 ;
  LAYER M2 ;
        RECT 36.38 13.72 47.04 14 ;
  LAYER M2 ;
        RECT 35.52 17.92 47.04 18.2 ;
  LAYER M2 ;
        RECT 35.52 14.14 46.18 14.42 ;
  LAYER M2 ;
        RECT 35.09 14.56 47.47 14.84 ;
  LAYER M2 ;
        RECT 35.52 19.6 46.18 19.88 ;
  LAYER M2 ;
        RECT 35.52 23.8 47.04 24.08 ;
  LAYER M2 ;
        RECT 36.38 20.02 47.04 20.3 ;
  LAYER M2 ;
        RECT 35.52 25.9 47.04 26.18 ;
  LAYER M2 ;
        RECT 35.09 20.44 47.47 20.72 ;
  LAYER M3 ;
        RECT 40.71 7.82 40.99 24.1 ;
  LAYER M3 ;
        RECT 41.14 8.24 41.42 20.32 ;
  LAYER M3 ;
        RECT 41.57 8.66 41.85 26.2 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 11.425 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 12.685 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 11.425 ;
  LAYER M1 ;
        RECT 12.345 11.675 12.595 12.685 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 14.785 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 14.785 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 11.425 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 12.685 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 14.785 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.365 11.675 18.615 12.685 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 14.785 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M2 ;
        RECT 1.12 7.84 18.66 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 19.52 12.32 ;
  LAYER M2 ;
        RECT 1.12 14.14 19.52 14.42 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 12.34 ;
  LAYER M2 ;
        RECT 1.98 8.26 19.52 8.54 ;
  LAYER M2 ;
        RECT 0.69 8.68 19.95 8.96 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 30.405 3.695 30.655 7.225 ;
  LAYER M1 ;
        RECT 30.405 2.435 30.655 3.445 ;
  LAYER M1 ;
        RECT 30.405 0.335 30.655 1.345 ;
  LAYER M1 ;
        RECT 30.835 3.695 31.085 7.225 ;
  LAYER M1 ;
        RECT 31.265 3.695 31.515 7.225 ;
  LAYER M1 ;
        RECT 31.265 2.435 31.515 3.445 ;
  LAYER M1 ;
        RECT 31.265 0.335 31.515 1.345 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 33.845 3.695 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.845 2.435 34.095 3.445 ;
  LAYER M1 ;
        RECT 33.845 0.335 34.095 1.345 ;
  LAYER M1 ;
        RECT 34.275 3.695 34.525 7.225 ;
  LAYER M1 ;
        RECT 34.705 3.695 34.955 7.225 ;
  LAYER M1 ;
        RECT 34.705 2.435 34.955 3.445 ;
  LAYER M1 ;
        RECT 34.705 0.335 34.955 1.345 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M1 ;
        RECT 35.565 3.695 35.815 7.225 ;
  LAYER M1 ;
        RECT 35.565 2.435 35.815 3.445 ;
  LAYER M1 ;
        RECT 35.565 0.335 35.815 1.345 ;
  LAYER M1 ;
        RECT 35.995 3.695 36.245 7.225 ;
  LAYER M1 ;
        RECT 36.425 3.695 36.675 7.225 ;
  LAYER M1 ;
        RECT 36.425 2.435 36.675 3.445 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 1.345 ;
  LAYER M1 ;
        RECT 36.855 3.695 37.105 7.225 ;
  LAYER M1 ;
        RECT 37.285 3.695 37.535 7.225 ;
  LAYER M1 ;
        RECT 37.285 2.435 37.535 3.445 ;
  LAYER M1 ;
        RECT 37.285 0.335 37.535 1.345 ;
  LAYER M1 ;
        RECT 37.715 3.695 37.965 7.225 ;
  LAYER M1 ;
        RECT 38.145 3.695 38.395 7.225 ;
  LAYER M1 ;
        RECT 38.145 2.435 38.395 3.445 ;
  LAYER M1 ;
        RECT 38.145 0.335 38.395 1.345 ;
  LAYER M1 ;
        RECT 38.575 3.695 38.825 7.225 ;
  LAYER M1 ;
        RECT 39.005 3.695 39.255 7.225 ;
  LAYER M1 ;
        RECT 39.005 2.435 39.255 3.445 ;
  LAYER M1 ;
        RECT 39.005 0.335 39.255 1.345 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.865 2.435 40.115 3.445 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 1.345 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M2 ;
        RECT 28.64 0.7 40.16 0.98 ;
  LAYER M2 ;
        RECT 28.64 7 39.3 7.28 ;
  LAYER M2 ;
        RECT 29.5 6.58 40.16 6.86 ;
  LAYER M2 ;
        RECT 28.64 2.8 39.3 3.08 ;
  LAYER M2 ;
        RECT 29.5 2.38 40.16 2.66 ;
  LAYER M2 ;
        RECT 28.21 6.16 40.59 6.44 ;
  END 
END CURRENT_MIRROR_OTA
