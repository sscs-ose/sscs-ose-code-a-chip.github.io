* SKY130 Spice File.
* Typical Varactor Parameters
.param
+ cnwvc_tox='41.6503*1'
+ cnwvc_cdepmult=1
+ cnwvc_cintmult=1
+ cnwvc_vt1=0.3333
+ cnwvc_vt2=0.2380952
+ cnwvc_vtr=0.16
+ cnwvc_dwc=0.0
+ cnwvc_dlc=0.0
+ cnwvc_dld=0.0
+ cnwvc2_tox='41.7642*1'
+ cnwvc2_cdepmult=1
+ cnwvc2_cintmult=1
+ cnwvc2_vt1=0.2
+ cnwvc2_vt2=0.33
+ cnwvc2_vtr=0.14
+ cnwvc2_dwc=0.0
+ cnwvc2_dlc=0.0
+ cnwvc2_dld=0.0
* sky130_fd_pr__model__parasitic__diode_ps2nw Parameters
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 1.000    $ Units: farad/meter^2
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 1.000    $ Units: farad/meter^2
* sky130_fd_pr__model__parasitic__diode_ps2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult = 1.000       $ Units: farad/meter
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 1.000       $ Units: farad/meter
* sky130_fd_pr__model__parasitic__diode_pw2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 1.0       $ Units: farad/meter
+ sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult = 1.0       $ Units: farad/meter
* sky130_fd_pr__diode_pw2nd_05v5  Parameters
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 1.0
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 1.0
* sky130_fd_pr__diode_pd2nw_05v5_hvt  Parameters
+ sky130_fd_pr__pfet_01v8_hvt__ajunction_mult = 1.0
+ sky130_fd_pr__pfet_01v8_hvt__pjunction_mult = 1.0
+ dkispp=1.000 dkbfpp=1.000 dknfpp = 1.000
+ dkispp5x=1.000 dkbfpp5x=1.000 dknfpp5x = 1.000 dkisepp5x=1.000
+ cvpp2_nhvnative10x4_cor=1.00
+ cvpp2_nhvnative10x4_sub=4.82e-15
+ cvpp2_phv5x4_cor=1.00
+ cvpp2_phv5x4_sub=4.82e-15
