# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_npn_05v5_W1p00L4p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_npn_05v5_W1p00L4p00 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  9.700000 BY  12.70000 ;
  OBS
    LAYER li1 ;
      RECT 0.170000  0.170000 9.790000  0.500000 ;
      RECT 0.170000  0.500000 0.500000 12.460000 ;
      RECT 0.170000 12.460000 9.790000 12.790000 ;
      RECT 1.300000  1.300000 8.660000  1.630000 ;
      RECT 1.300000  1.630000 1.630000 11.330000 ;
      RECT 1.300000 11.330000 8.660000 11.660000 ;
      RECT 3.310000  3.310000 6.650000  3.640000 ;
      RECT 3.310000  3.640000 3.640000  9.320000 ;
      RECT 3.310000  9.320000 6.650000  9.650000 ;
      RECT 4.475000  4.475000 5.485000  8.485000 ;
      RECT 6.320000  3.640000 6.650000  9.320000 ;
      RECT 8.330000  1.630000 8.660000 11.330000 ;
      RECT 9.460000  0.500000 9.790000 12.460000 ;
    LAYER mcon ;
      RECT 0.250000  0.250000 0.420000  0.420000 ;
      RECT 0.250000  0.635000 0.420000  0.805000 ;
      RECT 0.250000  0.995000 0.420000  1.165000 ;
      RECT 0.250000  1.355000 0.420000  1.525000 ;
      RECT 0.250000  1.715000 0.420000  1.885000 ;
      RECT 0.250000  2.075000 0.420000  2.245000 ;
      RECT 0.250000  2.435000 0.420000  2.605000 ;
      RECT 0.250000  2.795000 0.420000  2.965000 ;
      RECT 0.250000  3.155000 0.420000  3.325000 ;
      RECT 0.250000  3.515000 0.420000  3.685000 ;
      RECT 0.250000  3.875000 0.420000  4.045000 ;
      RECT 0.250000  4.235000 0.420000  4.405000 ;
      RECT 0.250000  4.595000 0.420000  4.765000 ;
      RECT 0.250000  4.955000 0.420000  5.125000 ;
      RECT 0.250000  5.315000 0.420000  5.485000 ;
      RECT 0.250000  5.675000 0.420000  5.845000 ;
      RECT 0.250000  6.035000 0.420000  6.205000 ;
      RECT 0.250000  6.395000 0.420000  6.565000 ;
      RECT 0.250000  6.755000 0.420000  6.925000 ;
      RECT 0.250000  7.115000 0.420000  7.285000 ;
      RECT 0.250000  7.475000 0.420000  7.645000 ;
      RECT 0.250000  7.835000 0.420000  8.005000 ;
      RECT 0.250000  8.195000 0.420000  8.365000 ;
      RECT 0.250000  8.555000 0.420000  8.725000 ;
      RECT 0.250000  8.915000 0.420000  9.085000 ;
      RECT 0.250000  9.275000 0.420000  9.445000 ;
      RECT 0.250000  9.635000 0.420000  9.805000 ;
      RECT 0.250000  9.995000 0.420000 10.165000 ;
      RECT 0.250000 10.355000 0.420000 10.525000 ;
      RECT 0.250000 10.715000 0.420000 10.885000 ;
      RECT 0.250000 11.075000 0.420000 11.245000 ;
      RECT 0.250000 11.435000 0.420000 11.605000 ;
      RECT 0.250000 11.795000 0.420000 11.965000 ;
      RECT 0.250000 12.155000 0.420000 12.325000 ;
      RECT 0.250000 12.540000 0.420000 12.710000 ;
      RECT 0.755000  0.250000 0.925000  0.420000 ;
      RECT 0.755000 12.540000 0.925000 12.710000 ;
      RECT 1.115000  0.250000 1.285000  0.420000 ;
      RECT 1.115000 12.540000 1.285000 12.710000 ;
      RECT 1.380000  1.380000 1.550000  1.550000 ;
      RECT 1.380000  1.895000 1.550000  2.065000 ;
      RECT 1.380000  2.255000 1.550000  2.425000 ;
      RECT 1.380000  2.615000 1.550000  2.785000 ;
      RECT 1.380000  2.975000 1.550000  3.145000 ;
      RECT 1.380000  3.335000 1.550000  3.505000 ;
      RECT 1.380000  3.695000 1.550000  3.865000 ;
      RECT 1.380000  4.055000 1.550000  4.225000 ;
      RECT 1.380000  4.415000 1.550000  4.585000 ;
      RECT 1.380000  4.775000 1.550000  4.945000 ;
      RECT 1.380000  5.135000 1.550000  5.305000 ;
      RECT 1.380000  5.495000 1.550000  5.665000 ;
      RECT 1.380000  5.855000 1.550000  6.025000 ;
      RECT 1.380000  6.215000 1.550000  6.385000 ;
      RECT 1.380000  6.575000 1.550000  6.745000 ;
      RECT 1.380000  6.935000 1.550000  7.105000 ;
      RECT 1.380000  7.295000 1.550000  7.465000 ;
      RECT 1.380000  7.655000 1.550000  7.825000 ;
      RECT 1.380000  8.015000 1.550000  8.185000 ;
      RECT 1.380000  8.375000 1.550000  8.545000 ;
      RECT 1.380000  8.735000 1.550000  8.905000 ;
      RECT 1.380000  9.095000 1.550000  9.265000 ;
      RECT 1.380000  9.455000 1.550000  9.625000 ;
      RECT 1.380000  9.815000 1.550000  9.985000 ;
      RECT 1.380000 10.175000 1.550000 10.345000 ;
      RECT 1.380000 10.535000 1.550000 10.705000 ;
      RECT 1.380000 10.895000 1.550000 11.065000 ;
      RECT 1.380000 11.410000 1.550000 11.580000 ;
      RECT 1.475000  0.250000 1.645000  0.420000 ;
      RECT 1.475000 12.540000 1.645000 12.710000 ;
      RECT 1.835000  0.250000 2.005000  0.420000 ;
      RECT 1.835000  1.380000 2.005000  1.550000 ;
      RECT 1.835000 11.410000 2.005000 11.580000 ;
      RECT 1.835000 12.540000 2.005000 12.710000 ;
      RECT 2.195000  0.250000 2.365000  0.420000 ;
      RECT 2.195000  1.380000 2.365000  1.550000 ;
      RECT 2.195000 11.410000 2.365000 11.580000 ;
      RECT 2.195000 12.540000 2.365000 12.710000 ;
      RECT 2.555000  0.250000 2.725000  0.420000 ;
      RECT 2.555000  1.380000 2.725000  1.550000 ;
      RECT 2.555000 11.410000 2.725000 11.580000 ;
      RECT 2.555000 12.540000 2.725000 12.710000 ;
      RECT 2.915000  0.250000 3.085000  0.420000 ;
      RECT 2.915000  1.380000 3.085000  1.550000 ;
      RECT 2.915000 11.410000 3.085000 11.580000 ;
      RECT 2.915000 12.540000 3.085000 12.710000 ;
      RECT 3.275000  0.250000 3.445000  0.420000 ;
      RECT 3.275000  1.380000 3.445000  1.550000 ;
      RECT 3.275000 11.410000 3.445000 11.580000 ;
      RECT 3.275000 12.540000 3.445000 12.710000 ;
      RECT 3.390000  3.390000 3.560000  3.560000 ;
      RECT 3.390000  3.875000 3.560000  4.045000 ;
      RECT 3.390000  4.235000 3.560000  4.405000 ;
      RECT 3.390000  4.595000 3.560000  4.765000 ;
      RECT 3.390000  4.955000 3.560000  5.125000 ;
      RECT 3.390000  5.315000 3.560000  5.485000 ;
      RECT 3.390000  5.675000 3.560000  5.845000 ;
      RECT 3.390000  6.035000 3.560000  6.205000 ;
      RECT 3.390000  6.395000 3.560000  6.565000 ;
      RECT 3.390000  6.755000 3.560000  6.925000 ;
      RECT 3.390000  7.115000 3.560000  7.285000 ;
      RECT 3.390000  7.475000 3.560000  7.645000 ;
      RECT 3.390000  7.835000 3.560000  8.005000 ;
      RECT 3.390000  8.195000 3.560000  8.365000 ;
      RECT 3.390000  8.555000 3.560000  8.725000 ;
      RECT 3.390000  8.915000 3.560000  9.085000 ;
      RECT 3.390000  9.400000 3.560000  9.570000 ;
      RECT 3.635000  0.250000 3.805000  0.420000 ;
      RECT 3.635000  1.380000 3.805000  1.550000 ;
      RECT 3.635000 11.410000 3.805000 11.580000 ;
      RECT 3.635000 12.540000 3.805000 12.710000 ;
      RECT 3.815000  3.390000 3.985000  3.560000 ;
      RECT 3.815000  9.400000 3.985000  9.570000 ;
      RECT 3.995000  0.250000 4.165000  0.420000 ;
      RECT 3.995000  1.380000 4.165000  1.550000 ;
      RECT 3.995000 11.410000 4.165000 11.580000 ;
      RECT 3.995000 12.540000 4.165000 12.710000 ;
      RECT 4.175000  3.390000 4.345000  3.560000 ;
      RECT 4.175000  9.400000 4.345000  9.570000 ;
      RECT 4.355000  0.250000 4.525000  0.420000 ;
      RECT 4.355000  1.380000 4.525000  1.550000 ;
      RECT 4.355000 11.410000 4.525000 11.580000 ;
      RECT 4.355000 12.540000 4.525000 12.710000 ;
      RECT 4.535000  3.390000 4.705000  3.560000 ;
      RECT 4.535000  4.595000 5.425000  8.365000 ;
      RECT 4.535000  9.400000 4.705000  9.570000 ;
      RECT 4.715000  0.250000 4.885000  0.420000 ;
      RECT 4.715000  1.380000 4.885000  1.550000 ;
      RECT 4.715000 11.410000 4.885000 11.580000 ;
      RECT 4.715000 12.540000 4.885000 12.710000 ;
      RECT 4.895000  3.390000 5.065000  3.560000 ;
      RECT 4.895000  9.400000 5.065000  9.570000 ;
      RECT 5.075000  0.250000 5.245000  0.420000 ;
      RECT 5.075000  1.380000 5.245000  1.550000 ;
      RECT 5.075000 11.410000 5.245000 11.580000 ;
      RECT 5.075000 12.540000 5.245000 12.710000 ;
      RECT 5.255000  3.390000 5.425000  3.560000 ;
      RECT 5.255000  9.400000 5.425000  9.570000 ;
      RECT 5.435000  0.250000 5.605000  0.420000 ;
      RECT 5.435000  1.380000 5.605000  1.550000 ;
      RECT 5.435000 11.410000 5.605000 11.580000 ;
      RECT 5.435000 12.540000 5.605000 12.710000 ;
      RECT 5.615000  3.390000 5.785000  3.560000 ;
      RECT 5.615000  9.400000 5.785000  9.570000 ;
      RECT 5.795000  0.250000 5.965000  0.420000 ;
      RECT 5.795000  1.380000 5.965000  1.550000 ;
      RECT 5.795000 11.410000 5.965000 11.580000 ;
      RECT 5.795000 12.540000 5.965000 12.710000 ;
      RECT 5.975000  3.390000 6.145000  3.560000 ;
      RECT 5.975000  9.400000 6.145000  9.570000 ;
      RECT 6.155000  0.250000 6.325000  0.420000 ;
      RECT 6.155000  1.380000 6.325000  1.550000 ;
      RECT 6.155000 11.410000 6.325000 11.580000 ;
      RECT 6.155000 12.540000 6.325000 12.710000 ;
      RECT 6.400000  3.390000 6.570000  3.560000 ;
      RECT 6.400000  3.875000 6.570000  4.045000 ;
      RECT 6.400000  4.235000 6.570000  4.405000 ;
      RECT 6.400000  4.595000 6.570000  4.765000 ;
      RECT 6.400000  4.955000 6.570000  5.125000 ;
      RECT 6.400000  5.315000 6.570000  5.485000 ;
      RECT 6.400000  5.675000 6.570000  5.845000 ;
      RECT 6.400000  6.035000 6.570000  6.205000 ;
      RECT 6.400000  6.395000 6.570000  6.565000 ;
      RECT 6.400000  6.755000 6.570000  6.925000 ;
      RECT 6.400000  7.115000 6.570000  7.285000 ;
      RECT 6.400000  7.475000 6.570000  7.645000 ;
      RECT 6.400000  7.835000 6.570000  8.005000 ;
      RECT 6.400000  8.195000 6.570000  8.365000 ;
      RECT 6.400000  8.555000 6.570000  8.725000 ;
      RECT 6.400000  8.915000 6.570000  9.085000 ;
      RECT 6.400000  9.400000 6.570000  9.570000 ;
      RECT 6.515000  0.250000 6.685000  0.420000 ;
      RECT 6.515000  1.380000 6.685000  1.550000 ;
      RECT 6.515000 11.410000 6.685000 11.580000 ;
      RECT 6.515000 12.540000 6.685000 12.710000 ;
      RECT 6.875000  0.250000 7.045000  0.420000 ;
      RECT 6.875000  1.380000 7.045000  1.550000 ;
      RECT 6.875000 11.410000 7.045000 11.580000 ;
      RECT 6.875000 12.540000 7.045000 12.710000 ;
      RECT 7.235000  0.250000 7.405000  0.420000 ;
      RECT 7.235000  1.380000 7.405000  1.550000 ;
      RECT 7.235000 11.410000 7.405000 11.580000 ;
      RECT 7.235000 12.540000 7.405000 12.710000 ;
      RECT 7.595000  0.250000 7.765000  0.420000 ;
      RECT 7.595000  1.380000 7.765000  1.550000 ;
      RECT 7.595000 11.410000 7.765000 11.580000 ;
      RECT 7.595000 12.540000 7.765000 12.710000 ;
      RECT 7.955000  0.250000 8.125000  0.420000 ;
      RECT 7.955000  1.380000 8.125000  1.550000 ;
      RECT 7.955000 11.410000 8.125000 11.580000 ;
      RECT 7.955000 12.540000 8.125000 12.710000 ;
      RECT 8.315000  0.250000 8.485000  0.420000 ;
      RECT 8.315000 12.540000 8.485000 12.710000 ;
      RECT 8.410000  1.380000 8.580000  1.550000 ;
      RECT 8.410000  1.895000 8.580000  2.065000 ;
      RECT 8.410000  2.255000 8.580000  2.425000 ;
      RECT 8.410000  2.615000 8.580000  2.785000 ;
      RECT 8.410000  2.975000 8.580000  3.145000 ;
      RECT 8.410000  3.335000 8.580000  3.505000 ;
      RECT 8.410000  3.695000 8.580000  3.865000 ;
      RECT 8.410000  4.055000 8.580000  4.225000 ;
      RECT 8.410000  4.415000 8.580000  4.585000 ;
      RECT 8.410000  4.775000 8.580000  4.945000 ;
      RECT 8.410000  5.135000 8.580000  5.305000 ;
      RECT 8.410000  5.495000 8.580000  5.665000 ;
      RECT 8.410000  5.855000 8.580000  6.025000 ;
      RECT 8.410000  6.215000 8.580000  6.385000 ;
      RECT 8.410000  6.575000 8.580000  6.745000 ;
      RECT 8.410000  6.935000 8.580000  7.105000 ;
      RECT 8.410000  7.295000 8.580000  7.465000 ;
      RECT 8.410000  7.655000 8.580000  7.825000 ;
      RECT 8.410000  8.015000 8.580000  8.185000 ;
      RECT 8.410000  8.375000 8.580000  8.545000 ;
      RECT 8.410000  8.735000 8.580000  8.905000 ;
      RECT 8.410000  9.095000 8.580000  9.265000 ;
      RECT 8.410000  9.455000 8.580000  9.625000 ;
      RECT 8.410000  9.815000 8.580000  9.985000 ;
      RECT 8.410000 10.175000 8.580000 10.345000 ;
      RECT 8.410000 10.535000 8.580000 10.705000 ;
      RECT 8.410000 10.895000 8.580000 11.065000 ;
      RECT 8.410000 11.410000 8.580000 11.580000 ;
      RECT 8.675000  0.250000 8.845000  0.420000 ;
      RECT 8.675000 12.540000 8.845000 12.710000 ;
      RECT 9.035000  0.250000 9.205000  0.420000 ;
      RECT 9.035000 12.540000 9.205000 12.710000 ;
      RECT 9.540000  0.250000 9.710000  0.420000 ;
      RECT 9.540000  0.635000 9.710000  0.805000 ;
      RECT 9.540000  0.995000 9.710000  1.165000 ;
      RECT 9.540000  1.355000 9.710000  1.525000 ;
      RECT 9.540000  1.715000 9.710000  1.885000 ;
      RECT 9.540000  2.075000 9.710000  2.245000 ;
      RECT 9.540000  2.435000 9.710000  2.605000 ;
      RECT 9.540000  2.795000 9.710000  2.965000 ;
      RECT 9.540000  3.155000 9.710000  3.325000 ;
      RECT 9.540000  3.515000 9.710000  3.685000 ;
      RECT 9.540000  3.875000 9.710000  4.045000 ;
      RECT 9.540000  4.235000 9.710000  4.405000 ;
      RECT 9.540000  4.595000 9.710000  4.765000 ;
      RECT 9.540000  4.955000 9.710000  5.125000 ;
      RECT 9.540000  5.315000 9.710000  5.485000 ;
      RECT 9.540000  5.675000 9.710000  5.845000 ;
      RECT 9.540000  6.035000 9.710000  6.205000 ;
      RECT 9.540000  6.395000 9.710000  6.565000 ;
      RECT 9.540000  6.755000 9.710000  6.925000 ;
      RECT 9.540000  7.115000 9.710000  7.285000 ;
      RECT 9.540000  7.475000 9.710000  7.645000 ;
      RECT 9.540000  7.835000 9.710000  8.005000 ;
      RECT 9.540000  8.195000 9.710000  8.365000 ;
      RECT 9.540000  8.555000 9.710000  8.725000 ;
      RECT 9.540000  8.915000 9.710000  9.085000 ;
      RECT 9.540000  9.275000 9.710000  9.445000 ;
      RECT 9.540000  9.635000 9.710000  9.805000 ;
      RECT 9.540000  9.995000 9.710000 10.165000 ;
      RECT 9.540000 10.355000 9.710000 10.525000 ;
      RECT 9.540000 10.715000 9.710000 10.885000 ;
      RECT 9.540000 11.075000 9.710000 11.245000 ;
      RECT 9.540000 11.435000 9.710000 11.605000 ;
      RECT 9.540000 11.795000 9.710000 11.965000 ;
      RECT 9.540000 12.155000 9.710000 12.325000 ;
      RECT 9.540000 12.540000 9.710000 12.710000 ;
    LAYER met1 ;
      RECT 0.190000  0.190000 9.770000  0.480000 ;
      RECT 0.190000  0.480000 0.480000 12.480000 ;
      RECT 0.190000 12.480000 9.770000 12.770000 ;
      RECT 1.320000  1.320000 8.640000  1.610000 ;
      RECT 1.320000  1.610000 1.610000 11.350000 ;
      RECT 1.320000 11.350000 8.640000 11.640000 ;
      RECT 3.330000  3.330000 6.630000  3.620000 ;
      RECT 3.330000  3.620000 3.620000  9.340000 ;
      RECT 3.330000  9.340000 6.630000  9.630000 ;
      RECT 4.475000  4.535000 5.485000  8.425000 ;
      RECT 6.340000  3.620000 6.630000  9.340000 ;
      RECT 8.350000  1.610000 8.640000 11.350000 ;
      RECT 9.480000  0.480000 9.770000 12.480000 ;
  END
END sky130_fd_pr__rf_npn_05v5_W1p00L4p00
END LIBRARY
