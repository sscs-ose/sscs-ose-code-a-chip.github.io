magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -276 -1779 276 1779
<< nmos >>
rect -80 -1631 80 1569
<< ndiff >>
rect -138 1557 -80 1569
rect -138 -1619 -126 1557
rect -92 -1619 -80 1557
rect -138 -1631 -80 -1619
rect 80 1557 138 1569
rect 80 -1619 92 1557
rect 126 -1619 138 1557
rect 80 -1631 138 -1619
<< ndiffc >>
rect -126 -1619 -92 1557
rect 92 -1619 126 1557
<< psubdiff >>
rect -240 1709 -144 1743
rect 144 1709 240 1743
rect -240 1647 -206 1709
rect 206 1647 240 1709
rect -240 -1709 -206 -1647
rect 206 -1709 240 -1647
rect -240 -1743 -144 -1709
rect 144 -1743 240 -1709
<< psubdiffcont >>
rect -144 1709 144 1743
rect -240 -1647 -206 1647
rect 206 -1647 240 1647
rect -144 -1743 144 -1709
<< poly >>
rect -80 1641 80 1657
rect -80 1607 -64 1641
rect 64 1607 80 1641
rect -80 1569 80 1607
rect -80 -1657 80 -1631
<< polycont >>
rect -64 1607 64 1641
<< locali >>
rect -240 1709 -144 1743
rect 144 1709 240 1743
rect -240 1647 -206 1709
rect 206 1647 240 1709
rect -80 1607 -64 1641
rect 64 1607 80 1641
rect -126 1557 -92 1573
rect -126 -1635 -92 -1619
rect 92 1557 126 1573
rect 92 -1635 126 -1619
rect -240 -1709 -206 -1647
rect 206 -1709 240 -1647
rect -240 -1743 -144 -1709
rect 144 -1743 240 -1709
<< viali >>
rect -64 1607 64 1641
rect -126 -1619 -92 1557
rect 92 -1619 126 1557
<< metal1 >>
rect -76 1641 76 1647
rect -76 1607 -64 1641
rect 64 1607 76 1641
rect -76 1601 76 1607
rect -132 1557 -86 1569
rect -132 -1619 -126 1557
rect -92 -1619 -86 1557
rect -132 -1631 -86 -1619
rect 86 1557 132 1569
rect 86 -1619 92 1557
rect 126 -1619 132 1557
rect 86 -1631 132 -1619
<< labels >>
rlabel psubdiffcont 0 -1726 0 -1726 0 B
port 1 nsew
rlabel ndiffc -109 -31 -109 -31 0 D
port 2 nsew
rlabel ndiffc 109 -31 109 -31 0 S
port 3 nsew
rlabel polycont 0 1624 0 1624 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -223 -1726 223 1726
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 16.0 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
