MACRO NMOS_S_7151189_X6_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_7151189_X6_Y2 0 0 ;
  SIZE 6880 BY 13440 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 260 3150 6460 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3300 4460 3580 10660 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3730 680 4010 12760 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 13105 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 13105 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 13105 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 13105 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 13105 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 13105 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M2 ;
      RECT 1120 280 5760 560 ;
    LAYER M2 ;
      RECT 1120 4480 5760 4760 ;
    LAYER M2 ;
      RECT 690 700 6190 980 ;
    LAYER M2 ;
      RECT 1120 6160 5760 6440 ;
    LAYER M2 ;
      RECT 1120 10360 5760 10640 ;
    LAYER M2 ;
      RECT 690 6580 6190 6860 ;
    LAYER M2 ;
      RECT 1120 12460 5760 12740 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12515 1375 12685 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12515 2235 12685 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12515 3095 12685 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12515 3955 12685 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12515 4815 12685 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12515 5675 12685 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V2 ;
      RECT 2935 345 3085 495 ;
    LAYER V2 ;
      RECT 2935 6225 3085 6375 ;
    LAYER V2 ;
      RECT 3365 4545 3515 4695 ;
    LAYER V2 ;
      RECT 3365 10425 3515 10575 ;
    LAYER V2 ;
      RECT 3795 765 3945 915 ;
    LAYER V2 ;
      RECT 3795 6645 3945 6795 ;
    LAYER V2 ;
      RECT 3795 12525 3945 12675 ;
  END
END NMOS_S_7151189_X6_Y2
