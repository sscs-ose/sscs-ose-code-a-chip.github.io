VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO myconfig
   CLASS BLOCK ;
   SIZE 276.46 BY 217.3 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.24 0.0 63.62 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  68.68 0.0 69.06 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  74.12 0.0 74.5 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.36 0.0 86.74 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.8 0.0 92.18 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.24 0.0 97.62 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.36 0.0 103.74 1.06 ;
      END
   END din0[7]
   PIN din1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 216.24 163.58 217.3 ;
      END
   END din1[0]
   PIN din1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 216.24 169.02 217.3 ;
      END
   END din1[1]
   PIN din1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 216.24 174.46 217.3 ;
      END
   END din1[2]
   PIN din1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 216.24 179.9 217.3 ;
      END
   END din1[3]
   PIN din1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 216.24 186.7 217.3 ;
      END
   END din1[4]
   PIN din1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 216.24 192.14 217.3 ;
      END
   END din1[5]
   PIN din1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 216.24 197.58 217.3 ;
      END
   END din1[6]
   PIN din1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 216.24 204.38 217.3 ;
      END
   END din1[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  56.44 0.0 56.82 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 111.52 1.06 111.9 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 119.68 1.06 120.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 125.8 1.06 126.18 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 133.28 1.06 133.66 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.72 1.06 139.1 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 216.24 213.22 217.3 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 73.44 276.46 73.82 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 65.28 276.46 65.66 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 61.2 276.46 61.58 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 50.32 276.46 50.7 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 45.56 276.46 45.94 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 19.04 1.06 19.42 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 197.88 276.46 198.26 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 27.2 1.06 27.58 ;
      END
   END web0
   PIN web1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  275.4 190.4 276.46 190.78 ;
      END
   END web1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.28 0.0 31.66 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 216.24 245.18 217.3 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  112.88 0.0 113.26 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 0.0 120.06 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  125.8 0.0 126.18 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  131.92 0.0 132.3 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 0.0 144.54 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 0.0 157.46 1.06 ;
      END
   END dout0[7]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  112.88 216.24 113.26 217.3 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 216.24 120.06 217.3 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  125.8 216.24 126.18 217.3 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  131.92 216.24 132.3 217.3 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 216.24 138.42 217.3 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 216.24 144.54 217.3 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 216.24 150.66 217.3 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 216.24 157.46 217.3 ;
      END
   END dout1[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  271.32 3.4 273.06 213.9 ;
         LAYER met3 ;
         RECT  3.4 3.4 273.06 5.14 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 213.9 ;
         LAYER met3 ;
         RECT  3.4 212.16 273.06 213.9 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 276.46 1.74 ;
         LAYER met4 ;
         RECT  274.72 0.0 276.46 217.3 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 217.3 ;
         LAYER met3 ;
         RECT  0.0 215.56 276.46 217.3 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 275.84 216.68 ;
   LAYER  met2 ;
      RECT  0.62 0.62 275.84 216.68 ;
   LAYER  met3 ;
      RECT  1.66 110.92 275.84 112.5 ;
      RECT  0.62 112.5 1.66 119.08 ;
      RECT  0.62 120.66 1.66 125.2 ;
      RECT  0.62 126.78 1.66 132.68 ;
      RECT  0.62 134.26 1.66 138.12 ;
      RECT  1.66 72.84 274.8 74.42 ;
      RECT  1.66 74.42 274.8 110.92 ;
      RECT  274.8 74.42 275.84 110.92 ;
      RECT  274.8 66.26 275.84 72.84 ;
      RECT  274.8 62.18 275.84 64.68 ;
      RECT  274.8 51.3 275.84 60.6 ;
      RECT  274.8 46.54 275.84 49.72 ;
      RECT  1.66 112.5 274.8 197.28 ;
      RECT  1.66 197.28 274.8 198.86 ;
      RECT  0.62 20.02 1.66 26.6 ;
      RECT  0.62 28.18 1.66 110.92 ;
      RECT  274.8 112.5 275.84 189.8 ;
      RECT  274.8 191.38 275.84 197.28 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 72.84 ;
      RECT  2.8 5.74 273.66 72.84 ;
      RECT  273.66 2.8 274.8 5.74 ;
      RECT  273.66 5.74 274.8 72.84 ;
      RECT  1.66 198.86 2.8 211.56 ;
      RECT  1.66 211.56 2.8 214.5 ;
      RECT  2.8 198.86 273.66 211.56 ;
      RECT  273.66 198.86 274.8 211.56 ;
      RECT  273.66 211.56 274.8 214.5 ;
      RECT  274.8 2.34 275.84 44.96 ;
      RECT  0.62 2.34 1.66 18.44 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 273.66 2.8 ;
      RECT  273.66 2.34 274.8 2.8 ;
      RECT  0.62 139.7 1.66 214.96 ;
      RECT  274.8 198.86 275.84 214.96 ;
      RECT  1.66 214.5 2.8 214.96 ;
      RECT  2.8 214.5 273.66 214.96 ;
      RECT  273.66 214.5 274.8 214.96 ;
   LAYER  met4 ;
      RECT  62.64 1.66 64.22 216.68 ;
      RECT  64.22 0.62 68.08 1.66 ;
      RECT  69.66 0.62 73.52 1.66 ;
      RECT  75.1 0.62 79.64 1.66 ;
      RECT  81.22 0.62 85.76 1.66 ;
      RECT  87.34 0.62 91.2 1.66 ;
      RECT  92.78 0.62 96.64 1.66 ;
      RECT  98.22 0.62 102.76 1.66 ;
      RECT  64.22 1.66 162.6 215.64 ;
      RECT  162.6 1.66 164.18 215.64 ;
      RECT  164.18 215.64 168.04 216.68 ;
      RECT  169.62 215.64 173.48 216.68 ;
      RECT  175.06 215.64 178.92 216.68 ;
      RECT  180.5 215.64 185.72 216.68 ;
      RECT  187.3 215.64 191.16 216.68 ;
      RECT  192.74 215.64 196.6 216.68 ;
      RECT  198.18 215.64 203.4 216.68 ;
      RECT  57.42 0.62 62.64 1.66 ;
      RECT  204.98 215.64 212.24 216.68 ;
      RECT  32.26 0.62 55.84 1.66 ;
      RECT  213.82 215.64 244.2 216.68 ;
      RECT  104.34 0.62 112.28 1.66 ;
      RECT  113.86 0.62 119.08 1.66 ;
      RECT  120.66 0.62 125.2 1.66 ;
      RECT  126.78 0.62 131.32 1.66 ;
      RECT  132.9 0.62 137.44 1.66 ;
      RECT  139.02 0.62 143.56 1.66 ;
      RECT  145.14 0.62 149.68 1.66 ;
      RECT  151.26 0.62 156.48 1.66 ;
      RECT  64.22 215.64 112.28 216.68 ;
      RECT  113.86 215.64 119.08 216.68 ;
      RECT  120.66 215.64 125.2 216.68 ;
      RECT  126.78 215.64 131.32 216.68 ;
      RECT  132.9 215.64 137.44 216.68 ;
      RECT  139.02 215.64 143.56 216.68 ;
      RECT  145.14 215.64 149.68 216.68 ;
      RECT  151.26 215.64 156.48 216.68 ;
      RECT  158.06 215.64 162.6 216.68 ;
      RECT  164.18 1.66 270.72 2.8 ;
      RECT  164.18 2.8 270.72 214.5 ;
      RECT  164.18 214.5 270.72 215.64 ;
      RECT  270.72 1.66 273.66 2.8 ;
      RECT  270.72 214.5 273.66 215.64 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 214.5 5.74 216.68 ;
      RECT  5.74 1.66 62.64 2.8 ;
      RECT  5.74 2.8 62.64 214.5 ;
      RECT  5.74 214.5 62.64 216.68 ;
      RECT  245.78 215.64 274.12 216.68 ;
      RECT  158.06 0.62 274.12 1.66 ;
      RECT  273.66 1.66 274.12 2.8 ;
      RECT  273.66 2.8 274.12 214.5 ;
      RECT  273.66 214.5 274.12 215.64 ;
      RECT  2.34 0.62 30.68 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 214.5 ;
      RECT  2.34 214.5 2.8 216.68 ;
   END
END    myconfig
END    LIBRARY
