# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_test_coil2
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_test_coil2 ;
  ORIGIN  132.5000  132.5000 ;
  SIZE  270.0000 BY  265.0000 ;
  OBS
    LAYER met2 ;
      POLYGON  -9.575000   77.500000  -8.725000   77.500000 -8.725000   76.650000 ;
      POLYGON  -9.575000  107.500000  -8.725000  107.500000 -8.725000  106.650000 ;
      POLYGON  -8.725000 -121.650000  -8.725000 -122.500000 -9.575000 -122.500000 ;
      POLYGON  -8.725000  -91.650000  -8.725000  -92.500000 -9.575000  -92.500000 ;
      POLYGON  -8.725000   76.650000   5.425000   76.650000  5.425000   62.500000 ;
      POLYGON  -8.725000  106.650000   5.425000  106.650000  5.425000   92.500000 ;
      POLYGON  -5.425000 -121.650000   5.425000 -121.650000 -5.425000 -132.500000 ;
      POLYGON  -5.425000  -91.650000   5.425000  -91.650000 -5.425000 -102.500000 ;
      POLYGON  -5.425000   87.500000   5.425000   76.650000 -5.425000   76.650000 ;
      POLYGON  -5.425000  117.500000   5.425000  106.650000 -5.425000  106.650000 ;
      POLYGON   5.425000 -117.500000   9.575000 -117.500000  5.425000 -121.650000 ;
      POLYGON   5.425000 -107.500000   5.425000 -121.650000 -8.725000 -121.650000 ;
      POLYGON   5.425000  -87.500000   9.575000  -87.500000  5.425000  -91.650000 ;
      POLYGON   5.425000  -77.500000   5.425000  -91.650000 -8.725000  -91.650000 ;
      POLYGON   5.425000   76.650000   9.575000   72.500000  5.425000   72.500000 ;
      POLYGON   5.425000  106.650000   9.575000  102.500000  5.425000  102.500000 ;
      RECT -31.155000 -132.500000  -5.425000 -122.500000 ;
      RECT -31.155000 -102.500000  -5.425000  -92.500000 ;
      RECT -31.155000   77.500000  -5.425000   87.500000 ;
      RECT -31.155000  107.500000  -5.425000  117.500000 ;
      RECT  -8.725000 -122.500000  -5.425000 -121.650000 ;
      RECT  -8.725000  -92.500000  -5.425000  -91.650000 ;
      RECT  -8.725000   76.650000  -5.425000   77.500000 ;
      RECT  -8.725000  106.650000  -5.425000  107.500000 ;
      RECT   5.425000 -117.500000  30.040000 -107.500000 ;
      RECT   5.425000  -87.500000  30.040000  -77.500000 ;
      RECT   5.425000   62.500000  30.040000   72.500000 ;
      RECT   5.425000   92.500000  30.040000  102.500000 ;
      RECT  49.540000   -5.000000 137.500000    5.000000 ;
    LAYER met3 ;
      POLYGON -132.500000  -54.890000 -125.590000  -54.890000 -125.590000  -61.800000 ;
      POLYGON -125.590000  -61.800000 -118.360000  -61.800000 -118.360000  -69.030000 ;
      POLYGON -125.590000   61.800000 -125.590000   54.890000 -132.500000   54.890000 ;
      POLYGON -122.500000  -50.750000 -117.500000  -55.750000 -122.500000  -55.750000 ;
      POLYGON -122.500000   54.890000 -118.360000   54.890000 -122.500000   50.750000 ;
      POLYGON -119.245000   68.145000 -119.245000   61.800000 -125.590000   61.800000 ;
      POLYGON -118.360000  -69.030000 -111.450000  -69.030000 -111.450000  -75.940000 ;
      POLYGON -118.360000   60.940000 -112.310000   60.940000 -118.360000   54.890000 ;
      POLYGON -117.500000  -55.750000 -110.430000  -62.820000 -117.500000  -62.820000 ;
      POLYGON -117.500000  -48.680000 -115.430000  -48.680000 -115.430000  -50.750000 ;
      POLYGON -115.430000  -50.750000 -110.430000  -50.750000 -110.430000  -55.750000 ;
      POLYGON -115.430000   50.750000 -115.430000   48.680000 -117.500000   48.680000 ;
      POLYGON -112.310000   68.010000 -105.240000   68.010000 -112.310000   60.940000 ;
      POLYGON -111.450000  -75.940000 -104.220000  -75.940000 -104.220000  -83.170000 ;
      POLYGON -111.450000   75.940000 -111.450000   68.145000 -119.245000   68.145000 ;
      POLYGON -111.290000   54.890000 -111.290000   50.750000 -115.430000   50.750000 ;
      POLYGON -110.430000  -62.820000 -103.360000  -69.890000 -110.430000  -69.890000 ;
      POLYGON -110.430000  -55.750000 -103.360000  -55.750000 -103.360000  -62.820000 ;
      POLYGON -107.500000  -44.540000 -102.500000  -49.540000 -107.500000  -49.540000 ;
      POLYGON -107.500000   45.940000 -106.100000   45.940000 -107.500000   44.540000 ;
      POLYGON -106.100000   53.015000  -99.025000   53.015000 -106.100000   45.940000 ;
      POLYGON -105.240000   60.940000 -105.240000   54.890000 -111.290000   54.890000 ;
      POLYGON -105.240000   75.080000  -98.170000   75.080000 -105.240000   68.010000 ;
      POLYGON -104.245000   83.145000 -104.245000   75.940000 -111.450000   75.940000 ;
      POLYGON -104.220000  -83.170000  -97.310000  -83.170000  -97.310000  -90.080000 ;
      POLYGON -103.360000  -69.890000  -96.290000  -76.960000 -103.360000  -76.960000 ;
      POLYGON -103.360000  -62.820000  -96.290000  -62.820000  -96.290000  -69.890000 ;
      POLYGON -102.500000  -49.540000  -95.435000  -56.605000 -102.500000  -56.605000 ;
      POLYGON -102.500000  -42.465000 -100.425000  -42.465000 -100.425000  -44.540000 ;
      POLYGON -100.425000  -44.540000  -95.425000  -44.540000  -95.425000  -49.540000 ;
      POLYGON -100.425000   44.540000 -100.425000   42.465000 -102.500000   42.465000 ;
      POLYGON  -99.025000   45.940000  -99.025000   44.540000 -100.425000   44.540000 ;
      POLYGON  -99.025000   60.080000  -91.960000   60.080000  -99.025000   53.015000 ;
      POLYGON  -98.170000   68.010000  -98.170000   60.940000 -105.240000   60.940000 ;
      POLYGON  -98.170000   82.150000  -91.100000   82.150000  -98.170000   75.080000 ;
      POLYGON  -97.310000  -90.080000  -89.250000  -90.080000  -89.250000  -98.140000 ;
      POLYGON  -97.310000   90.080000  -97.310000   83.145000 -104.245000   83.145000 ;
      POLYGON  -96.290000  -76.960000  -89.220000  -84.030000  -96.290000  -84.030000 ;
      POLYGON  -96.290000  -69.890000  -89.220000  -69.890000  -89.220000  -76.960000 ;
      POLYGON  -95.435000  -56.605000  -88.360000  -63.680000  -95.435000  -63.680000 ;
      POLYGON  -95.425000  -49.540000  -88.360000  -49.540000  -88.360000  -56.605000 ;
      POLYGON  -92.500000  -38.325000  -87.500000  -43.325000  -92.500000  -43.325000 ;
      POLYGON  -92.500000   45.080000  -85.745000   45.080000  -92.500000   38.325000 ;
      POLYGON  -91.960000   67.155000  -84.885000   67.155000  -91.960000   60.080000 ;
      POLYGON  -91.950000   53.015000  -91.950000   45.940000  -99.025000   45.940000 ;
      POLYGON  -91.100000   75.080000  -91.100000   68.010000  -98.170000   68.010000 ;
      POLYGON  -91.100000   89.220000  -84.030000   89.220000  -91.100000   82.150000 ;
      POLYGON  -90.535000   96.855000  -90.535000   90.080000  -97.310000   90.080000 ;
      POLYGON  -89.250000  -98.140000  -83.170000  -98.140000  -83.170000 -104.220000 ;
      POLYGON  -89.220000  -84.030000  -82.150000  -91.100000  -89.220000  -91.100000 ;
      POLYGON  -89.220000  -76.960000  -82.150000  -76.960000  -82.150000  -84.030000 ;
      POLYGON  -88.360000  -63.680000  -81.295000  -70.745000  -88.360000  -70.745000 ;
      POLYGON  -88.360000  -56.605000  -81.285000  -56.605000  -81.285000  -63.680000 ;
      POLYGON  -87.500000  -43.325000  -80.430000  -50.395000  -87.500000  -50.395000 ;
      POLYGON  -87.500000  -36.255000  -85.430000  -36.255000  -85.430000  -38.325000 ;
      POLYGON  -85.745000   52.150000  -78.675000   52.150000  -85.745000   45.080000 ;
      POLYGON  -85.430000  -38.325000  -80.430000  -38.325000  -80.430000  -43.325000 ;
      POLYGON  -85.430000   38.325000  -85.430000   36.255000  -87.500000   36.255000 ;
      POLYGON  -84.885000   60.080000  -84.885000   53.015000  -91.950000   53.015000 ;
      POLYGON  -84.885000   74.220000  -77.820000   74.220000  -84.885000   67.155000 ;
      POLYGON  -84.315000   81.865000  -84.315000   75.080000  -91.100000   75.080000 ;
      POLYGON  -84.030000   82.150000  -84.030000   81.865000  -84.315000   81.865000 ;
      POLYGON  -84.030000   94.235000  -79.015000   94.235000  -84.030000   89.220000 ;
      POLYGON  -83.170000 -104.220000  -75.530000 -104.220000  -75.530000 -111.860000 ;
      POLYGON  -83.170000  104.220000  -83.170000   96.855000  -90.535000   96.855000 ;
      POLYGON  -82.150000  -91.100000  -75.080000  -98.170000  -82.150000  -98.170000 ;
      POLYGON  -82.150000  -84.030000  -75.080000  -84.030000  -75.080000  -91.100000 ;
      POLYGON  -81.295000  -70.745000  -74.220000  -77.820000  -81.295000  -77.820000 ;
      POLYGON  -81.285000  -63.680000  -74.220000  -63.680000  -74.220000  -70.745000 ;
      POLYGON  -80.430000  -50.395000  -73.360000  -57.465000  -80.430000  -57.465000 ;
      POLYGON  -80.430000  -43.325000  -73.360000  -43.325000  -73.360000  -50.395000 ;
      POLYGON  -79.215000   44.540000  -79.215000   38.325000  -85.430000   38.325000 ;
      POLYGON  -79.015000   99.475000  -73.775000   99.475000  -79.015000   94.235000 ;
      POLYGON  -78.675000   45.080000  -78.675000   44.540000  -79.215000   44.540000 ;
      POLYGON  -78.675000   59.220000  -71.605000   59.220000  -78.675000   52.150000 ;
      POLYGON  -78.100000   66.865000  -78.100000   60.080000  -84.885000   60.080000 ;
      POLYGON  -77.820000   81.295000  -70.745000   81.295000  -77.820000   74.220000 ;
      POLYGON  -77.810000   67.155000  -77.810000   66.865000  -78.100000   66.865000 ;
      POLYGON  -77.500000  -32.115000  -72.500000  -37.115000  -77.500000  -37.115000 ;
      POLYGON  -77.500000   37.155000  -72.460000   37.155000  -77.500000   32.115000 ;
      POLYGON  -76.960000   89.220000  -76.960000   82.150000  -84.030000   82.150000 ;
      POLYGON  -76.870000  110.520000  -76.870000  104.220000  -83.170000  104.220000 ;
      POLYGON  -75.530000 -111.860000  -69.030000 -111.860000  -69.030000 -118.360000 ;
      POLYGON  -75.080000  -98.170000  -68.010000 -105.240000  -75.080000 -105.240000 ;
      POLYGON  -75.080000  -91.100000  -68.010000  -91.100000  -68.010000  -98.170000 ;
      POLYGON  -74.220000  -77.820000  -67.155000  -84.885000  -74.220000  -84.885000 ;
      POLYGON  -74.220000  -70.745000  -67.145000  -70.745000  -67.145000  -77.820000 ;
      POLYGON  -73.775000  105.240000  -68.010000  105.240000  -73.775000   99.475000 ;
      POLYGON  -73.360000  -57.465000  -66.290000  -64.535000  -73.360000  -64.535000 ;
      POLYGON  -73.360000  -50.395000  -66.290000  -50.395000  -66.290000  -57.465000 ;
      POLYGON  -72.500000  -37.115000  -65.435000  -44.180000  -72.500000  -44.180000 ;
      POLYGON  -72.500000  -30.040000  -70.425000  -30.040000  -70.425000  -32.115000 ;
      POLYGON  -72.460000   30.080000  -72.460000   30.040000  -72.500000   30.040000 ;
      POLYGON  -72.460000   44.220000  -65.395000   44.220000  -72.460000   37.155000 ;
      POLYGON  -71.945000   94.235000  -71.945000   89.220000  -76.960000   89.220000 ;
      POLYGON  -71.605000   52.150000  -71.605000   45.080000  -78.675000   45.080000 ;
      POLYGON  -71.605000   66.290000  -64.535000   66.290000  -71.605000   59.220000 ;
      POLYGON  -70.745000   74.220000  -70.745000   67.155000  -77.810000   67.155000 ;
      POLYGON  -70.745000   88.360000  -63.680000   88.360000  -70.745000   81.295000 ;
      POLYGON  -70.665000   95.515000  -70.665000   94.235000  -71.945000   94.235000 ;
      POLYGON  -70.425000  -32.115000  -65.425000  -32.115000  -65.425000  -37.115000 ;
      POLYGON  -70.425000   32.115000  -70.425000   30.080000  -72.460000   30.080000 ;
      POLYGON  -69.030000 -118.360000  -54.890000 -118.360000  -54.890000 -132.500000 ;
      POLYGON  -69.030000  118.360000  -69.030000  110.520000  -76.870000  110.520000 ;
      POLYGON  -68.010000 -105.240000  -60.940000 -112.310000  -68.010000 -112.310000 ;
      POLYGON  -68.010000  -98.170000  -60.940000  -98.170000  -60.940000 -105.240000 ;
      POLYGON  -68.010000  111.450000  -61.800000  111.450000  -68.010000  105.240000 ;
      POLYGON  -67.155000  -84.885000  -60.080000  -91.960000  -67.155000  -91.960000 ;
      POLYGON  -67.145000  -77.820000  -60.080000  -77.820000  -60.080000  -84.885000 ;
      POLYGON  -66.705000   99.475000  -66.705000   95.515000  -70.665000   95.515000 ;
      POLYGON  -66.290000  -64.535000  -59.220000  -71.605000  -66.290000  -71.605000 ;
      POLYGON  -66.290000  -57.465000  -59.220000  -57.465000  -59.220000  -64.535000 ;
      POLYGON  -65.435000  -44.180000  -64.535000  -45.080000  -65.435000  -45.080000 ;
      POLYGON  -65.425000  -37.115000  -64.215000  -37.115000  -64.215000  -38.325000 ;
      POLYGON  -65.395000   51.295000  -58.320000   51.295000  -65.395000   44.220000 ;
      POLYGON  -65.385000   37.155000  -65.385000   32.115000  -70.425000   32.115000 ;
      POLYGON  -64.535000  -45.080000  -58.360000  -51.255000  -64.535000  -51.255000 ;
      POLYGON  -64.535000   59.220000  -64.535000   52.150000  -71.605000   52.150000 ;
      POLYGON  -64.535000   73.360000  -57.465000   73.360000  -64.535000   66.290000 ;
      POLYGON  -64.440000   80.525000  -64.440000   74.220000  -70.745000   74.220000 ;
      POLYGON  -64.215000  -38.325000  -58.360000  -38.325000  -58.360000  -44.180000 ;
      POLYGON  -63.680000   94.235000  -57.805000   94.235000  -63.680000   88.360000 ;
      POLYGON  -63.670000   81.295000  -63.670000   80.525000  -64.440000   80.525000 ;
      POLYGON  -62.820000  103.360000  -62.820000   99.475000  -66.705000   99.475000 ;
      POLYGON  -62.500000  -25.900000  -50.075000  -38.325000  -62.500000  -38.325000 ;
      POLYGON  -62.500000   30.080000  -58.320000   30.080000  -62.500000   25.900000 ;
      POLYGON  -61.800000  118.360000  -54.890000  118.360000  -61.800000  111.450000 ;
      POLYGON  -60.940000 -112.310000  -54.890000 -118.360000  -60.940000 -118.360000 ;
      POLYGON  -60.940000 -105.240000  -53.870000 -105.240000  -53.870000 -112.310000 ;
      POLYGON  -60.940000  105.240000  -60.940000  103.360000  -62.820000  103.360000 ;
      POLYGON  -60.080000  -91.960000  -53.015000  -99.025000  -60.080000  -99.025000 ;
      POLYGON  -60.080000  -84.885000  -53.005000  -84.885000  -53.005000  -91.960000 ;
      POLYGON  -59.220000  -71.605000  -52.150000  -78.675000  -59.220000  -78.675000 ;
      POLYGON  -59.220000  -64.535000  -52.150000  -64.535000  -52.150000  -71.605000 ;
      POLYGON  -58.360000  -51.255000  -51.295000  -58.320000  -58.360000  -58.320000 ;
      POLYGON  -58.360000  -44.180000  -57.460000  -44.180000  -57.460000  -45.080000 ;
      POLYGON  -58.320000   38.325000  -50.075000   38.325000  -58.320000   30.080000 ;
      POLYGON  -58.320000   44.220000  -58.320000   37.155000  -65.385000   37.155000 ;
      POLYGON  -58.320000   58.320000  -51.295000   58.320000  -58.320000   51.295000 ;
      POLYGON  -58.230000   65.525000  -58.230000   59.220000  -64.535000   59.220000 ;
      POLYGON  -57.805000  100.755000  -51.285000  100.755000  -57.805000   94.235000 ;
      POLYGON  -57.465000   66.290000  -57.465000   65.525000  -58.230000   65.525000 ;
      POLYGON  -57.465000   79.245000  -51.580000   79.245000  -57.465000   73.360000 ;
      POLYGON  -57.460000  -45.080000  -51.285000  -45.080000  -51.285000  -51.255000 ;
      POLYGON  -56.940000  109.240000  -56.940000  105.240000  -60.940000  105.240000 ;
      POLYGON  -56.605000   88.360000  -56.605000   81.295000  -63.670000   81.295000 ;
      POLYGON  -54.890000 -118.360000  -50.750000 -122.500000  -54.890000 -122.500000 ;
      POLYGON  -54.890000  122.500000  -50.750000  122.500000  -54.890000  118.360000 ;
      POLYGON  -54.890000  132.500000  -54.890000  118.360000  -69.030000  118.360000 ;
      POLYGON  -54.730000  111.450000  -54.730000  109.240000  -56.940000  109.240000 ;
      POLYGON  -53.870000 -112.310000  -48.680000 -112.310000  -48.680000 -117.500000 ;
      POLYGON  -53.015000  -99.025000  -46.800000 -105.240000  -53.015000 -105.240000 ;
      POLYGON  -53.005000  -91.960000  -45.940000  -91.960000  -45.940000  -99.025000 ;
      POLYGON  -52.150000  -78.675000  -45.080000  -85.745000  -52.150000  -85.745000 ;
      POLYGON  -52.150000  -71.605000  -45.080000  -71.605000  -45.080000  -78.675000 ;
      POLYGON  -51.580000   85.765000  -45.060000   85.765000  -51.580000   79.245000 ;
      POLYGON  -51.295000  -58.320000  -44.220000  -65.395000  -51.295000  -65.395000 ;
      POLYGON  -51.295000   64.245000  -45.370000   64.245000  -51.295000   58.320000 ;
      POLYGON  -51.285000  -51.255000  -44.220000  -51.255000  -44.220000  -58.320000 ;
      POLYGON  -51.285000  107.500000  -44.540000  107.500000  -51.285000  100.755000 ;
      POLYGON  -51.245000   51.295000  -51.245000   44.220000  -58.320000   44.220000 ;
      POLYGON  -50.730000   94.235000  -50.730000   88.360000  -56.605000   88.360000 ;
      POLYGON  -50.395000   73.360000  -50.395000   66.290000  -57.465000   66.290000 ;
      POLYGON  -50.075000  -38.325000  -37.650000  -50.750000  -50.075000  -50.750000 ;
      POLYGON  -50.075000   50.395000  -38.005000   50.395000  -50.075000   38.325000 ;
      POLYGON  -48.680000  117.500000  -48.680000  111.450000  -54.730000  111.450000 ;
      POLYGON  -46.800000 -105.240000  -44.540000 -107.500000  -46.800000 -107.500000 ;
      POLYGON  -45.940000  -99.025000  -42.465000  -99.025000  -42.465000 -102.500000 ;
      POLYGON  -45.370000   70.745000  -38.870000   70.745000  -45.370000   64.245000 ;
      POLYGON  -45.080000  -85.745000  -38.325000  -92.500000  -45.080000  -92.500000 ;
      POLYGON  -45.080000  -78.675000  -38.010000  -78.675000  -38.010000  -85.745000 ;
      POLYGON  -45.060000   92.500000  -38.325000   92.500000  -45.060000   85.765000 ;
      POLYGON  -44.510000   79.245000  -44.510000   73.360000  -50.395000   73.360000 ;
      POLYGON  -44.220000  -65.395000  -38.870000  -70.745000  -44.220000  -70.745000 ;
      POLYGON  -44.220000  -58.320000  -38.005000  -58.320000  -38.005000  -64.535000 ;
      POLYGON  -44.220000   58.320000  -44.220000   51.295000  -51.245000   51.295000 ;
      POLYGON  -44.210000  100.755000  -44.210000   94.235000  -50.730000   94.235000 ;
      POLYGON  -42.465000  102.500000  -42.465000  100.755000  -44.210000  100.755000 ;
      POLYGON  -38.870000  -70.745000  -32.115000  -77.500000  -38.870000  -77.500000 ;
      POLYGON  -38.870000   77.500000  -32.115000   77.500000  -38.870000   70.745000 ;
      POLYGON  -38.295000   64.245000  -38.295000   58.320000  -44.220000   58.320000 ;
      POLYGON  -38.010000  -85.745000  -36.255000  -85.745000  -36.255000  -87.500000 ;
      POLYGON  -38.005000  -64.535000  -37.145000  -64.535000  -37.145000  -65.395000 ;
      POLYGON  -38.005000   62.500000  -25.900000   62.500000  -38.005000   50.395000 ;
      POLYGON  -37.990000   85.765000  -37.990000   79.245000  -44.510000   79.245000 ;
      POLYGON  -37.650000  -50.750000  -25.900000  -62.500000  -37.650000  -62.500000 ;
      POLYGON  -37.145000  -65.395000  -31.795000  -65.395000  -31.795000  -70.745000 ;
      POLYGON  -36.255000   87.500000  -36.255000   85.765000  -37.990000   85.765000 ;
      POLYGON  -31.795000  -70.745000  -30.040000  -70.745000  -30.040000  -72.500000 ;
      POLYGON  -31.795000   70.745000  -31.795000   64.245000  -38.295000   64.245000 ;
      POLYGON  -30.040000   72.500000  -30.040000   70.745000  -31.795000   70.745000 ;
      POLYGON  -11.010000 -131.265000   -9.775000 -131.265000  -11.010000 -132.500000 ;
      POLYGON  -11.010000 -122.500000   -9.775000 -123.735000  -11.010000 -123.735000 ;
      POLYGON  -11.010000 -101.265000   -9.775000 -101.265000  -11.010000 -102.500000 ;
      POLYGON  -11.010000  -92.500000   -9.775000  -93.735000  -11.010000  -93.735000 ;
      POLYGON  -11.010000   78.735000   -9.775000   78.735000  -11.010000   77.500000 ;
      POLYGON  -11.010000   87.500000   -9.775000   86.265000  -11.010000   86.265000 ;
      POLYGON  -11.010000  108.735000   -9.775000  108.735000  -11.010000  107.500000 ;
      POLYGON  -11.010000  117.500000   -9.775000  116.265000  -11.010000  116.265000 ;
      POLYGON   -9.575000 -117.500000   -8.715000 -117.500000   -8.715000 -118.360000 ;
      POLYGON   -9.575000  -87.500000   -5.975000  -87.500000   -5.975000  -91.100000 ;
      POLYGON   -8.725000   73.350000   -8.725000   72.500000   -9.575000   72.500000 ;
      POLYGON   -8.725000  103.350000   -8.725000  102.500000   -9.575000  102.500000 ;
      POLYGON   -8.715000 -118.360000   -4.575000 -118.360000   -4.575000 -122.500000 ;
      POLYGON   -5.975000  -91.100000   -4.575000  -91.100000   -4.575000  -92.500000 ;
      POLYGON   -5.425000 -107.500000    5.435000 -118.360000   -5.425000 -118.360000 ;
      POLYGON   -5.425000  -77.500000    7.155000  -90.080000   -5.425000  -90.080000 ;
      POLYGON   -5.425000   73.350000    5.425000   73.350000   -5.425000   62.500000 ;
      POLYGON   -5.425000  103.350000    5.425000  103.350000   -5.425000   92.500000 ;
      POLYGON   -4.575000 -122.500000    5.425000 -122.500000    5.425000 -132.500000 ;
      POLYGON   -4.575000  -92.500000    5.425000  -92.500000    5.425000 -102.500000 ;
      POLYGON   -4.575000   77.500000   -4.575000   73.350000   -8.725000   73.350000 ;
      POLYGON   -4.575000  107.500000   -4.575000  103.350000   -8.725000  103.350000 ;
      POLYGON    5.425000   77.500000    9.575000   77.500000    5.425000   73.350000 ;
      POLYGON    5.425000   87.500000    5.425000   77.500000   -4.575000   77.500000 ;
      POLYGON    5.425000  107.500000    9.575000  107.500000    5.425000  103.350000 ;
      POLYGON    5.425000  117.500000    5.425000  107.500000   -4.575000  107.500000 ;
      POLYGON    5.435000 -118.360000    9.575000 -122.500000    5.435000 -122.500000 ;
      POLYGON    7.155000  -90.080000    9.575000  -92.500000    7.155000  -92.500000 ;
      POLYGON    8.660000 -116.265000    9.895000 -116.265000    9.895000 -117.500000 ;
      POLYGON    8.660000  -86.265000    9.895000  -86.265000    9.895000  -87.500000 ;
      POLYGON    8.660000   63.735000    9.895000   63.735000    9.895000   62.500000 ;
      POLYGON    8.660000   93.735000    9.895000   93.735000    9.895000   92.500000 ;
      POLYGON    9.895000 -107.500000    9.895000 -108.735000    8.660000 -108.735000 ;
      POLYGON    9.895000  -77.500000    9.895000  -78.735000    8.660000  -78.735000 ;
      POLYGON    9.895000   72.500000    9.895000   71.265000    8.660000   71.265000 ;
      POLYGON    9.895000  102.500000    9.895000  101.265000    8.660000  101.265000 ;
      POLYGON   25.900000   62.500000   38.005000   62.500000   38.005000   50.395000 ;
      POLYGON   30.040000  -69.030000   33.510000  -69.030000   30.040000  -72.500000 ;
      POLYGON   30.040000   72.500000   31.795000   70.745000   30.040000   70.745000 ;
      POLYGON   31.795000   70.745000   38.005000   64.535000   31.795000   64.535000 ;
      POLYGON   32.115000   77.500000   36.265000   77.500000   36.265000   73.350000 ;
      POLYGON   33.510000  -62.820000   39.720000  -62.820000   33.510000  -69.030000 ;
      POLYGON   33.675000  -75.940000   33.675000  -77.500000   32.115000  -77.500000 ;
      POLYGON   36.255000  -80.430000   43.325000  -80.430000   36.255000  -87.500000 ;
      POLYGON   36.255000   87.500000   38.010000   85.745000   36.255000   85.745000 ;
      POLYGON   36.265000   73.350000   37.115000   73.350000   37.115000   72.500000 ;
      POLYGON   37.115000  -72.500000   37.115000  -75.940000   33.675000  -75.940000 ;
      POLYGON   37.115000   72.500000   38.870000   72.500000   38.870000   70.745000 ;
      POLYGON   37.650000  -50.750000   37.650000  -62.500000   25.900000  -62.500000 ;
      POLYGON   38.005000  -50.395000   38.005000  -50.750000   37.650000  -50.750000 ;
      POLYGON   38.005000   50.395000   50.075000   50.395000   50.075000   38.325000 ;
      POLYGON   38.005000   64.535000   44.220000   58.320000   38.005000   58.320000 ;
      POLYGON   38.010000   85.745000   45.080000   78.675000   38.010000   78.675000 ;
      POLYGON   38.325000   92.500000   43.325000   92.500000   43.325000   87.500000 ;
      POLYGON   38.870000   70.745000   45.080000   70.745000   45.080000   64.535000 ;
      POLYGON   39.720000  -56.605000   45.935000  -56.605000   39.720000  -62.820000 ;
      POLYGON   40.585000  -69.030000   40.585000  -72.500000   37.115000  -72.500000 ;
      POLYGON   40.745000  -90.080000   40.745000  -92.500000   38.325000  -92.500000 ;
      POLYGON   42.465000  -95.435000   49.530000  -95.435000   42.465000 -102.500000 ;
      POLYGON   42.465000  102.500000   47.655000   97.310000   42.465000   97.310000 ;
      POLYGON   43.325000  -87.500000   43.325000  -90.080000   40.745000  -90.080000 ;
      POLYGON   43.325000  -73.360000   50.395000  -73.360000   43.325000  -80.430000 ;
      POLYGON   43.325000   87.500000   45.080000   87.500000   45.080000   85.745000 ;
      POLYGON   44.180000  -65.435000   44.180000  -69.030000   40.585000  -69.030000 ;
      POLYGON   44.220000   58.320000   51.285000   51.255000   44.220000   51.255000 ;
      POLYGON   44.540000  107.500000   48.690000  107.500000   48.690000  103.350000 ;
      POLYGON   45.080000   64.535000   51.295000   64.535000   51.295000   58.320000 ;
      POLYGON   45.080000   78.675000   52.150000   71.605000   45.080000   71.605000 ;
      POLYGON   45.080000   85.745000   52.150000   85.745000   52.150000   78.675000 ;
      POLYGON   45.935000  -50.395000   52.145000  -50.395000   45.935000  -56.605000 ;
      POLYGON   46.795000  -62.820000   46.795000  -65.435000   44.180000  -65.435000 ;
      POLYGON   46.800000 -105.240000   46.800000 -107.500000   44.540000 -107.500000 ;
      POLYGON   47.655000   97.310000   53.865000   91.100000   47.655000   91.100000 ;
      POLYGON   48.680000 -110.430000   55.750000 -110.430000   48.680000 -117.500000 ;
      POLYGON   48.680000  117.500000   54.730000  111.450000   48.680000  111.450000 ;
      POLYGON   48.690000  103.350000   49.540000  103.350000   49.540000  102.500000 ;
      POLYGON   49.530000  -88.360000   56.605000  -88.360000   49.530000  -95.435000 ;
      POLYGON   49.540000 -102.500000   49.540000 -105.240000   46.800000 -105.240000 ;
      POLYGON   49.540000  102.500000   54.730000  102.500000   54.730000   97.310000 ;
      POLYGON   50.075000  -38.325000   50.075000  -50.395000   38.005000  -50.395000 ;
      POLYGON   50.075000   38.325000   58.320000   38.325000   58.320000   30.080000 ;
      POLYGON   50.395000  -80.430000   50.395000  -87.500000   43.325000  -87.500000 ;
      POLYGON   50.395000  -66.290000   57.465000  -66.290000   50.395000  -73.360000 ;
      POLYGON   50.750000  122.500000   54.890000  122.500000   54.890000  118.360000 ;
      POLYGON   51.285000   51.255000   58.360000   44.180000   51.285000   44.180000 ;
      POLYGON   51.295000   58.320000   58.360000   58.320000   58.360000   51.255000 ;
      POLYGON   52.145000  -48.680000   53.860000  -48.680000   52.145000  -50.395000 ;
      POLYGON   52.145000  -36.255000   52.145000  -38.325000   50.075000  -38.325000 ;
      POLYGON   52.150000   71.605000   59.220000   64.535000   52.150000   64.535000 ;
      POLYGON   52.150000   78.675000   59.220000   78.675000   59.220000   71.605000 ;
      POLYGON   53.010000  -56.605000   53.010000  -62.820000   46.795000  -62.820000 ;
      POLYGON   53.860000  -42.465000   60.075000  -42.465000   53.860000  -48.680000 ;
      POLYGON   53.865000   91.100000   60.080000   84.885000   53.865000   84.885000 ;
      POLYGON   54.730000   97.310000   60.940000   97.310000   60.940000   91.100000 ;
      POLYGON   54.730000  111.450000   60.940000  105.240000   54.730000  105.240000 ;
      POLYGON   54.890000 -118.360000   54.890000 -122.500000   50.750000 -122.500000 ;
      POLYGON   54.890000 -118.360000   69.030000 -118.360000   54.890000 -132.500000 ;
      POLYGON   54.890000  118.360000   55.750000  118.360000   55.750000  117.500000 ;
      POLYGON   54.890000  132.500000   64.890000  122.500000   54.890000  122.500000 ;
      POLYGON   55.750000 -117.500000   55.750000 -118.360000   54.890000 -118.360000 ;
      POLYGON   55.750000 -103.360000   62.820000 -103.360000   55.750000 -110.430000 ;
      POLYGON   55.750000  117.500000   61.800000  117.500000   61.800000  111.450000 ;
      POLYGON   56.605000  -95.435000   56.605000 -102.500000   49.540000 -102.500000 ;
      POLYGON   56.605000  -81.295000   63.670000  -81.295000   56.605000  -88.360000 ;
      POLYGON   57.465000  -73.360000   57.465000  -80.430000   50.395000  -80.430000 ;
      POLYGON   57.465000  -61.800000   61.955000  -61.800000   57.465000  -66.290000 ;
      POLYGON   58.320000  -51.295000   58.320000  -56.605000   53.010000  -56.605000 ;
      POLYGON   58.320000   30.080000   58.360000   30.080000   58.360000   30.040000 ;
      POLYGON   58.360000   30.040000   62.500000   30.040000   62.500000   25.900000 ;
      POLYGON   58.360000   44.180000   65.425000   37.115000   58.360000   37.115000 ;
      POLYGON   58.360000   51.255000   65.435000   51.255000   65.435000   44.180000 ;
      POLYGON   59.220000  -50.395000   59.220000  -51.295000   58.320000  -51.295000 ;
      POLYGON   59.220000   64.535000   66.290000   57.465000   59.220000   57.465000 ;
      POLYGON   59.220000   71.605000   66.290000   71.605000   66.290000   64.535000 ;
      POLYGON   60.075000  -36.255000   66.285000  -36.255000   60.075000  -42.465000 ;
      POLYGON   60.080000   84.885000   67.145000   77.820000   60.080000   77.820000 ;
      POLYGON   60.935000  -48.680000   60.935000  -50.395000   59.220000  -50.395000 ;
      POLYGON   60.940000   91.100000   67.155000   91.100000   67.155000   84.885000 ;
      POLYGON   60.940000  105.240000   68.010000   98.170000   60.940000   98.170000 ;
      POLYGON   61.800000  111.450000   68.010000  111.450000   68.010000  105.240000 ;
      POLYGON   61.955000  -54.890000   68.865000  -54.890000   61.955000  -61.800000 ;
      POLYGON   62.500000  -25.900000   62.500000  -36.255000   52.145000  -36.255000 ;
      POLYGON   62.820000 -110.430000   62.820000 -117.500000   55.750000 -117.500000 ;
      POLYGON   62.820000  -96.290000   69.890000  -96.290000   62.820000 -103.360000 ;
      POLYGON   63.670000  -74.220000   70.745000  -74.220000   63.670000  -81.295000 ;
      POLYGON   63.680000  -88.360000   63.680000  -95.435000   56.605000  -95.435000 ;
      POLYGON   64.535000  -66.290000   64.535000  -73.360000   57.465000  -73.360000 ;
      POLYGON   64.890000  122.500000   75.940000  111.450000   64.890000  111.450000 ;
      POLYGON   65.425000   37.115000   72.500000   30.040000   65.425000   30.040000 ;
      POLYGON   65.435000   44.180000   72.500000   44.180000   72.500000   37.115000 ;
      POLYGON   66.285000  -30.040000   72.500000  -30.040000   66.285000  -36.255000 ;
      POLYGON   66.290000   57.465000   73.360000   50.395000   66.290000   50.395000 ;
      POLYGON   66.290000   64.535000   73.360000   64.535000   73.360000   57.465000 ;
      POLYGON   67.145000   77.820000   74.220000   70.745000   67.145000   70.745000 ;
      POLYGON   67.150000  -42.465000   67.150000  -48.680000   60.935000  -48.680000 ;
      POLYGON   67.155000   84.885000   74.220000   84.885000   74.220000   77.820000 ;
      POLYGON   68.010000   98.170000   75.080000   91.100000   68.010000   91.100000 ;
      POLYGON   68.010000  105.240000   75.080000  105.240000   75.080000   98.170000 ;
      POLYGON   68.865000  -48.680000   75.075000  -48.680000   68.865000  -54.890000 ;
      POLYGON   69.025000  -61.800000   69.025000  -66.290000   64.535000  -66.290000 ;
      POLYGON   69.030000 -104.220000   69.030000 -110.430000   62.820000 -110.430000 ;
      POLYGON   69.030000 -104.220000   83.170000 -104.220000   69.030000 -118.360000 ;
      POLYGON   69.890000 -103.360000   69.890000 -104.220000   69.030000 -104.220000 ;
      POLYGON   69.890000  -89.220000   76.960000  -89.220000   69.890000  -96.290000 ;
      POLYGON   70.745000  -81.295000   70.745000  -88.360000   63.680000  -88.360000 ;
      POLYGON   70.745000  -67.155000   77.810000  -67.155000   70.745000  -74.220000 ;
      POLYGON   72.500000   37.115000   77.500000   37.115000   77.500000   32.115000 ;
      POLYGON   73.360000  -36.255000   73.360000  -42.465000   67.150000  -42.465000 ;
      POLYGON   73.360000   50.395000   80.430000   43.325000   73.360000   43.325000 ;
      POLYGON   73.360000   57.465000   80.430000   57.465000   80.430000   50.395000 ;
      POLYGON   74.220000   70.745000   81.285000   63.680000   74.220000   63.680000 ;
      POLYGON   74.220000   77.820000   81.295000   77.820000   81.295000   70.745000 ;
      POLYGON   75.075000  -43.325000   80.430000  -43.325000   75.075000  -48.680000 ;
      POLYGON   75.080000   91.100000   82.150000   84.030000   75.080000   84.030000 ;
      POLYGON   75.080000   98.170000   75.940000   98.170000   75.940000   97.310000 ;
      POLYGON   75.935000  -54.890000   75.935000  -61.800000   69.025000  -61.800000 ;
      POLYGON   75.940000   97.310000   82.150000   97.310000   82.150000   91.100000 ;
      POLYGON   75.940000  111.450000   90.080000   97.310000   75.940000   97.310000 ;
      POLYGON   76.960000  -96.290000   76.960000 -103.360000   69.890000 -103.360000 ;
      POLYGON   76.960000  -82.150000   84.030000  -82.150000   76.960000  -89.220000 ;
      POLYGON   77.500000  -32.115000   77.500000  -36.255000   73.360000  -36.255000 ;
      POLYGON   77.810000  -61.800000   83.165000  -61.800000   77.810000  -67.155000 ;
      POLYGON   77.820000  -74.220000   77.820000  -81.295000   70.745000  -81.295000 ;
      POLYGON   78.675000  -52.150000   78.675000  -54.890000   75.935000  -54.890000 ;
      POLYGON   80.430000  -36.255000   87.500000  -36.255000   80.430000  -43.325000 ;
      POLYGON   80.430000   43.325000   87.500000   36.255000   80.430000   36.255000 ;
      POLYGON   80.430000   50.395000   87.500000   50.395000   87.500000   43.325000 ;
      POLYGON   81.285000   63.680000   88.360000   56.605000   81.285000   56.605000 ;
      POLYGON   81.295000   70.745000   88.360000   70.745000   88.360000   63.680000 ;
      POLYGON   82.145000  -48.680000   82.145000  -52.150000   78.675000  -52.150000 ;
      POLYGON   82.150000   84.030000   89.220000   76.960000   82.150000   76.960000 ;
      POLYGON   82.150000   91.100000   89.220000   91.100000   89.220000   84.030000 ;
      POLYGON   83.165000  -54.890000   90.075000  -54.890000   83.165000  -61.800000 ;
      POLYGON   83.170000  -90.080000   83.170000  -96.290000   76.960000  -96.290000 ;
      POLYGON   83.170000  -90.080000   97.310000  -90.080000   83.170000 -104.220000 ;
      POLYGON   84.030000  -89.220000   84.030000  -90.080000   83.170000  -90.080000 ;
      POLYGON   84.030000  -75.080000   91.100000  -75.080000   84.030000  -82.150000 ;
      POLYGON   84.885000  -67.155000   84.885000  -74.220000   77.820000  -74.220000 ;
      POLYGON   87.500000  -43.325000   87.500000  -48.680000   82.145000  -48.680000 ;
      POLYGON   87.500000   43.325000   92.500000   43.325000   92.500000   38.325000 ;
      POLYGON   88.360000   56.605000   95.425000   49.540000   88.360000   49.540000 ;
      POLYGON   88.360000   63.680000   95.435000   63.680000   95.435000   56.605000 ;
      POLYGON   89.220000   76.960000   96.290000   69.890000   89.220000   69.890000 ;
      POLYGON   89.220000   84.030000   90.080000   84.030000   90.080000   83.170000 ;
      POLYGON   90.075000  -48.680000   96.285000  -48.680000   90.075000  -54.890000 ;
      POLYGON   90.080000   83.170000   96.290000   83.170000   96.290000   76.960000 ;
      POLYGON   90.080000   97.310000  104.220000   83.170000   90.080000   83.170000 ;
      POLYGON   90.240000  -61.800000   90.240000  -67.155000   84.885000  -67.155000 ;
      POLYGON   91.100000  -82.150000   91.100000  -89.220000   84.030000  -89.220000 ;
      POLYGON   91.100000  -68.010000   98.170000  -68.010000   91.100000  -75.080000 ;
      POLYGON   92.500000  -38.325000   92.500000  -43.325000   87.500000  -43.325000 ;
      POLYGON   95.425000   49.540000  102.500000   42.465000   95.425000   42.465000 ;
      POLYGON   95.435000   56.605000  102.500000   56.605000  102.500000   49.540000 ;
      POLYGON   96.285000  -42.465000  102.500000  -42.465000   96.285000  -48.680000 ;
      POLYGON   96.290000   69.890000  103.360000   62.820000   96.290000   62.820000 ;
      POLYGON   96.290000   76.960000  103.360000   76.960000  103.360000   69.890000 ;
      POLYGON   97.150000  -54.890000   97.150000  -61.800000   90.240000  -61.800000 ;
      POLYGON   97.310000  -75.940000   97.310000  -82.150000   91.100000  -82.150000 ;
      POLYGON   97.310000  -75.940000  111.450000  -75.940000   97.310000  -90.080000 ;
      POLYGON   98.170000  -75.080000   98.170000  -75.940000   97.310000  -75.940000 ;
      POLYGON   98.170000  -61.800000  104.380000  -61.800000   98.170000  -68.010000 ;
      POLYGON  102.500000   49.540000  107.500000   49.540000  107.500000   44.540000 ;
      POLYGON  103.360000  -48.680000  103.360000  -54.890000   97.150000  -54.890000 ;
      POLYGON  103.360000   62.820000  110.430000   55.750000  103.360000   55.750000 ;
      POLYGON  103.360000   69.890000  104.220000   69.890000  104.220000   69.030000 ;
      POLYGON  104.220000   69.030000  110.430000   69.030000  110.430000   62.820000 ;
      POLYGON  104.220000   83.170000  118.360000   69.030000  104.220000   69.030000 ;
      POLYGON  104.380000  -55.750000  110.430000  -55.750000  104.380000  -61.800000 ;
      POLYGON  105.240000  -68.010000  105.240000  -75.080000   98.170000  -75.080000 ;
      POLYGON  107.500000  -44.540000  107.500000  -48.680000  103.360000  -48.680000 ;
      POLYGON  110.430000  -48.680000  117.500000  -48.680000  110.430000  -55.750000 ;
      POLYGON  110.430000   55.750000  117.500000   48.680000  110.430000   48.680000 ;
      POLYGON  110.430000   62.820000  117.500000   62.820000  117.500000   55.750000 ;
      POLYGON  111.450000  -61.800000  111.450000  -68.010000  105.240000  -68.010000 ;
      POLYGON  111.450000  -61.800000  125.590000  -61.800000  111.450000  -75.940000 ;
      POLYGON  117.500000  -55.750000  117.500000  -61.800000  111.450000  -61.800000 ;
      POLYGON  117.500000   55.750000  118.360000   55.750000  118.360000   54.890000 ;
      POLYGON  118.360000   54.890000  122.500000   54.890000  122.500000   50.750000 ;
      POLYGON  118.360000   69.030000  132.500000   54.890000  118.360000   54.890000 ;
      POLYGON  122.500000  -50.750000  122.500000  -55.750000  117.500000  -55.750000 ;
      POLYGON  125.590000  -54.890000  132.500000  -54.890000  125.590000  -61.800000 ;
      RECT -132.500000  -54.890000 -122.500000   54.890000 ;
      RECT -125.590000  -61.800000 -117.500000  -55.750000 ;
      RECT -125.590000  -55.750000 -122.500000  -54.890000 ;
      RECT -125.590000   54.890000 -118.360000   60.940000 ;
      RECT -125.590000   60.940000 -112.310000   61.800000 ;
      RECT -119.245000   61.800000 -112.310000   68.010000 ;
      RECT -119.245000   68.010000 -105.240000   68.145000 ;
      RECT -118.360000  -69.030000 -110.430000  -62.820000 ;
      RECT -118.360000  -62.820000 -117.500000  -61.800000 ;
      RECT -117.500000  -48.680000 -107.500000   45.940000 ;
      RECT -117.500000   45.940000 -106.100000   48.680000 ;
      RECT -115.430000  -50.750000 -102.500000  -49.540000 ;
      RECT -115.430000  -49.540000 -107.500000  -48.680000 ;
      RECT -115.430000   48.680000 -106.100000   50.750000 ;
      RECT -111.450000  -75.940000 -103.360000  -69.890000 ;
      RECT -111.450000  -69.890000 -110.430000  -69.030000 ;
      RECT -111.450000   68.145000 -105.240000   75.080000 ;
      RECT -111.450000   75.080000  -98.170000   75.940000 ;
      RECT -111.290000   50.750000 -106.100000   53.015000 ;
      RECT -111.290000   53.015000  -99.025000   54.890000 ;
      RECT -110.430000  -55.750000 -102.500000  -50.750000 ;
      RECT -105.240000   54.890000  -99.025000   60.080000 ;
      RECT -105.240000   60.080000  -91.960000   60.940000 ;
      RECT -104.245000   75.940000  -98.170000   82.150000 ;
      RECT -104.245000   82.150000  -91.100000   83.145000 ;
      RECT -104.220000  -83.170000  -96.290000  -76.960000 ;
      RECT -104.220000  -76.960000 -103.360000  -75.940000 ;
      RECT -103.360000  -62.820000  -95.435000  -56.605000 ;
      RECT -103.360000  -56.605000 -102.500000  -55.750000 ;
      RECT -102.500000  -42.465000  -92.500000   42.465000 ;
      RECT -100.425000  -44.540000  -87.500000  -43.325000 ;
      RECT -100.425000  -43.325000  -92.500000  -42.465000 ;
      RECT -100.425000   42.465000  -92.500000   44.540000 ;
      RECT  -99.025000   44.540000  -92.500000   45.080000 ;
      RECT  -99.025000   45.080000  -85.745000   45.940000 ;
      RECT  -98.170000   60.940000  -91.960000   67.155000 ;
      RECT  -98.170000   67.155000  -84.885000   68.010000 ;
      RECT  -97.310000  -90.080000  -89.220000  -84.030000 ;
      RECT  -97.310000  -84.030000  -96.290000  -83.170000 ;
      RECT  -97.310000   83.145000  -91.100000   89.220000 ;
      RECT  -97.310000   89.220000  -84.030000   90.080000 ;
      RECT  -96.290000  -69.890000  -88.360000  -63.680000 ;
      RECT  -96.290000  -63.680000  -95.435000  -62.820000 ;
      RECT  -95.425000  -49.540000  -87.500000  -44.540000 ;
      RECT  -91.950000   45.940000  -85.745000   52.150000 ;
      RECT  -91.950000   52.150000  -78.675000   53.015000 ;
      RECT  -91.100000   68.010000  -84.885000   74.220000 ;
      RECT  -91.100000   74.220000  -77.820000   75.080000 ;
      RECT  -90.535000   90.080000  -84.030000   94.235000 ;
      RECT  -90.535000   94.235000  -79.015000   96.855000 ;
      RECT  -89.250000  -98.140000  -82.150000  -91.100000 ;
      RECT  -89.250000  -91.100000  -89.220000  -90.080000 ;
      RECT  -89.220000  -76.960000  -81.295000  -70.745000 ;
      RECT  -89.220000  -70.745000  -88.360000  -69.890000 ;
      RECT  -88.360000  -56.605000  -80.430000  -50.395000 ;
      RECT  -88.360000  -50.395000  -87.500000  -49.540000 ;
      RECT  -87.500000  -36.255000  -77.500000   36.255000 ;
      RECT  -85.430000  -38.325000  -72.500000  -37.115000 ;
      RECT  -85.430000  -37.115000  -77.500000  -36.255000 ;
      RECT  -85.430000   36.255000  -77.500000   37.155000 ;
      RECT  -85.430000   37.155000  -72.460000   38.325000 ;
      RECT  -84.885000   53.015000  -78.675000   59.220000 ;
      RECT  -84.885000   59.220000  -71.605000   60.080000 ;
      RECT  -84.315000   75.080000  -77.820000   81.295000 ;
      RECT  -84.315000   81.295000  -70.745000   81.865000 ;
      RECT  -84.030000   81.865000  -70.745000   82.150000 ;
      RECT  -83.170000 -104.220000  -75.080000  -98.170000 ;
      RECT  -83.170000  -98.170000  -82.150000  -98.140000 ;
      RECT  -83.170000   96.855000  -79.015000   99.475000 ;
      RECT  -83.170000   99.475000  -73.775000  104.220000 ;
      RECT  -82.150000  -84.030000  -74.220000  -77.820000 ;
      RECT  -82.150000  -77.820000  -81.295000  -76.960000 ;
      RECT  -81.285000  -63.680000  -73.360000  -57.465000 ;
      RECT  -81.285000  -57.465000  -80.430000  -56.605000 ;
      RECT  -80.430000  -43.325000  -72.500000  -38.325000 ;
      RECT  -79.215000   38.325000  -72.460000   44.220000 ;
      RECT  -79.215000   44.220000  -65.395000   44.540000 ;
      RECT  -78.675000   44.540000  -65.395000   45.080000 ;
      RECT  -78.100000   60.080000  -71.605000   66.290000 ;
      RECT  -78.100000   66.290000  -64.535000   66.865000 ;
      RECT  -77.810000   66.865000  -64.535000   67.155000 ;
      RECT  -76.960000   82.150000  -70.745000   88.360000 ;
      RECT  -76.960000   88.360000  -63.680000   89.220000 ;
      RECT  -76.870000  104.220000  -73.775000  105.240000 ;
      RECT  -76.870000  105.240000  -68.010000  110.520000 ;
      RECT  -75.530000 -111.860000  -68.010000 -105.240000 ;
      RECT  -75.530000 -105.240000  -75.080000 -104.220000 ;
      RECT  -75.080000  -91.100000  -67.155000  -84.885000 ;
      RECT  -75.080000  -84.885000  -74.220000  -84.030000 ;
      RECT  -74.220000  -70.745000  -66.290000  -64.535000 ;
      RECT  -74.220000  -64.535000  -73.360000  -63.680000 ;
      RECT  -73.360000  -50.395000  -64.535000  -45.080000 ;
      RECT  -73.360000  -45.080000  -65.435000  -44.180000 ;
      RECT  -73.360000  -44.180000  -72.500000  -43.325000 ;
      RECT  -72.500000  -30.040000  -62.500000   -5.000000 ;
      RECT  -72.500000   -5.000000   57.500000    5.000000 ;
      RECT  -72.500000    5.000000  -62.500000   30.040000 ;
      RECT  -72.460000   30.040000  -62.500000   30.080000 ;
      RECT  -71.945000   89.220000  -63.680000   94.235000 ;
      RECT  -71.605000   45.080000  -65.395000   51.295000 ;
      RECT  -71.605000   51.295000  -58.320000   52.150000 ;
      RECT  -70.745000   67.155000  -64.535000   73.360000 ;
      RECT  -70.745000   73.360000  -57.465000   74.220000 ;
      RECT  -70.665000   94.235000  -57.805000   95.515000 ;
      RECT  -70.425000  -32.115000  -62.500000  -30.040000 ;
      RECT  -70.425000   30.080000  -58.320000   32.115000 ;
      RECT  -69.030000 -118.360000  -60.940000 -112.310000 ;
      RECT  -69.030000 -112.310000  -68.010000 -111.860000 ;
      RECT  -69.030000  110.520000  -68.010000  111.450000 ;
      RECT  -69.030000  111.450000  -61.800000  118.360000 ;
      RECT  -68.010000  -98.170000  -60.080000  -91.960000 ;
      RECT  -68.010000  -91.960000  -67.155000  -91.100000 ;
      RECT  -67.145000  -77.820000  -59.220000  -71.605000 ;
      RECT  -67.145000  -71.605000  -66.290000  -70.745000 ;
      RECT  -66.705000   95.515000  -57.805000   99.475000 ;
      RECT  -66.290000  -57.465000  -58.360000  -51.255000 ;
      RECT  -66.290000  -51.255000  -64.535000  -50.395000 ;
      RECT  -65.425000  -37.115000  -62.500000  -32.115000 ;
      RECT  -65.385000   32.115000  -58.320000   37.155000 ;
      RECT  -64.535000   52.150000  -58.320000   58.320000 ;
      RECT  -64.535000   58.320000  -51.295000   59.220000 ;
      RECT  -64.440000   74.220000  -57.465000   79.245000 ;
      RECT  -64.440000   79.245000  -51.580000   80.525000 ;
      RECT  -64.215000  -38.325000  -62.500000  -37.115000 ;
      RECT  -63.670000   80.525000  -51.580000   81.295000 ;
      RECT  -62.820000   99.475000  -57.805000  100.755000 ;
      RECT  -62.820000  100.755000  -51.285000  103.360000 ;
      RECT  -60.940000 -105.240000  -53.015000  -99.025000 ;
      RECT  -60.940000  -99.025000  -60.080000  -98.170000 ;
      RECT  -60.940000  103.360000  -51.285000  105.240000 ;
      RECT  -60.080000  -84.885000  -52.150000  -78.675000 ;
      RECT  -60.080000  -78.675000  -59.220000  -77.820000 ;
      RECT  -59.220000  -64.535000  -51.295000  -58.320000 ;
      RECT  -59.220000  -58.320000  -58.360000  -57.465000 ;
      RECT  -58.360000  -44.180000  -50.075000  -38.325000 ;
      RECT  -58.320000   38.325000  -50.075000   44.220000 ;
      RECT  -58.230000   59.220000  -51.295000   64.245000 ;
      RECT  -58.230000   64.245000  -45.370000   65.525000 ;
      RECT  -57.465000   65.525000  -45.370000   66.290000 ;
      RECT  -57.460000  -45.080000  -50.075000  -44.180000 ;
      RECT  -56.940000  105.240000  -51.285000  107.500000 ;
      RECT  -56.940000  107.500000  -11.010000  108.735000 ;
      RECT  -56.940000  108.735000   -9.775000  109.240000 ;
      RECT  -56.605000   81.295000  -51.580000   85.765000 ;
      RECT  -56.605000   85.765000  -45.060000   88.360000 ;
      RECT  -54.890000 -132.500000  -11.010000 -131.265000 ;
      RECT  -54.890000 -131.265000   -9.775000 -123.735000 ;
      RECT  -54.890000 -123.735000  -11.010000 -122.500000 ;
      RECT  -54.890000  122.500000   54.890000  132.500000 ;
      RECT  -54.730000  109.240000   -9.775000  111.450000 ;
      RECT  -53.870000 -112.310000   -5.425000 -107.500000 ;
      RECT  -53.870000 -107.500000  -46.800000 -105.240000 ;
      RECT  -53.005000  -91.960000  -45.080000  -85.745000 ;
      RECT  -53.005000  -85.745000  -52.150000  -84.885000 ;
      RECT  -52.150000  -71.605000  -38.870000  -70.745000 ;
      RECT  -52.150000  -70.745000  -44.220000  -65.395000 ;
      RECT  -52.150000  -65.395000  -51.295000  -64.535000 ;
      RECT  -51.285000  -51.255000  -37.650000  -50.750000 ;
      RECT  -51.285000  -50.750000  -50.075000  -45.080000 ;
      RECT  -51.245000   44.220000  -50.075000   50.395000 ;
      RECT  -51.245000   50.395000  -38.005000   51.295000 ;
      RECT  -50.730000   88.360000  -45.060000   92.500000 ;
      RECT  -50.730000   92.500000   -5.425000   94.235000 ;
      RECT  -50.395000   66.290000  -45.370000   70.745000 ;
      RECT  -50.395000   70.745000  -38.870000   73.360000 ;
      RECT  -48.680000 -117.500000   -5.425000 -112.310000 ;
      RECT  -48.680000  111.450000   -9.775000  116.265000 ;
      RECT  -48.680000  116.265000  -11.010000  117.500000 ;
      RECT  -45.940000  -99.025000   -9.775000  -93.735000 ;
      RECT  -45.940000  -93.735000  -11.010000  -92.500000 ;
      RECT  -45.940000  -92.500000  -45.080000  -91.960000 ;
      RECT  -45.080000  -78.675000   -5.425000  -77.500000 ;
      RECT  -45.080000  -77.500000  -38.870000  -71.605000 ;
      RECT  -44.510000   73.360000  -38.870000   77.500000 ;
      RECT  -44.510000   77.500000  -11.010000   78.735000 ;
      RECT  -44.510000   78.735000   -9.775000   79.245000 ;
      RECT  -44.220000  -58.320000  -37.650000  -51.255000 ;
      RECT  -44.220000   51.295000  -38.005000   58.320000 ;
      RECT  -44.210000   94.235000   -5.425000  100.755000 ;
      RECT  -42.465000 -102.500000  -11.010000 -101.265000 ;
      RECT  -42.465000 -101.265000   -9.775000  -99.025000 ;
      RECT  -42.465000  100.755000   -5.425000  102.500000 ;
      RECT  -38.295000   58.320000  -38.005000   62.500000 ;
      RECT  -38.295000   62.500000   -5.425000   64.245000 ;
      RECT  -38.010000  -85.745000   -5.425000  -78.675000 ;
      RECT  -38.005000  -64.535000   33.510000  -62.820000 ;
      RECT  -38.005000  -62.820000   39.720000  -62.500000 ;
      RECT  -38.005000  -62.500000  -37.650000  -58.320000 ;
      RECT  -37.990000   79.245000   -9.775000   85.765000 ;
      RECT  -37.145000  -65.395000   33.510000  -64.535000 ;
      RECT  -36.255000  -87.500000   -5.425000  -85.745000 ;
      RECT  -36.255000   85.765000   -9.775000   86.265000 ;
      RECT  -36.255000   86.265000  -11.010000   87.500000 ;
      RECT  -31.795000  -70.745000   30.040000  -69.030000 ;
      RECT  -31.795000  -69.030000   33.510000  -65.395000 ;
      RECT  -31.795000   64.245000   -5.425000   70.745000 ;
      RECT  -30.040000  -72.500000   30.040000  -70.745000 ;
      RECT  -30.040000   70.745000   -5.425000   72.500000 ;
      RECT   -8.725000   72.500000   -5.425000   73.350000 ;
      RECT   -8.725000  102.500000   -5.425000  103.350000 ;
      RECT   -8.715000 -118.360000   -5.425000 -117.500000 ;
      RECT   -5.975000  -91.100000    7.155000  -90.080000 ;
      RECT   -5.975000  -90.080000   -5.425000  -87.500000 ;
      RECT   -4.575000 -122.500000    5.435000 -118.360000 ;
      RECT   -4.575000  -92.500000    7.155000  -91.100000 ;
      RECT   -4.575000   73.350000    5.425000   77.500000 ;
      RECT   -4.575000  103.350000    5.425000  107.500000 ;
      RECT    5.425000 -132.500000   54.890000 -122.500000 ;
      RECT    5.425000 -102.500000   42.465000  -95.435000 ;
      RECT    5.425000  -95.435000   49.530000  -92.500000 ;
      RECT    5.425000   77.500000   45.080000   78.675000 ;
      RECT    5.425000   78.675000   38.010000   85.745000 ;
      RECT    5.425000   85.745000   36.255000   87.500000 ;
      RECT    5.425000  107.500000   54.730000  111.450000 ;
      RECT    5.425000  111.450000   48.680000  117.500000 ;
      RECT    8.660000 -116.265000   48.680000 -110.430000 ;
      RECT    8.660000 -110.430000   55.750000 -108.735000 ;
      RECT    8.660000  -86.265000   36.255000  -80.430000 ;
      RECT    8.660000  -80.430000   43.325000  -78.735000 ;
      RECT    8.660000   63.735000   38.005000   64.535000 ;
      RECT    8.660000   64.535000   31.795000   70.745000 ;
      RECT    8.660000   70.745000   30.040000   71.265000 ;
      RECT    8.660000   93.735000   47.655000   97.310000 ;
      RECT    8.660000   97.310000   42.465000  101.265000 ;
      RECT    9.895000 -117.500000   48.680000 -116.265000 ;
      RECT    9.895000 -108.735000   55.750000 -107.500000 ;
      RECT    9.895000  -87.500000   36.255000  -86.265000 ;
      RECT    9.895000  -78.735000   43.325000  -77.500000 ;
      RECT    9.895000   62.500000   38.005000   63.735000 ;
      RECT    9.895000   71.265000   30.040000   72.500000 ;
      RECT    9.895000   92.500000   47.655000   93.735000 ;
      RECT    9.895000  101.265000   42.465000  102.500000 ;
      RECT   33.675000  -77.500000   43.325000  -75.940000 ;
      RECT   36.265000   73.350000   45.080000   77.500000 ;
      RECT   37.115000  -75.940000   43.325000  -73.360000 ;
      RECT   37.115000  -73.360000   50.395000  -72.500000 ;
      RECT   37.115000   72.500000   45.080000   73.350000 ;
      RECT   37.650000  -62.500000   39.720000  -56.605000 ;
      RECT   37.650000  -56.605000   45.935000  -50.750000 ;
      RECT   38.005000  -50.750000   45.935000  -50.395000 ;
      RECT   38.005000   50.395000   51.285000   51.255000 ;
      RECT   38.005000   51.255000   44.220000   58.320000 ;
      RECT   38.870000   70.745000   52.150000   71.605000 ;
      RECT   38.870000   71.605000   45.080000   72.500000 ;
      RECT   40.585000  -72.500000   50.395000  -69.030000 ;
      RECT   40.745000  -92.500000   49.530000  -90.080000 ;
      RECT   43.325000  -90.080000   49.530000  -88.360000 ;
      RECT   43.325000  -88.360000   56.605000  -87.500000 ;
      RECT   43.325000   87.500000   53.865000   91.100000 ;
      RECT   43.325000   91.100000   47.655000   92.500000 ;
      RECT   44.180000  -69.030000   50.395000  -66.290000 ;
      RECT   44.180000  -66.290000   57.465000  -65.435000 ;
      RECT   45.080000   64.535000   52.150000   70.745000 ;
      RECT   45.080000   85.745000   53.865000   87.500000 ;
      RECT   46.795000  -65.435000   57.465000  -62.820000 ;
      RECT   46.800000 -107.500000   55.750000 -105.240000 ;
      RECT   48.690000  103.350000   60.940000  105.240000 ;
      RECT   48.690000  105.240000   54.730000  107.500000 ;
      RECT   49.540000 -105.240000   55.750000 -103.360000 ;
      RECT   49.540000 -103.360000   62.820000 -102.500000 ;
      RECT   49.540000  102.500000   60.940000  103.350000 ;
      RECT   50.075000  -50.395000   52.145000  -48.680000 ;
      RECT   50.075000  -48.680000   53.860000  -42.465000 ;
      RECT   50.075000  -42.465000   60.075000  -38.325000 ;
      RECT   50.075000   38.325000   58.360000   44.180000 ;
      RECT   50.075000   44.180000   51.285000   50.395000 ;
      RECT   50.395000  -87.500000   56.605000  -81.295000 ;
      RECT   50.395000  -81.295000   63.670000  -80.430000 ;
      RECT   51.295000   58.320000   59.220000   64.535000 ;
      RECT   52.145000  -38.325000   60.075000  -36.255000 ;
      RECT   52.150000   78.675000   60.080000   84.885000 ;
      RECT   52.150000   84.885000   53.865000   85.745000 ;
      RECT   53.010000  -62.820000   57.465000  -61.800000 ;
      RECT   53.010000  -61.800000   61.955000  -56.605000 ;
      RECT   54.730000   97.310000   68.010000   98.170000 ;
      RECT   54.730000   98.170000   60.940000  102.500000 ;
      RECT   54.890000  118.360000   64.890000  122.500000 ;
      RECT   55.750000 -118.360000   69.030000 -117.500000 ;
      RECT   55.750000  117.500000   64.890000  118.360000 ;
      RECT   56.605000 -102.500000   62.820000  -96.290000 ;
      RECT   56.605000  -96.290000   69.890000  -95.435000 ;
      RECT   57.465000  -80.430000   63.670000  -74.220000 ;
      RECT   57.465000  -74.220000   70.745000  -73.360000 ;
      RECT   58.320000  -56.605000   61.955000  -54.890000 ;
      RECT   58.320000  -54.890000   68.865000  -51.295000 ;
      RECT   58.320000   30.080000   65.425000   37.115000 ;
      RECT   58.320000   37.115000   58.360000   38.325000 ;
      RECT   58.360000   30.040000   65.425000   30.080000 ;
      RECT   58.360000   51.255000   66.290000   57.465000 ;
      RECT   58.360000   57.465000   59.220000   58.320000 ;
      RECT   59.220000  -51.295000   68.865000  -50.395000 ;
      RECT   59.220000   71.605000   67.145000   77.820000 ;
      RECT   59.220000   77.820000   60.080000   78.675000 ;
      RECT   60.935000  -50.395000   68.865000  -48.680000 ;
      RECT   60.940000   91.100000   68.010000   97.310000 ;
      RECT   61.800000  111.450000   64.890000  117.500000 ;
      RECT   62.500000  -36.255000   66.285000  -30.040000 ;
      RECT   62.500000  -30.040000   72.500000   30.040000 ;
      RECT   62.820000 -117.500000   69.030000 -110.430000 ;
      RECT   63.680000  -95.435000   69.890000  -89.220000 ;
      RECT   63.680000  -89.220000   76.960000  -88.360000 ;
      RECT   64.535000  -73.360000   70.745000  -67.155000 ;
      RECT   64.535000  -67.155000   77.810000  -66.290000 ;
      RECT   65.435000   44.180000   73.360000   50.395000 ;
      RECT   65.435000   50.395000   66.290000   51.255000 ;
      RECT   66.290000   64.535000   74.220000   70.745000 ;
      RECT   66.290000   70.745000   67.145000   71.605000 ;
      RECT   67.150000  -48.680000   75.075000  -43.325000 ;
      RECT   67.150000  -43.325000   80.430000  -42.465000 ;
      RECT   67.155000   84.885000   75.080000   91.100000 ;
      RECT   68.010000  105.240000   75.940000  111.450000 ;
      RECT   69.025000  -66.290000   77.810000  -61.800000 ;
      RECT   69.890000 -104.220000   83.170000 -103.360000 ;
      RECT   70.745000  -88.360000   76.960000  -82.150000 ;
      RECT   70.745000  -82.150000   84.030000  -81.295000 ;
      RECT   72.500000   37.115000   80.430000   43.325000 ;
      RECT   72.500000   43.325000   73.360000   44.180000 ;
      RECT   73.360000  -42.465000   80.430000  -36.255000 ;
      RECT   73.360000   57.465000   81.285000   63.680000 ;
      RECT   73.360000   63.680000   74.220000   64.535000 ;
      RECT   74.220000   77.820000   82.150000   84.030000 ;
      RECT   74.220000   84.030000   75.080000   84.885000 ;
      RECT   75.080000   98.170000   75.940000  105.240000 ;
      RECT   75.935000  -61.800000   83.165000  -54.890000 ;
      RECT   76.960000 -103.360000   83.170000  -96.290000 ;
      RECT   77.500000  -36.255000   87.500000   36.255000 ;
      RECT   77.500000   36.255000   80.430000   37.115000 ;
      RECT   77.820000  -81.295000   84.030000  -75.080000 ;
      RECT   77.820000  -75.080000   91.100000  -74.220000 ;
      RECT   78.675000  -54.890000   90.075000  -52.150000 ;
      RECT   80.430000   50.395000   88.360000   56.605000 ;
      RECT   80.430000   56.605000   81.285000   57.465000 ;
      RECT   81.295000   70.745000   89.220000   76.960000 ;
      RECT   81.295000   76.960000   82.150000   77.820000 ;
      RECT   82.145000  -52.150000   90.075000  -48.680000 ;
      RECT   82.150000   91.100000   90.080000   97.310000 ;
      RECT   84.030000  -90.080000   97.310000  -89.220000 ;
      RECT   84.885000  -74.220000   91.100000  -68.010000 ;
      RECT   84.885000  -68.010000   98.170000  -67.155000 ;
      RECT   87.500000  -48.680000   96.285000  -43.325000 ;
      RECT   87.500000   43.325000   95.425000   49.540000 ;
      RECT   87.500000   49.540000   88.360000   50.395000 ;
      RECT   88.360000   63.680000   96.290000   69.890000 ;
      RECT   88.360000   69.890000   89.220000   70.745000 ;
      RECT   89.220000   84.030000   90.080000   91.100000 ;
      RECT   90.240000  -67.155000   98.170000  -61.800000 ;
      RECT   91.100000  -89.220000   97.310000  -82.150000 ;
      RECT   92.500000  -43.325000   96.285000  -42.465000 ;
      RECT   92.500000  -42.465000  102.500000   42.465000 ;
      RECT   92.500000   42.465000   95.425000   43.325000 ;
      RECT   95.435000   56.605000  103.360000   62.820000 ;
      RECT   95.435000   62.820000   96.290000   63.680000 ;
      RECT   96.290000   76.960000  104.220000   83.170000 ;
      RECT   97.150000  -61.800000  104.380000  -55.750000 ;
      RECT   97.150000  -55.750000  110.430000  -54.890000 ;
      RECT   98.170000  -75.940000  111.450000  -75.080000 ;
      RECT  102.500000   49.540000  110.430000   55.750000 ;
      RECT  102.500000   55.750000  103.360000   56.605000 ;
      RECT  103.360000  -54.890000  110.430000  -48.680000 ;
      RECT  103.360000   69.890000  104.220000   76.960000 ;
      RECT  105.240000  -75.080000  111.450000  -68.010000 ;
      RECT  107.500000  -48.680000  117.500000   48.680000 ;
      RECT  107.500000   48.680000  110.430000   49.540000 ;
      RECT  110.430000   62.820000  118.360000   69.030000 ;
      RECT  117.500000  -61.800000  125.590000  -55.750000 ;
      RECT  117.500000   55.750000  118.360000   62.820000 ;
      RECT  122.500000  -55.750000  125.590000  -54.890000 ;
      RECT  122.500000  -54.890000  132.500000  -25.000000 ;
      RECT  122.500000  -25.000000  137.500000  -15.000000 ;
      RECT  122.500000   15.000000  137.500000   25.000000 ;
      RECT  122.500000   25.000000  132.500000   54.890000 ;
    LAYER via2 ;
      RECT -30.655000   79.245000 -29.375000   80.525000 ;
      RECT -30.655000   81.865000 -29.375000   83.145000 ;
      RECT -30.655000   84.485000 -29.375000   85.765000 ;
      RECT -30.650000 -130.760000 -29.370000 -129.480000 ;
      RECT -30.650000 -128.140000 -29.370000 -126.860000 ;
      RECT -30.650000 -125.520000 -29.370000 -124.240000 ;
      RECT -30.650000 -100.760000 -29.370000  -99.480000 ;
      RECT -30.650000  -98.140000 -29.370000  -96.860000 ;
      RECT -30.650000  -95.520000 -29.370000  -94.240000 ;
      RECT -30.650000  109.240000 -29.370000  110.520000 ;
      RECT -30.650000  111.860000 -29.370000  113.140000 ;
      RECT -30.650000  114.480000 -29.370000  115.760000 ;
      RECT -28.035000   79.245000 -26.755000   80.525000 ;
      RECT -28.035000   81.865000 -26.755000   83.145000 ;
      RECT -28.035000   84.485000 -26.755000   85.765000 ;
      RECT -28.030000 -130.760000 -26.750000 -129.480000 ;
      RECT -28.030000 -128.140000 -26.750000 -126.860000 ;
      RECT -28.030000 -125.520000 -26.750000 -124.240000 ;
      RECT -28.030000 -100.760000 -26.750000  -99.480000 ;
      RECT -28.030000  -98.140000 -26.750000  -96.860000 ;
      RECT -28.030000  -95.520000 -26.750000  -94.240000 ;
      RECT -28.030000  109.240000 -26.750000  110.520000 ;
      RECT -28.030000  111.860000 -26.750000  113.140000 ;
      RECT -28.030000  114.480000 -26.750000  115.760000 ;
      RECT -25.265000   79.245000 -23.985000   80.525000 ;
      RECT -25.265000   81.865000 -23.985000   83.145000 ;
      RECT -25.265000   84.485000 -23.985000   85.765000 ;
      RECT -25.260000 -130.760000 -23.980000 -129.480000 ;
      RECT -25.260000 -128.140000 -23.980000 -126.860000 ;
      RECT -25.260000 -125.520000 -23.980000 -124.240000 ;
      RECT -25.260000 -100.760000 -23.980000  -99.480000 ;
      RECT -25.260000  -98.140000 -23.980000  -96.860000 ;
      RECT -25.260000  -95.520000 -23.980000  -94.240000 ;
      RECT -25.260000  109.240000 -23.980000  110.520000 ;
      RECT -25.260000  111.860000 -23.980000  113.140000 ;
      RECT -25.260000  114.480000 -23.980000  115.760000 ;
      RECT -22.495000   79.245000 -21.215000   80.525000 ;
      RECT -22.495000   81.865000 -21.215000   83.145000 ;
      RECT -22.495000   84.485000 -21.215000   85.765000 ;
      RECT -22.490000 -130.760000 -21.210000 -129.480000 ;
      RECT -22.490000 -128.140000 -21.210000 -126.860000 ;
      RECT -22.490000 -125.520000 -21.210000 -124.240000 ;
      RECT -22.490000 -100.760000 -21.210000  -99.480000 ;
      RECT -22.490000  -98.140000 -21.210000  -96.860000 ;
      RECT -22.490000  -95.520000 -21.210000  -94.240000 ;
      RECT -22.490000  109.240000 -21.210000  110.520000 ;
      RECT -22.490000  111.860000 -21.210000  113.140000 ;
      RECT -22.490000  114.480000 -21.210000  115.760000 ;
      RECT -19.725000   79.245000 -18.445000   80.525000 ;
      RECT -19.725000   81.865000 -18.445000   83.145000 ;
      RECT -19.725000   84.485000 -18.445000   85.765000 ;
      RECT -19.720000 -130.760000 -18.440000 -129.480000 ;
      RECT -19.720000 -128.140000 -18.440000 -126.860000 ;
      RECT -19.720000 -125.520000 -18.440000 -124.240000 ;
      RECT -19.720000 -100.760000 -18.440000  -99.480000 ;
      RECT -19.720000  -98.140000 -18.440000  -96.860000 ;
      RECT -19.720000  -95.520000 -18.440000  -94.240000 ;
      RECT -19.720000  109.240000 -18.440000  110.520000 ;
      RECT -19.720000  111.860000 -18.440000  113.140000 ;
      RECT -19.720000  114.480000 -18.440000  115.760000 ;
      RECT -16.955000   79.245000 -15.675000   80.525000 ;
      RECT -16.955000   81.865000 -15.675000   83.145000 ;
      RECT -16.955000   84.485000 -15.675000   85.765000 ;
      RECT -16.950000 -130.760000 -15.670000 -129.480000 ;
      RECT -16.950000 -128.140000 -15.670000 -126.860000 ;
      RECT -16.950000 -125.520000 -15.670000 -124.240000 ;
      RECT -16.950000 -100.760000 -15.670000  -99.480000 ;
      RECT -16.950000  -98.140000 -15.670000  -96.860000 ;
      RECT -16.950000  -95.520000 -15.670000  -94.240000 ;
      RECT -16.950000  109.240000 -15.670000  110.520000 ;
      RECT -16.950000  111.860000 -15.670000  113.140000 ;
      RECT -16.950000  114.480000 -15.670000  115.760000 ;
      RECT -14.185000   79.245000 -12.905000   80.525000 ;
      RECT -14.185000   81.865000 -12.905000   83.145000 ;
      RECT -14.185000   84.485000 -12.905000   85.765000 ;
      RECT -14.180000 -130.760000 -12.900000 -129.480000 ;
      RECT -14.180000 -128.140000 -12.900000 -126.860000 ;
      RECT -14.180000 -125.520000 -12.900000 -124.240000 ;
      RECT -14.180000 -100.760000 -12.900000  -99.480000 ;
      RECT -14.180000  -98.140000 -12.900000  -96.860000 ;
      RECT -14.180000  -95.520000 -12.900000  -94.240000 ;
      RECT -14.180000  109.240000 -12.900000  110.520000 ;
      RECT -14.180000  111.860000 -12.900000  113.140000 ;
      RECT -14.180000  114.480000 -12.900000  115.760000 ;
      RECT -11.565000   79.245000 -10.285000   80.525000 ;
      RECT -11.565000   81.865000 -10.285000   83.145000 ;
      RECT -11.565000   84.485000 -10.285000   85.765000 ;
      RECT -11.560000 -130.760000 -10.280000 -129.480000 ;
      RECT -11.560000 -128.140000 -10.280000 -126.860000 ;
      RECT -11.560000 -125.520000 -10.280000 -124.240000 ;
      RECT -11.560000 -100.760000 -10.280000  -99.480000 ;
      RECT -11.560000  -98.140000 -10.280000  -96.860000 ;
      RECT -11.560000  -95.520000 -10.280000  -94.240000 ;
      RECT -11.560000  109.240000 -10.280000  110.520000 ;
      RECT -11.560000  111.860000 -10.280000  113.140000 ;
      RECT -11.560000  114.480000 -10.280000  115.760000 ;
      RECT   9.160000  -85.765000  10.440000  -84.485000 ;
      RECT   9.160000  -83.145000  10.440000  -81.865000 ;
      RECT   9.160000  -80.525000  10.440000  -79.245000 ;
      RECT   9.165000 -115.760000  10.445000 -114.480000 ;
      RECT   9.165000 -113.140000  10.445000 -111.860000 ;
      RECT   9.165000 -110.520000  10.445000 -109.240000 ;
      RECT   9.165000   64.245000  10.445000   65.525000 ;
      RECT   9.165000   66.865000  10.445000   68.145000 ;
      RECT   9.165000   69.485000  10.445000   70.765000 ;
      RECT   9.165000   94.235000  10.445000   95.515000 ;
      RECT   9.165000   96.855000  10.445000   98.135000 ;
      RECT   9.165000   99.475000  10.445000  100.755000 ;
      RECT  11.780000  -85.765000  13.060000  -84.485000 ;
      RECT  11.780000  -83.145000  13.060000  -81.865000 ;
      RECT  11.780000  -80.525000  13.060000  -79.245000 ;
      RECT  11.785000 -115.760000  13.065000 -114.480000 ;
      RECT  11.785000 -113.140000  13.065000 -111.860000 ;
      RECT  11.785000 -110.520000  13.065000 -109.240000 ;
      RECT  11.785000   64.245000  13.065000   65.525000 ;
      RECT  11.785000   66.865000  13.065000   68.145000 ;
      RECT  11.785000   69.485000  13.065000   70.765000 ;
      RECT  11.785000   94.235000  13.065000   95.515000 ;
      RECT  11.785000   96.855000  13.065000   98.135000 ;
      RECT  11.785000   99.475000  13.065000  100.755000 ;
      RECT  14.550000  -85.765000  15.830000  -84.485000 ;
      RECT  14.550000  -83.145000  15.830000  -81.865000 ;
      RECT  14.550000  -80.525000  15.830000  -79.245000 ;
      RECT  14.555000 -115.760000  15.835000 -114.480000 ;
      RECT  14.555000 -113.140000  15.835000 -111.860000 ;
      RECT  14.555000 -110.520000  15.835000 -109.240000 ;
      RECT  14.555000   64.245000  15.835000   65.525000 ;
      RECT  14.555000   66.865000  15.835000   68.145000 ;
      RECT  14.555000   69.485000  15.835000   70.765000 ;
      RECT  14.555000   94.235000  15.835000   95.515000 ;
      RECT  14.555000   96.855000  15.835000   98.135000 ;
      RECT  14.555000   99.475000  15.835000  100.755000 ;
      RECT  17.320000  -85.765000  18.600000  -84.485000 ;
      RECT  17.320000  -83.145000  18.600000  -81.865000 ;
      RECT  17.320000  -80.525000  18.600000  -79.245000 ;
      RECT  17.325000 -115.760000  18.605000 -114.480000 ;
      RECT  17.325000 -113.140000  18.605000 -111.860000 ;
      RECT  17.325000 -110.520000  18.605000 -109.240000 ;
      RECT  17.325000   64.245000  18.605000   65.525000 ;
      RECT  17.325000   66.865000  18.605000   68.145000 ;
      RECT  17.325000   69.485000  18.605000   70.765000 ;
      RECT  17.325000   94.235000  18.605000   95.515000 ;
      RECT  17.325000   96.855000  18.605000   98.135000 ;
      RECT  17.325000   99.475000  18.605000  100.755000 ;
      RECT  20.090000  -85.765000  21.370000  -84.485000 ;
      RECT  20.090000  -83.145000  21.370000  -81.865000 ;
      RECT  20.090000  -80.525000  21.370000  -79.245000 ;
      RECT  20.095000 -115.760000  21.375000 -114.480000 ;
      RECT  20.095000 -113.140000  21.375000 -111.860000 ;
      RECT  20.095000 -110.520000  21.375000 -109.240000 ;
      RECT  20.095000   64.245000  21.375000   65.525000 ;
      RECT  20.095000   66.865000  21.375000   68.145000 ;
      RECT  20.095000   69.485000  21.375000   70.765000 ;
      RECT  20.095000   94.235000  21.375000   95.515000 ;
      RECT  20.095000   96.855000  21.375000   98.135000 ;
      RECT  20.095000   99.475000  21.375000  100.755000 ;
      RECT  22.860000  -85.765000  24.140000  -84.485000 ;
      RECT  22.860000  -83.145000  24.140000  -81.865000 ;
      RECT  22.860000  -80.525000  24.140000  -79.245000 ;
      RECT  22.865000 -115.760000  24.145000 -114.480000 ;
      RECT  22.865000 -113.140000  24.145000 -111.860000 ;
      RECT  22.865000 -110.520000  24.145000 -109.240000 ;
      RECT  22.865000   64.245000  24.145000   65.525000 ;
      RECT  22.865000   66.865000  24.145000   68.145000 ;
      RECT  22.865000   69.485000  24.145000   70.765000 ;
      RECT  22.865000   94.235000  24.145000   95.515000 ;
      RECT  22.865000   96.855000  24.145000   98.135000 ;
      RECT  22.865000   99.475000  24.145000  100.755000 ;
      RECT  25.630000  -85.765000  26.910000  -84.485000 ;
      RECT  25.630000  -83.145000  26.910000  -81.865000 ;
      RECT  25.630000  -80.525000  26.910000  -79.245000 ;
      RECT  25.635000 -115.760000  26.915000 -114.480000 ;
      RECT  25.635000 -113.140000  26.915000 -111.860000 ;
      RECT  25.635000 -110.520000  26.915000 -109.240000 ;
      RECT  25.635000   64.245000  26.915000   65.525000 ;
      RECT  25.635000   66.865000  26.915000   68.145000 ;
      RECT  25.635000   69.485000  26.915000   70.765000 ;
      RECT  25.635000   94.235000  26.915000   95.515000 ;
      RECT  25.635000   96.855000  26.915000   98.135000 ;
      RECT  25.635000   99.475000  26.915000  100.755000 ;
      RECT  28.250000  -85.765000  29.530000  -84.485000 ;
      RECT  28.250000  -83.145000  29.530000  -81.865000 ;
      RECT  28.250000  -80.525000  29.530000  -79.245000 ;
      RECT  28.255000 -115.760000  29.535000 -114.480000 ;
      RECT  28.255000 -113.140000  29.535000 -111.860000 ;
      RECT  28.255000 -110.520000  29.535000 -109.240000 ;
      RECT  28.255000   64.245000  29.535000   65.525000 ;
      RECT  28.255000   66.865000  29.535000   68.145000 ;
      RECT  28.255000   69.485000  29.535000   70.765000 ;
      RECT  28.255000   94.235000  29.535000   95.515000 ;
      RECT  28.255000   96.855000  29.535000   98.135000 ;
      RECT  28.255000   99.475000  29.535000  100.755000 ;
      RECT  50.260000   -3.260000  51.540000   -1.980000 ;
      RECT  50.260000   -0.640000  51.540000    0.640000 ;
      RECT  50.260000    1.980000  51.540000    3.260000 ;
      RECT  52.880000   -3.260000  54.160000   -1.980000 ;
      RECT  52.880000   -0.640000  54.160000    0.640000 ;
      RECT  52.880000    1.980000  54.160000    3.260000 ;
      RECT  55.650000   -3.260000  56.930000   -1.980000 ;
      RECT  55.650000   -0.640000  56.930000    0.640000 ;
      RECT  55.650000    1.980000  56.930000    3.260000 ;
  END
END sky130_fd_pr__rf_test_coil2
END LIBRARY
