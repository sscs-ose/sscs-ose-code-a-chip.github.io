* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0






.subckt sky130_fd_pr__rf_aura_blocking B_P D_N2 D_P D_P2 G G_N2 G_P G_P2 NWELL S S_N2
+ S_P S_P2 VGND VPWR
Xsky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15_0 D_P2 S_P2 G_P2 B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0 D_N2 G_N2 S_N2 SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
Xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_0 D_P S_P G_P B_P SUBS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
Xsky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0 VPWR G S SUBS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15
.ends
