# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF04W2p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF04W2p00L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  2.330000 BY  3.120000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.120000 ;
    PORT
      LAYER met3 ;
        RECT 0.570000 1.375000 0.900000 1.815000 ;
        RECT 0.570000 1.815000 1.760000 2.145000 ;
        RECT 1.430000 1.375000 1.760000 1.815000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.200000 ;
    PORT
      LAYER met1 ;
        RECT 0.480000 2.365000 1.850000 2.655000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.620000 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.445000 2.140000 -0.145000 ;
        RECT 0.190000 -0.145000 0.420000  2.105000 ;
        RECT 1.050000 -0.145000 1.280000  2.105000 ;
        RECT 1.910000 -0.145000 2.140000  2.105000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.255000 0.390000 2.105000 ;
      RECT 0.490000 2.335000 1.840000 2.675000 ;
      RECT 0.650000 0.255000 0.820000 2.105000 ;
      RECT 1.080000 0.255000 1.250000 2.105000 ;
      RECT 1.510000 0.255000 1.680000 2.105000 ;
      RECT 1.940000 0.255000 2.110000 2.105000 ;
    LAYER mcon ;
      RECT 0.220000 0.375000 0.390000 0.545000 ;
      RECT 0.220000 0.735000 0.390000 0.905000 ;
      RECT 0.220000 1.095000 0.390000 1.265000 ;
      RECT 0.220000 1.455000 0.390000 1.625000 ;
      RECT 0.220000 1.815000 0.390000 1.985000 ;
      RECT 0.540000 2.425000 0.710000 2.595000 ;
      RECT 0.650000 0.375000 0.820000 0.545000 ;
      RECT 0.650000 0.735000 0.820000 0.905000 ;
      RECT 0.650000 1.095000 0.820000 1.265000 ;
      RECT 0.650000 1.455000 0.820000 1.625000 ;
      RECT 0.650000 1.815000 0.820000 1.985000 ;
      RECT 0.900000 2.425000 1.070000 2.595000 ;
      RECT 1.080000 0.375000 1.250000 0.545000 ;
      RECT 1.080000 0.735000 1.250000 0.905000 ;
      RECT 1.080000 1.095000 1.250000 1.265000 ;
      RECT 1.080000 1.455000 1.250000 1.625000 ;
      RECT 1.080000 1.815000 1.250000 1.985000 ;
      RECT 1.260000 2.425000 1.430000 2.595000 ;
      RECT 1.510000 0.375000 1.680000 0.545000 ;
      RECT 1.510000 0.735000 1.680000 0.905000 ;
      RECT 1.510000 1.095000 1.680000 1.265000 ;
      RECT 1.510000 1.455000 1.680000 1.625000 ;
      RECT 1.510000 1.815000 1.680000 1.985000 ;
      RECT 1.620000 2.425000 1.790000 2.595000 ;
      RECT 1.940000 0.375000 2.110000 0.545000 ;
      RECT 1.940000 0.735000 2.110000 0.905000 ;
      RECT 1.940000 1.095000 2.110000 1.265000 ;
      RECT 1.940000 1.455000 2.110000 1.625000 ;
      RECT 1.940000 1.815000 2.110000 1.985000 ;
    LAYER met1 ;
      RECT 0.605000 0.255000 0.865000 2.105000 ;
      RECT 1.465000 0.255000 1.725000 2.105000 ;
    LAYER met2 ;
      RECT 0.570000 1.375000 0.900000 2.145000 ;
      RECT 1.430000 1.375000 1.760000 2.145000 ;
    LAYER via ;
      RECT 0.605000 1.470000 0.865000 1.730000 ;
      RECT 0.605000 1.790000 0.865000 2.050000 ;
      RECT 1.465000 1.470000 1.725000 1.730000 ;
      RECT 1.465000 1.790000 1.725000 2.050000 ;
    LAYER via2 ;
      RECT 0.595000 1.420000 0.875000 1.700000 ;
      RECT 0.595000 1.820000 0.875000 2.100000 ;
      RECT 1.455000 1.420000 1.735000 1.700000 ;
      RECT 1.455000 1.820000 1.735000 2.100000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF04W2p00L0p15
END LIBRARY
