MACRO SCM_NMOS_B_85279373_X8_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_85279373_X8_Y1 0 0 ;
  SIZE 29240 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 6580 27690 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 14050 260 14330 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3270 700 25970 980 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 28550 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 4115 1845 5125 ;
    LAYER M1 ;
      RECT 1595 6215 1845 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 4115 3565 5125 ;
    LAYER M1 ;
      RECT 3315 6215 3565 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 4115 5285 5125 ;
    LAYER M1 ;
      RECT 5035 6215 5285 7225 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 4115 7005 5125 ;
    LAYER M1 ;
      RECT 6755 6215 7005 7225 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 4115 8725 5125 ;
    LAYER M1 ;
      RECT 8475 6215 8725 7225 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 4115 10445 5125 ;
    LAYER M1 ;
      RECT 10195 6215 10445 7225 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 11915 4115 12165 5125 ;
    LAYER M1 ;
      RECT 11915 6215 12165 7225 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 13635 4115 13885 5125 ;
    LAYER M1 ;
      RECT 13635 6215 13885 7225 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15355 4115 15605 5125 ;
    LAYER M1 ;
      RECT 15355 6215 15605 7225 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17075 4115 17325 5125 ;
    LAYER M1 ;
      RECT 17075 6215 17325 7225 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 18795 4115 19045 5125 ;
    LAYER M1 ;
      RECT 18795 6215 19045 7225 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20515 4115 20765 5125 ;
    LAYER M1 ;
      RECT 20515 6215 20765 7225 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22235 4115 22485 5125 ;
    LAYER M1 ;
      RECT 22235 6215 22485 7225 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 23955 4115 24205 5125 ;
    LAYER M1 ;
      RECT 23955 6215 24205 7225 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M1 ;
      RECT 25675 335 25925 3865 ;
    LAYER M1 ;
      RECT 25675 4115 25925 5125 ;
    LAYER M1 ;
      RECT 25675 6215 25925 7225 ;
    LAYER M1 ;
      RECT 26535 335 26785 3865 ;
    LAYER M1 ;
      RECT 27395 335 27645 3865 ;
    LAYER M1 ;
      RECT 27395 4115 27645 5125 ;
    LAYER M1 ;
      RECT 27395 6215 27645 7225 ;
    LAYER M1 ;
      RECT 28255 335 28505 3865 ;
    LAYER M2 ;
      RECT 1550 4480 27690 4760 ;
    LAYER M2 ;
      RECT 1550 280 27690 560 ;
    LAYER V1 ;
      RECT 13675 335 13845 505 ;
    LAYER V1 ;
      RECT 13675 4535 13845 4705 ;
    LAYER V1 ;
      RECT 13675 6635 13845 6805 ;
    LAYER V1 ;
      RECT 27435 335 27605 505 ;
    LAYER V1 ;
      RECT 27435 4535 27605 4705 ;
    LAYER V1 ;
      RECT 27435 6635 27605 6805 ;
    LAYER V1 ;
      RECT 15395 335 15565 505 ;
    LAYER V1 ;
      RECT 15395 4535 15565 4705 ;
    LAYER V1 ;
      RECT 15395 6635 15565 6805 ;
    LAYER V1 ;
      RECT 1635 335 1805 505 ;
    LAYER V1 ;
      RECT 1635 4535 1805 4705 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 4535 3525 4705 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17115 4535 17285 4705 ;
    LAYER V1 ;
      RECT 17115 6635 17285 6805 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 4535 5245 4705 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 18835 4535 19005 4705 ;
    LAYER V1 ;
      RECT 18835 6635 19005 6805 ;
    LAYER V1 ;
      RECT 6795 335 6965 505 ;
    LAYER V1 ;
      RECT 6795 4535 6965 4705 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 20555 335 20725 505 ;
    LAYER V1 ;
      RECT 20555 4535 20725 4705 ;
    LAYER V1 ;
      RECT 20555 6635 20725 6805 ;
    LAYER V1 ;
      RECT 25715 755 25885 925 ;
    LAYER V1 ;
      RECT 25715 4535 25885 4705 ;
    LAYER V1 ;
      RECT 25715 6635 25885 6805 ;
    LAYER V1 ;
      RECT 22275 335 22445 505 ;
    LAYER V1 ;
      RECT 22275 4535 22445 4705 ;
    LAYER V1 ;
      RECT 22275 6635 22445 6805 ;
    LAYER V1 ;
      RECT 8515 335 8685 505 ;
    LAYER V1 ;
      RECT 8515 4535 8685 4705 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 23995 4535 24165 4705 ;
    LAYER V1 ;
      RECT 23995 6635 24165 6805 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 11955 4535 12125 4705 ;
    LAYER V1 ;
      RECT 11955 6635 12125 6805 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 10235 4535 10405 4705 ;
    LAYER V1 ;
      RECT 10235 6635 10405 6805 ;
    LAYER V1 ;
      RECT 28295 1175 28465 1345 ;
    LAYER V1 ;
      RECT 14535 1175 14705 1345 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 16255 1175 16425 1345 ;
    LAYER V1 ;
      RECT 24855 1175 25025 1345 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 17975 1175 18145 1345 ;
    LAYER V1 ;
      RECT 19695 1175 19865 1345 ;
    LAYER V1 ;
      RECT 5935 1175 6105 1345 ;
    LAYER V1 ;
      RECT 21415 1175 21585 1345 ;
    LAYER V1 ;
      RECT 7655 1175 7825 1345 ;
    LAYER V1 ;
      RECT 23135 1175 23305 1345 ;
    LAYER V1 ;
      RECT 9375 1175 9545 1345 ;
    LAYER V1 ;
      RECT 11095 1175 11265 1345 ;
    LAYER V1 ;
      RECT 12815 1175 12985 1345 ;
    LAYER V1 ;
      RECT 26575 1175 26745 1345 ;
    LAYER V2 ;
      RECT 14115 345 14265 495 ;
    LAYER V2 ;
      RECT 14115 4545 14265 4695 ;
  END
END SCM_NMOS_B_85279373_X8_Y1
