# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  4.050000 BY  2.800000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.881600 ;
    PORT
      LAYER met3 ;
        RECT 0.570000 1.055000 0.900000 1.495000 ;
        RECT 0.570000 1.495000 3.480000 1.825000 ;
        RECT 1.430000 1.055000 1.760000 1.495000 ;
        RECT 2.290000 1.055000 2.620000 1.495000 ;
        RECT 3.150000 1.055000 3.480000 1.495000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  2.016000 ;
    PORT
      LAYER met1 ;
        RECT 0.620000 2.045000 3.430000 2.335000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.301600 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.445000 3.860000 -0.145000 ;
        RECT 0.190000 -0.145000 0.420000  1.785000 ;
        RECT 1.050000 -0.145000 1.280000  1.785000 ;
        RECT 1.910000 -0.145000 2.140000  1.785000 ;
        RECT 2.770000 -0.145000 3.000000  1.785000 ;
        RECT 3.630000 -0.145000 3.860000  1.785000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.255000 0.390000 1.785000 ;
      RECT 0.650000 0.255000 0.820000 1.785000 ;
      RECT 0.670000 2.015000 3.380000 2.355000 ;
      RECT 1.080000 0.255000 1.250000 1.785000 ;
      RECT 1.510000 0.255000 1.680000 1.785000 ;
      RECT 1.940000 0.255000 2.110000 1.785000 ;
      RECT 2.370000 0.255000 2.540000 1.785000 ;
      RECT 2.800000 0.255000 2.970000 1.785000 ;
      RECT 3.230000 0.255000 3.400000 1.785000 ;
      RECT 3.660000 0.255000 3.830000 1.785000 ;
    LAYER mcon ;
      RECT 0.220000 0.395000 0.390000 0.565000 ;
      RECT 0.220000 0.755000 0.390000 0.925000 ;
      RECT 0.220000 1.115000 0.390000 1.285000 ;
      RECT 0.220000 1.475000 0.390000 1.645000 ;
      RECT 0.650000 0.395000 0.820000 0.565000 ;
      RECT 0.650000 0.755000 0.820000 0.925000 ;
      RECT 0.650000 1.115000 0.820000 1.285000 ;
      RECT 0.650000 1.475000 0.820000 1.645000 ;
      RECT 0.680000 2.105000 0.850000 2.275000 ;
      RECT 1.040000 2.105000 1.210000 2.275000 ;
      RECT 1.080000 0.395000 1.250000 0.565000 ;
      RECT 1.080000 0.755000 1.250000 0.925000 ;
      RECT 1.080000 1.115000 1.250000 1.285000 ;
      RECT 1.080000 1.475000 1.250000 1.645000 ;
      RECT 1.400000 2.105000 1.570000 2.275000 ;
      RECT 1.510000 0.395000 1.680000 0.565000 ;
      RECT 1.510000 0.755000 1.680000 0.925000 ;
      RECT 1.510000 1.115000 1.680000 1.285000 ;
      RECT 1.510000 1.475000 1.680000 1.645000 ;
      RECT 1.760000 2.105000 1.930000 2.275000 ;
      RECT 1.940000 0.395000 2.110000 0.565000 ;
      RECT 1.940000 0.755000 2.110000 0.925000 ;
      RECT 1.940000 1.115000 2.110000 1.285000 ;
      RECT 1.940000 1.475000 2.110000 1.645000 ;
      RECT 2.120000 2.105000 2.290000 2.275000 ;
      RECT 2.370000 0.395000 2.540000 0.565000 ;
      RECT 2.370000 0.755000 2.540000 0.925000 ;
      RECT 2.370000 1.115000 2.540000 1.285000 ;
      RECT 2.370000 1.475000 2.540000 1.645000 ;
      RECT 2.480000 2.105000 2.650000 2.275000 ;
      RECT 2.800000 0.395000 2.970000 0.565000 ;
      RECT 2.800000 0.755000 2.970000 0.925000 ;
      RECT 2.800000 1.115000 2.970000 1.285000 ;
      RECT 2.800000 1.475000 2.970000 1.645000 ;
      RECT 2.840000 2.105000 3.010000 2.275000 ;
      RECT 3.200000 2.105000 3.370000 2.275000 ;
      RECT 3.230000 0.395000 3.400000 0.565000 ;
      RECT 3.230000 0.755000 3.400000 0.925000 ;
      RECT 3.230000 1.115000 3.400000 1.285000 ;
      RECT 3.230000 1.475000 3.400000 1.645000 ;
      RECT 3.660000 0.395000 3.830000 0.565000 ;
      RECT 3.660000 0.755000 3.830000 0.925000 ;
      RECT 3.660000 1.115000 3.830000 1.285000 ;
      RECT 3.660000 1.475000 3.830000 1.645000 ;
    LAYER met1 ;
      RECT 0.605000 0.255000 0.865000 1.785000 ;
      RECT 1.465000 0.255000 1.725000 1.785000 ;
      RECT 2.325000 0.255000 2.585000 1.785000 ;
      RECT 3.185000 0.255000 3.445000 1.785000 ;
    LAYER met2 ;
      RECT 0.570000 1.055000 0.900000 1.825000 ;
      RECT 1.430000 1.055000 1.760000 1.825000 ;
      RECT 2.290000 1.055000 2.620000 1.825000 ;
      RECT 3.150000 1.055000 3.480000 1.825000 ;
    LAYER via ;
      RECT 0.605000 1.150000 0.865000 1.410000 ;
      RECT 0.605000 1.470000 0.865000 1.730000 ;
      RECT 1.465000 1.150000 1.725000 1.410000 ;
      RECT 1.465000 1.470000 1.725000 1.730000 ;
      RECT 2.325000 1.150000 2.585000 1.410000 ;
      RECT 2.325000 1.470000 2.585000 1.730000 ;
      RECT 3.185000 1.150000 3.445000 1.410000 ;
      RECT 3.185000 1.470000 3.445000 1.730000 ;
    LAYER via2 ;
      RECT 0.595000 1.100000 0.875000 1.380000 ;
      RECT 0.595000 1.500000 0.875000 1.780000 ;
      RECT 1.455000 1.100000 1.735000 1.380000 ;
      RECT 1.455000 1.500000 1.735000 1.780000 ;
      RECT 2.315000 1.100000 2.595000 1.380000 ;
      RECT 2.315000 1.500000 2.595000 1.780000 ;
      RECT 3.175000 1.100000 3.455000 1.380000 ;
      RECT 3.175000 1.500000 3.455000 1.780000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15
END LIBRARY
