# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.680000 BY  6.070000 ;
  PIN BULK
    ANTENNADIFFAREA  2.929000 ;
    PORT
      LAYER li1 ;
        RECT 0.240000 0.610000 0.410000 5.460000 ;
        RECT 2.270000 0.610000 2.440000 5.460000 ;
      LAYER mcon ;
        RECT 0.240000 0.970000 0.410000 1.140000 ;
        RECT 0.240000 1.330000 0.410000 1.500000 ;
        RECT 0.240000 1.690000 0.410000 1.860000 ;
        RECT 0.240000 2.050000 0.410000 2.220000 ;
        RECT 0.240000 2.410000 0.410000 2.580000 ;
        RECT 0.240000 2.770000 0.410000 2.940000 ;
        RECT 0.240000 3.130000 0.410000 3.300000 ;
        RECT 0.240000 3.490000 0.410000 3.660000 ;
        RECT 0.240000 3.850000 0.410000 4.020000 ;
        RECT 0.240000 4.210000 0.410000 4.380000 ;
        RECT 0.240000 4.570000 0.410000 4.740000 ;
        RECT 0.240000 4.930000 0.410000 5.100000 ;
        RECT 0.240000 5.290000 0.410000 5.460000 ;
        RECT 2.270000 0.970000 2.440000 1.140000 ;
        RECT 2.270000 1.330000 2.440000 1.500000 ;
        RECT 2.270000 1.690000 2.440000 1.860000 ;
        RECT 2.270000 2.050000 2.440000 2.220000 ;
        RECT 2.270000 2.410000 2.440000 2.580000 ;
        RECT 2.270000 2.770000 2.440000 2.940000 ;
        RECT 2.270000 3.130000 2.440000 3.300000 ;
        RECT 2.270000 3.490000 2.440000 3.660000 ;
        RECT 2.270000 3.850000 2.440000 4.020000 ;
        RECT 2.270000 4.210000 2.440000 4.380000 ;
        RECT 2.270000 4.570000 2.440000 4.740000 ;
        RECT 2.270000 4.930000 2.440000 5.100000 ;
        RECT 2.270000 5.290000 2.440000 5.460000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.180000 0.550000 0.470000 5.520000 ;
        RECT 2.210000 0.550000 2.500000 5.520000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  1.414000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 3.160000 2.630000 5.520000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.818000 ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.100000 1.845000 0.270000 ;
        RECT 0.835000 5.800000 1.845000 5.970000 ;
      LAYER mcon ;
        RECT 0.895000 0.100000 1.065000 0.270000 ;
        RECT 0.895000 5.800000 1.065000 5.970000 ;
        RECT 1.255000 0.100000 1.425000 0.270000 ;
        RECT 1.255000 5.800000 1.425000 5.970000 ;
        RECT 1.615000 0.100000 1.785000 0.270000 ;
        RECT 1.615000 5.800000 1.785000 5.970000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.835000 0.000000 1.845000 0.330000 ;
        RECT 0.835000 5.740000 1.845000 6.070000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.550000 2.630000 2.910000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.795000 0.490000 0.965000 5.580000 ;
      RECT 1.255000 0.490000 1.425000 5.580000 ;
      RECT 1.715000 0.490000 1.885000 5.580000 ;
    LAYER mcon ;
      RECT 0.795000 0.610000 0.965000 0.780000 ;
      RECT 0.795000 0.970000 0.965000 1.140000 ;
      RECT 0.795000 1.330000 0.965000 1.500000 ;
      RECT 0.795000 1.690000 0.965000 1.860000 ;
      RECT 0.795000 2.050000 0.965000 2.220000 ;
      RECT 0.795000 2.410000 0.965000 2.580000 ;
      RECT 0.795000 2.770000 0.965000 2.940000 ;
      RECT 0.795000 3.130000 0.965000 3.300000 ;
      RECT 0.795000 3.490000 0.965000 3.660000 ;
      RECT 0.795000 3.850000 0.965000 4.020000 ;
      RECT 0.795000 4.210000 0.965000 4.380000 ;
      RECT 0.795000 4.570000 0.965000 4.740000 ;
      RECT 0.795000 4.930000 0.965000 5.100000 ;
      RECT 0.795000 5.290000 0.965000 5.460000 ;
      RECT 1.255000 0.610000 1.425000 0.780000 ;
      RECT 1.255000 0.970000 1.425000 1.140000 ;
      RECT 1.255000 1.330000 1.425000 1.500000 ;
      RECT 1.255000 1.690000 1.425000 1.860000 ;
      RECT 1.255000 2.050000 1.425000 2.220000 ;
      RECT 1.255000 2.410000 1.425000 2.580000 ;
      RECT 1.255000 2.770000 1.425000 2.940000 ;
      RECT 1.255000 3.130000 1.425000 3.300000 ;
      RECT 1.255000 3.490000 1.425000 3.660000 ;
      RECT 1.255000 3.850000 1.425000 4.020000 ;
      RECT 1.255000 4.210000 1.425000 4.380000 ;
      RECT 1.255000 4.570000 1.425000 4.740000 ;
      RECT 1.255000 4.930000 1.425000 5.100000 ;
      RECT 1.255000 5.290000 1.425000 5.460000 ;
      RECT 1.715000 0.610000 1.885000 0.780000 ;
      RECT 1.715000 0.970000 1.885000 1.140000 ;
      RECT 1.715000 1.330000 1.885000 1.500000 ;
      RECT 1.715000 1.690000 1.885000 1.860000 ;
      RECT 1.715000 2.050000 1.885000 2.220000 ;
      RECT 1.715000 2.410000 1.885000 2.580000 ;
      RECT 1.715000 2.770000 1.885000 2.940000 ;
      RECT 1.715000 3.130000 1.885000 3.300000 ;
      RECT 1.715000 3.490000 1.885000 3.660000 ;
      RECT 1.715000 3.850000 1.885000 4.020000 ;
      RECT 1.715000 4.210000 1.885000 4.380000 ;
      RECT 1.715000 4.570000 1.885000 4.740000 ;
      RECT 1.715000 4.930000 1.885000 5.100000 ;
      RECT 1.715000 5.290000 1.885000 5.460000 ;
    LAYER met1 ;
      RECT 0.750000 0.550000 1.010000 5.520000 ;
      RECT 1.210000 0.550000 1.470000 5.520000 ;
      RECT 1.670000 0.550000 1.930000 5.520000 ;
    LAYER via ;
      RECT 0.750000 0.580000 1.010000 0.840000 ;
      RECT 0.750000 0.900000 1.010000 1.160000 ;
      RECT 0.750000 1.220000 1.010000 1.480000 ;
      RECT 0.750000 1.540000 1.010000 1.800000 ;
      RECT 0.750000 1.860000 1.010000 2.120000 ;
      RECT 0.750000 2.180000 1.010000 2.440000 ;
      RECT 0.750000 2.500000 1.010000 2.760000 ;
      RECT 1.210000 3.310000 1.470000 3.570000 ;
      RECT 1.210000 3.630000 1.470000 3.890000 ;
      RECT 1.210000 3.950000 1.470000 4.210000 ;
      RECT 1.210000 4.270000 1.470000 4.530000 ;
      RECT 1.210000 4.590000 1.470000 4.850000 ;
      RECT 1.210000 4.910000 1.470000 5.170000 ;
      RECT 1.210000 5.230000 1.470000 5.490000 ;
      RECT 1.670000 0.580000 1.930000 0.840000 ;
      RECT 1.670000 0.900000 1.930000 1.160000 ;
      RECT 1.670000 1.220000 1.930000 1.480000 ;
      RECT 1.670000 1.540000 1.930000 1.800000 ;
      RECT 1.670000 1.860000 1.930000 2.120000 ;
      RECT 1.670000 2.180000 1.930000 2.440000 ;
      RECT 1.670000 2.500000 1.930000 2.760000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18
END LIBRARY
