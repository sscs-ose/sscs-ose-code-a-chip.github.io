MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 29.83 BY 27.64 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 12.76 2.78 13.04 13.18 ;
      LAYER M3 ;
        RECT 16.2 2.78 16.48 8.98 ;
      LAYER M3 ;
        RECT 12.76 6.115 13.04 6.485 ;
      LAYER M2 ;
        RECT 12.9 6.16 16.34 6.44 ;
      LAYER M3 ;
        RECT 16.2 6.115 16.48 6.485 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 18.35 20.42 18.63 26.62 ;
      LAYER M3 ;
        RECT 24.8 14.54 25.08 26.62 ;
      LAYER M3 ;
        RECT 18.35 21.655 18.63 22.025 ;
      LAYER M2 ;
        RECT 18.49 21.7 24.94 21.98 ;
      LAYER M3 ;
        RECT 24.8 21.655 25.08 22.025 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 19.64 2.78 19.92 8.98 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 9.32 2.78 9.6 8.98 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 4.16 14.54 4.44 26.62 ;
  LAYER M3 ;
        RECT 11.04 16.22 11.32 26.62 ;
  LAYER M3 ;
        RECT 17.92 16.22 18.2 22.42 ;
  LAYER M3 ;
        RECT 4.16 19.975 4.44 20.345 ;
  LAYER M4 ;
        RECT 4.3 19.76 11.18 20.56 ;
  LAYER M3 ;
        RECT 11.04 19.975 11.32 20.345 ;
  LAYER M4 ;
        RECT 11.18 19.76 18.06 20.56 ;
  LAYER M3 ;
        RECT 17.92 19.975 18.2 20.345 ;
  LAYER M3 ;
        RECT 4.16 19.975 4.44 20.345 ;
  LAYER M4 ;
        RECT 4.135 19.76 4.465 20.56 ;
  LAYER M3 ;
        RECT 11.04 19.975 11.32 20.345 ;
  LAYER M4 ;
        RECT 11.015 19.76 11.345 20.56 ;
  LAYER M3 ;
        RECT 4.16 19.975 4.44 20.345 ;
  LAYER M4 ;
        RECT 4.135 19.76 4.465 20.56 ;
  LAYER M3 ;
        RECT 11.04 19.975 11.32 20.345 ;
  LAYER M4 ;
        RECT 11.015 19.76 11.345 20.56 ;
  LAYER M3 ;
        RECT 4.16 19.975 4.44 20.345 ;
  LAYER M4 ;
        RECT 4.135 19.76 4.465 20.56 ;
  LAYER M3 ;
        RECT 11.04 19.975 11.32 20.345 ;
  LAYER M4 ;
        RECT 11.015 19.76 11.345 20.56 ;
  LAYER M3 ;
        RECT 17.92 19.975 18.2 20.345 ;
  LAYER M4 ;
        RECT 17.895 19.76 18.225 20.56 ;
  LAYER M3 ;
        RECT 4.16 19.975 4.44 20.345 ;
  LAYER M4 ;
        RECT 4.135 19.76 4.465 20.56 ;
  LAYER M3 ;
        RECT 11.04 19.975 11.32 20.345 ;
  LAYER M4 ;
        RECT 11.015 19.76 11.345 20.56 ;
  LAYER M3 ;
        RECT 17.92 19.975 18.2 20.345 ;
  LAYER M4 ;
        RECT 17.895 19.76 18.225 20.56 ;
  LAYER M3 ;
        RECT 24.8 2.78 25.08 7.3 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 13.18 ;
  LAYER M3 ;
        RECT 25.23 10.34 25.51 22.42 ;
  LAYER M3 ;
        RECT 24.8 7.14 25.08 7.56 ;
  LAYER M2 ;
        RECT 20.21 7.42 24.94 7.7 ;
  LAYER M3 ;
        RECT 20.07 7.375 20.35 7.745 ;
  LAYER M2 ;
        RECT 24.94 7.42 25.37 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.56 25.51 10.5 ;
  LAYER M2 ;
        RECT 20.05 7.42 20.37 7.7 ;
  LAYER M3 ;
        RECT 20.07 7.4 20.35 7.72 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 20.05 7.42 20.37 7.7 ;
  LAYER M3 ;
        RECT 20.07 7.4 20.35 7.72 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 20.05 7.42 20.37 7.7 ;
  LAYER M3 ;
        RECT 20.07 7.4 20.35 7.72 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 20.05 7.42 20.37 7.7 ;
  LAYER M3 ;
        RECT 20.07 7.4 20.35 7.72 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M3 ;
        RECT 4.16 2.78 4.44 7.3 ;
  LAYER M3 ;
        RECT 8.89 6.98 9.17 13.18 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 22.42 ;
  LAYER M3 ;
        RECT 4.16 7.14 4.44 7.56 ;
  LAYER M2 ;
        RECT 4.3 7.42 9.03 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.375 9.17 7.745 ;
  LAYER M2 ;
        RECT 3.87 7.42 4.3 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.56 4.01 10.5 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M2 ;
        RECT 3.71 7.42 4.03 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.4 4.01 7.72 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M2 ;
        RECT 3.71 7.42 4.03 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.4 4.01 7.72 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 8.87 7.42 9.19 7.7 ;
  LAYER M3 ;
        RECT 8.89 7.4 9.17 7.72 ;
  LAYER M3 ;
        RECT 9.75 6.56 10.03 12.76 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M3 ;
        RECT 19.21 6.56 19.49 12.76 ;
  LAYER M3 ;
        RECT 9.75 9.475 10.03 9.845 ;
  LAYER M2 ;
        RECT 9.89 9.52 15.91 9.8 ;
  LAYER M3 ;
        RECT 15.77 9.475 16.05 9.845 ;
  LAYER M2 ;
        RECT 15.91 9.52 19.35 9.8 ;
  LAYER M3 ;
        RECT 19.21 9.475 19.49 9.845 ;
  LAYER M2 ;
        RECT 9.73 9.52 10.05 9.8 ;
  LAYER M3 ;
        RECT 9.75 9.5 10.03 9.82 ;
  LAYER M2 ;
        RECT 15.75 9.52 16.07 9.8 ;
  LAYER M3 ;
        RECT 15.77 9.5 16.05 9.82 ;
  LAYER M2 ;
        RECT 9.73 9.52 10.05 9.8 ;
  LAYER M3 ;
        RECT 9.75 9.5 10.03 9.82 ;
  LAYER M2 ;
        RECT 15.75 9.52 16.07 9.8 ;
  LAYER M3 ;
        RECT 15.77 9.5 16.05 9.82 ;
  LAYER M2 ;
        RECT 9.73 9.52 10.05 9.8 ;
  LAYER M3 ;
        RECT 9.75 9.5 10.03 9.82 ;
  LAYER M2 ;
        RECT 15.75 9.52 16.07 9.8 ;
  LAYER M3 ;
        RECT 15.77 9.5 16.05 9.82 ;
  LAYER M2 ;
        RECT 19.19 9.52 19.51 9.8 ;
  LAYER M3 ;
        RECT 19.21 9.5 19.49 9.82 ;
  LAYER M2 ;
        RECT 9.73 9.52 10.05 9.8 ;
  LAYER M3 ;
        RECT 9.75 9.5 10.03 9.82 ;
  LAYER M2 ;
        RECT 15.75 9.52 16.07 9.8 ;
  LAYER M3 ;
        RECT 15.77 9.5 16.05 9.82 ;
  LAYER M2 ;
        RECT 19.19 9.52 19.51 9.8 ;
  LAYER M3 ;
        RECT 19.21 9.5 19.49 9.82 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 9.575 12.595 13.105 ;
  LAYER M1 ;
        RECT 12.345 8.315 12.595 9.325 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 9.575 12.165 13.105 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M2 ;
        RECT 12.3 8.68 13.5 8.96 ;
  LAYER M2 ;
        RECT 12.3 12.88 13.5 13.16 ;
  LAYER M2 ;
        RECT 11.87 12.46 13.93 12.74 ;
  LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 11.87 6.58 13.93 6.86 ;
  LAYER M2 ;
        RECT 12.3 0.7 13.5 0.98 ;
  LAYER M3 ;
        RECT 12.76 2.78 13.04 13.18 ;
  LAYER M3 ;
        RECT 12.33 0.68 12.61 12.76 ;
  LAYER M1 ;
        RECT 8.905 23.015 9.155 26.545 ;
  LAYER M1 ;
        RECT 8.905 21.755 9.155 22.765 ;
  LAYER M1 ;
        RECT 8.905 17.135 9.155 20.665 ;
  LAYER M1 ;
        RECT 8.905 15.875 9.155 16.885 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 23.015 8.725 26.545 ;
  LAYER M1 ;
        RECT 8.475 17.135 8.725 20.665 ;
  LAYER M1 ;
        RECT 9.335 23.015 9.585 26.545 ;
  LAYER M1 ;
        RECT 9.335 17.135 9.585 20.665 ;
  LAYER M1 ;
        RECT 9.765 23.015 10.015 26.545 ;
  LAYER M1 ;
        RECT 9.765 21.755 10.015 22.765 ;
  LAYER M1 ;
        RECT 9.765 17.135 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.765 15.875 10.015 16.885 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 23.015 10.445 26.545 ;
  LAYER M1 ;
        RECT 10.195 17.135 10.445 20.665 ;
  LAYER M1 ;
        RECT 10.625 23.015 10.875 26.545 ;
  LAYER M1 ;
        RECT 10.625 21.755 10.875 22.765 ;
  LAYER M1 ;
        RECT 10.625 17.135 10.875 20.665 ;
  LAYER M1 ;
        RECT 10.625 15.875 10.875 16.885 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 23.015 11.305 26.545 ;
  LAYER M1 ;
        RECT 11.055 17.135 11.305 20.665 ;
  LAYER M1 ;
        RECT 11.485 23.015 11.735 26.545 ;
  LAYER M1 ;
        RECT 11.485 21.755 11.735 22.765 ;
  LAYER M1 ;
        RECT 11.485 17.135 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.485 15.875 11.735 16.885 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 23.015 12.165 26.545 ;
  LAYER M1 ;
        RECT 11.915 17.135 12.165 20.665 ;
  LAYER M1 ;
        RECT 12.345 23.015 12.595 26.545 ;
  LAYER M1 ;
        RECT 12.345 21.755 12.595 22.765 ;
  LAYER M1 ;
        RECT 12.345 17.135 12.595 20.665 ;
  LAYER M1 ;
        RECT 12.345 15.875 12.595 16.885 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 14.785 ;
  LAYER M1 ;
        RECT 12.775 23.015 13.025 26.545 ;
  LAYER M1 ;
        RECT 12.775 17.135 13.025 20.665 ;
  LAYER M1 ;
        RECT 13.205 23.015 13.455 26.545 ;
  LAYER M1 ;
        RECT 13.205 21.755 13.455 22.765 ;
  LAYER M1 ;
        RECT 13.205 17.135 13.455 20.665 ;
  LAYER M1 ;
        RECT 13.205 15.875 13.455 16.885 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.635 23.015 13.885 26.545 ;
  LAYER M1 ;
        RECT 13.635 17.135 13.885 20.665 ;
  LAYER M2 ;
        RECT 8.86 22.12 13.5 22.4 ;
  LAYER M2 ;
        RECT 8.86 26.32 13.5 26.6 ;
  LAYER M2 ;
        RECT 8.43 25.9 13.93 26.18 ;
  LAYER M2 ;
        RECT 8.86 16.24 13.5 16.52 ;
  LAYER M2 ;
        RECT 8.86 20.44 13.5 20.72 ;
  LAYER M2 ;
        RECT 8.43 20.02 13.93 20.3 ;
  LAYER M2 ;
        RECT 8.86 14.14 13.5 14.42 ;
  LAYER M3 ;
        RECT 11.04 16.22 11.32 26.62 ;
  LAYER M3 ;
        RECT 11.47 14.12 11.75 26.2 ;
  LAYER M1 ;
        RECT 26.965 3.695 27.215 7.225 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 1.345 ;
  LAYER M1 ;
        RECT 27.395 3.695 27.645 7.225 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 23.525 3.695 23.775 7.225 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.525 0.335 23.775 1.345 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M2 ;
        RECT 22.62 2.8 27.26 3.08 ;
  LAYER M2 ;
        RECT 22.62 7 27.26 7.28 ;
  LAYER M2 ;
        RECT 22.19 6.58 27.69 6.86 ;
  LAYER M2 ;
        RECT 22.62 0.7 27.26 0.98 ;
  LAYER M3 ;
        RECT 24.8 2.78 25.08 7.3 ;
  LAYER M3 ;
        RECT 24.37 0.68 24.65 6.88 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 1.98 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 1.98 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 1.55 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 1.98 0.7 6.62 0.98 ;
  LAYER M3 ;
        RECT 4.16 2.78 4.44 7.3 ;
  LAYER M3 ;
        RECT 4.59 0.68 4.87 6.88 ;
  LAYER M1 ;
        RECT 20.085 23.015 20.335 26.545 ;
  LAYER M1 ;
        RECT 20.085 21.755 20.335 22.765 ;
  LAYER M1 ;
        RECT 20.085 17.135 20.335 20.665 ;
  LAYER M1 ;
        RECT 20.085 15.875 20.335 16.885 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 14.785 ;
  LAYER M1 ;
        RECT 20.515 23.015 20.765 26.545 ;
  LAYER M1 ;
        RECT 20.515 17.135 20.765 20.665 ;
  LAYER M1 ;
        RECT 19.655 23.015 19.905 26.545 ;
  LAYER M1 ;
        RECT 19.655 17.135 19.905 20.665 ;
  LAYER M1 ;
        RECT 19.225 23.015 19.475 26.545 ;
  LAYER M1 ;
        RECT 19.225 21.755 19.475 22.765 ;
  LAYER M1 ;
        RECT 19.225 17.135 19.475 20.665 ;
  LAYER M1 ;
        RECT 19.225 15.875 19.475 16.885 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 18.795 23.015 19.045 26.545 ;
  LAYER M1 ;
        RECT 18.795 17.135 19.045 20.665 ;
  LAYER M1 ;
        RECT 18.365 23.015 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.365 21.755 18.615 22.765 ;
  LAYER M1 ;
        RECT 18.365 17.135 18.615 20.665 ;
  LAYER M1 ;
        RECT 18.365 15.875 18.615 16.885 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 14.785 ;
  LAYER M1 ;
        RECT 17.935 23.015 18.185 26.545 ;
  LAYER M1 ;
        RECT 17.935 17.135 18.185 20.665 ;
  LAYER M1 ;
        RECT 17.505 23.015 17.755 26.545 ;
  LAYER M1 ;
        RECT 17.505 21.755 17.755 22.765 ;
  LAYER M1 ;
        RECT 17.505 17.135 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.505 15.875 17.755 16.885 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.075 23.015 17.325 26.545 ;
  LAYER M1 ;
        RECT 17.075 17.135 17.325 20.665 ;
  LAYER M1 ;
        RECT 16.645 23.015 16.895 26.545 ;
  LAYER M1 ;
        RECT 16.645 21.755 16.895 22.765 ;
  LAYER M1 ;
        RECT 16.645 17.135 16.895 20.665 ;
  LAYER M1 ;
        RECT 16.645 15.875 16.895 16.885 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 16.215 23.015 16.465 26.545 ;
  LAYER M1 ;
        RECT 16.215 17.135 16.465 20.665 ;
  LAYER M1 ;
        RECT 15.785 23.015 16.035 26.545 ;
  LAYER M1 ;
        RECT 15.785 21.755 16.035 22.765 ;
  LAYER M1 ;
        RECT 15.785 17.135 16.035 20.665 ;
  LAYER M1 ;
        RECT 15.785 15.875 16.035 16.885 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 14.785 ;
  LAYER M1 ;
        RECT 15.355 23.015 15.605 26.545 ;
  LAYER M1 ;
        RECT 15.355 17.135 15.605 20.665 ;
  LAYER M2 ;
        RECT 15.74 26.32 20.38 26.6 ;
  LAYER M2 ;
        RECT 15.74 22.12 20.38 22.4 ;
  LAYER M2 ;
        RECT 15.31 25.9 20.81 26.18 ;
  LAYER M2 ;
        RECT 15.74 20.44 20.38 20.72 ;
  LAYER M2 ;
        RECT 15.74 16.24 20.38 16.52 ;
  LAYER M2 ;
        RECT 15.31 20.02 20.81 20.3 ;
  LAYER M2 ;
        RECT 15.74 14.14 20.38 14.42 ;
  LAYER M3 ;
        RECT 18.35 20.42 18.63 26.62 ;
  LAYER M3 ;
        RECT 17.92 16.22 18.2 22.42 ;
  LAYER M3 ;
        RECT 17.49 14.12 17.77 26.2 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 16.645 9.575 16.895 13.105 ;
  LAYER M1 ;
        RECT 16.645 8.315 16.895 9.325 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M2 ;
        RECT 15.74 12.88 16.94 13.16 ;
  LAYER M2 ;
        RECT 15.74 8.68 16.94 8.96 ;
  LAYER M2 ;
        RECT 15.31 12.46 17.37 12.74 ;
  LAYER M2 ;
        RECT 15.74 7 16.94 7.28 ;
  LAYER M2 ;
        RECT 15.74 2.8 16.94 3.08 ;
  LAYER M2 ;
        RECT 15.31 6.58 17.37 6.86 ;
  LAYER M2 ;
        RECT 15.74 0.7 16.94 0.98 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M3 ;
        RECT 16.2 2.78 16.48 8.98 ;
  LAYER M3 ;
        RECT 16.63 0.68 16.91 12.76 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 6.325 21.755 6.575 22.765 ;
  LAYER M1 ;
        RECT 6.325 17.135 6.575 20.665 ;
  LAYER M1 ;
        RECT 6.325 15.875 6.575 16.885 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 6.755 17.135 7.005 20.665 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M1 ;
        RECT 5.895 17.135 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 5.465 23.015 5.715 26.545 ;
  LAYER M1 ;
        RECT 5.465 21.755 5.715 22.765 ;
  LAYER M1 ;
        RECT 5.465 17.135 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.465 15.875 5.715 16.885 ;
  LAYER M1 ;
        RECT 5.465 11.255 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.465 9.995 5.715 11.005 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.905 ;
  LAYER M1 ;
        RECT 5.035 23.015 5.285 26.545 ;
  LAYER M1 ;
        RECT 5.035 17.135 5.285 20.665 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 26.545 ;
  LAYER M1 ;
        RECT 4.605 21.755 4.855 22.765 ;
  LAYER M1 ;
        RECT 4.605 17.135 4.855 20.665 ;
  LAYER M1 ;
        RECT 4.605 15.875 4.855 16.885 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M1 ;
        RECT 4.175 17.135 4.425 20.665 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 21.755 3.995 22.765 ;
  LAYER M1 ;
        RECT 3.745 17.135 3.995 20.665 ;
  LAYER M1 ;
        RECT 3.745 15.875 3.995 16.885 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M1 ;
        RECT 3.315 17.135 3.565 20.665 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 2.885 23.015 3.135 26.545 ;
  LAYER M1 ;
        RECT 2.885 21.755 3.135 22.765 ;
  LAYER M1 ;
        RECT 2.885 17.135 3.135 20.665 ;
  LAYER M1 ;
        RECT 2.885 15.875 3.135 16.885 ;
  LAYER M1 ;
        RECT 2.885 11.255 3.135 14.785 ;
  LAYER M1 ;
        RECT 2.885 9.995 3.135 11.005 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.905 ;
  LAYER M1 ;
        RECT 2.455 23.015 2.705 26.545 ;
  LAYER M1 ;
        RECT 2.455 17.135 2.705 20.665 ;
  LAYER M1 ;
        RECT 2.455 11.255 2.705 14.785 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 26.545 ;
  LAYER M1 ;
        RECT 2.025 21.755 2.275 22.765 ;
  LAYER M1 ;
        RECT 2.025 17.135 2.275 20.665 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.885 ;
  LAYER M1 ;
        RECT 2.025 11.255 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.905 ;
  LAYER M1 ;
        RECT 1.595 23.015 1.845 26.545 ;
  LAYER M1 ;
        RECT 1.595 17.135 1.845 20.665 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M1 ;
        RECT 1.165 23.015 1.415 26.545 ;
  LAYER M1 ;
        RECT 1.165 21.755 1.415 22.765 ;
  LAYER M1 ;
        RECT 1.165 17.135 1.415 20.665 ;
  LAYER M1 ;
        RECT 1.165 15.875 1.415 16.885 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.165 9.995 1.415 11.005 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 8.905 ;
  LAYER M1 ;
        RECT 0.735 23.015 0.985 26.545 ;
  LAYER M1 ;
        RECT 0.735 17.135 0.985 20.665 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 1.12 26.32 6.62 26.6 ;
  LAYER M2 ;
        RECT 1.12 22.12 6.62 22.4 ;
  LAYER M2 ;
        RECT 0.69 25.9 7.05 26.18 ;
  LAYER M2 ;
        RECT 1.12 20.44 6.62 20.72 ;
  LAYER M2 ;
        RECT 1.12 16.24 6.62 16.52 ;
  LAYER M2 ;
        RECT 0.69 20.02 7.05 20.3 ;
  LAYER M2 ;
        RECT 1.12 14.56 6.62 14.84 ;
  LAYER M2 ;
        RECT 1.12 10.36 6.62 10.64 ;
  LAYER M2 ;
        RECT 0.69 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 1.12 8.26 6.62 8.54 ;
  LAYER M3 ;
        RECT 4.16 14.54 4.44 26.62 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 22.42 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 26.2 ;
  LAYER M1 ;
        RECT 22.665 23.015 22.915 26.545 ;
  LAYER M1 ;
        RECT 22.665 21.755 22.915 22.765 ;
  LAYER M1 ;
        RECT 22.665 17.135 22.915 20.665 ;
  LAYER M1 ;
        RECT 22.665 15.875 22.915 16.885 ;
  LAYER M1 ;
        RECT 22.665 11.255 22.915 14.785 ;
  LAYER M1 ;
        RECT 22.665 9.995 22.915 11.005 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 8.905 ;
  LAYER M1 ;
        RECT 22.235 23.015 22.485 26.545 ;
  LAYER M1 ;
        RECT 22.235 17.135 22.485 20.665 ;
  LAYER M1 ;
        RECT 22.235 11.255 22.485 14.785 ;
  LAYER M1 ;
        RECT 23.095 23.015 23.345 26.545 ;
  LAYER M1 ;
        RECT 23.095 17.135 23.345 20.665 ;
  LAYER M1 ;
        RECT 23.095 11.255 23.345 14.785 ;
  LAYER M1 ;
        RECT 23.525 23.015 23.775 26.545 ;
  LAYER M1 ;
        RECT 23.525 21.755 23.775 22.765 ;
  LAYER M1 ;
        RECT 23.525 17.135 23.775 20.665 ;
  LAYER M1 ;
        RECT 23.525 15.875 23.775 16.885 ;
  LAYER M1 ;
        RECT 23.525 11.255 23.775 14.785 ;
  LAYER M1 ;
        RECT 23.525 9.995 23.775 11.005 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 8.905 ;
  LAYER M1 ;
        RECT 23.955 23.015 24.205 26.545 ;
  LAYER M1 ;
        RECT 23.955 17.135 24.205 20.665 ;
  LAYER M1 ;
        RECT 23.955 11.255 24.205 14.785 ;
  LAYER M1 ;
        RECT 24.385 23.015 24.635 26.545 ;
  LAYER M1 ;
        RECT 24.385 21.755 24.635 22.765 ;
  LAYER M1 ;
        RECT 24.385 17.135 24.635 20.665 ;
  LAYER M1 ;
        RECT 24.385 15.875 24.635 16.885 ;
  LAYER M1 ;
        RECT 24.385 11.255 24.635 14.785 ;
  LAYER M1 ;
        RECT 24.385 9.995 24.635 11.005 ;
  LAYER M1 ;
        RECT 24.385 7.895 24.635 8.905 ;
  LAYER M1 ;
        RECT 24.815 23.015 25.065 26.545 ;
  LAYER M1 ;
        RECT 24.815 17.135 25.065 20.665 ;
  LAYER M1 ;
        RECT 24.815 11.255 25.065 14.785 ;
  LAYER M1 ;
        RECT 25.245 23.015 25.495 26.545 ;
  LAYER M1 ;
        RECT 25.245 21.755 25.495 22.765 ;
  LAYER M1 ;
        RECT 25.245 17.135 25.495 20.665 ;
  LAYER M1 ;
        RECT 25.245 15.875 25.495 16.885 ;
  LAYER M1 ;
        RECT 25.245 11.255 25.495 14.785 ;
  LAYER M1 ;
        RECT 25.245 9.995 25.495 11.005 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 8.905 ;
  LAYER M1 ;
        RECT 25.675 23.015 25.925 26.545 ;
  LAYER M1 ;
        RECT 25.675 17.135 25.925 20.665 ;
  LAYER M1 ;
        RECT 25.675 11.255 25.925 14.785 ;
  LAYER M1 ;
        RECT 26.105 23.015 26.355 26.545 ;
  LAYER M1 ;
        RECT 26.105 21.755 26.355 22.765 ;
  LAYER M1 ;
        RECT 26.105 17.135 26.355 20.665 ;
  LAYER M1 ;
        RECT 26.105 15.875 26.355 16.885 ;
  LAYER M1 ;
        RECT 26.105 11.255 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.105 9.995 26.355 11.005 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 8.905 ;
  LAYER M1 ;
        RECT 26.535 23.015 26.785 26.545 ;
  LAYER M1 ;
        RECT 26.535 17.135 26.785 20.665 ;
  LAYER M1 ;
        RECT 26.535 11.255 26.785 14.785 ;
  LAYER M1 ;
        RECT 26.965 23.015 27.215 26.545 ;
  LAYER M1 ;
        RECT 26.965 21.755 27.215 22.765 ;
  LAYER M1 ;
        RECT 26.965 17.135 27.215 20.665 ;
  LAYER M1 ;
        RECT 26.965 15.875 27.215 16.885 ;
  LAYER M1 ;
        RECT 26.965 11.255 27.215 14.785 ;
  LAYER M1 ;
        RECT 26.965 9.995 27.215 11.005 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 8.905 ;
  LAYER M1 ;
        RECT 27.395 23.015 27.645 26.545 ;
  LAYER M1 ;
        RECT 27.395 17.135 27.645 20.665 ;
  LAYER M1 ;
        RECT 27.395 11.255 27.645 14.785 ;
  LAYER M1 ;
        RECT 27.825 23.015 28.075 26.545 ;
  LAYER M1 ;
        RECT 27.825 21.755 28.075 22.765 ;
  LAYER M1 ;
        RECT 27.825 17.135 28.075 20.665 ;
  LAYER M1 ;
        RECT 27.825 15.875 28.075 16.885 ;
  LAYER M1 ;
        RECT 27.825 11.255 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.825 9.995 28.075 11.005 ;
  LAYER M1 ;
        RECT 27.825 7.895 28.075 8.905 ;
  LAYER M1 ;
        RECT 28.255 23.015 28.505 26.545 ;
  LAYER M1 ;
        RECT 28.255 17.135 28.505 20.665 ;
  LAYER M1 ;
        RECT 28.255 11.255 28.505 14.785 ;
  LAYER M2 ;
        RECT 22.62 26.32 28.12 26.6 ;
  LAYER M2 ;
        RECT 22.62 22.12 28.12 22.4 ;
  LAYER M2 ;
        RECT 22.19 25.9 28.55 26.18 ;
  LAYER M2 ;
        RECT 22.62 20.44 28.12 20.72 ;
  LAYER M2 ;
        RECT 22.62 16.24 28.12 16.52 ;
  LAYER M2 ;
        RECT 22.19 20.02 28.55 20.3 ;
  LAYER M2 ;
        RECT 22.62 14.56 28.12 14.84 ;
  LAYER M2 ;
        RECT 22.62 10.36 28.12 10.64 ;
  LAYER M2 ;
        RECT 22.19 14.14 28.55 14.42 ;
  LAYER M2 ;
        RECT 22.62 8.26 28.12 8.54 ;
  LAYER M3 ;
        RECT 24.8 14.54 25.08 26.62 ;
  LAYER M3 ;
        RECT 25.23 10.34 25.51 22.42 ;
  LAYER M3 ;
        RECT 25.66 8.24 25.94 26.2 ;
  LAYER M1 ;
        RECT 20.085 9.575 20.335 13.105 ;
  LAYER M1 ;
        RECT 20.085 8.315 20.335 9.325 ;
  LAYER M1 ;
        RECT 20.085 3.695 20.335 7.225 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 1.345 ;
  LAYER M1 ;
        RECT 20.515 9.575 20.765 13.105 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 19.655 9.575 19.905 13.105 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 19.225 9.575 19.475 13.105 ;
  LAYER M1 ;
        RECT 19.225 8.315 19.475 9.325 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 9.575 19.045 13.105 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M2 ;
        RECT 19.18 12.88 20.38 13.16 ;
  LAYER M2 ;
        RECT 19.18 8.68 20.38 8.96 ;
  LAYER M2 ;
        RECT 18.75 12.46 20.81 12.74 ;
  LAYER M2 ;
        RECT 19.18 7 20.38 7.28 ;
  LAYER M2 ;
        RECT 19.18 2.8 20.38 3.08 ;
  LAYER M2 ;
        RECT 18.75 6.58 20.81 6.86 ;
  LAYER M2 ;
        RECT 19.18 0.7 20.38 0.98 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 13.18 ;
  LAYER M3 ;
        RECT 19.64 2.78 19.92 8.98 ;
  LAYER M3 ;
        RECT 19.21 6.56 19.49 12.76 ;
  LAYER M1 ;
        RECT 8.905 9.575 9.155 13.105 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 9.325 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M2 ;
        RECT 8.86 12.88 10.06 13.16 ;
  LAYER M2 ;
        RECT 8.86 8.68 10.06 8.96 ;
  LAYER M2 ;
        RECT 8.43 12.46 10.49 12.74 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 8.43 6.58 10.49 6.86 ;
  LAYER M2 ;
        RECT 8.86 0.7 10.06 0.98 ;
  LAYER M3 ;
        RECT 8.89 6.98 9.17 13.18 ;
  LAYER M3 ;
        RECT 9.32 2.78 9.6 8.98 ;
  LAYER M3 ;
        RECT 9.75 6.56 10.03 12.76 ;
  END 
END CURRENT_MIRROR_OTA
