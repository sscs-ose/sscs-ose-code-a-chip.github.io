* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__pfet_g5v0d16v0 d g s b  w=5.0 l=0.66 ad=0 as=0 pd=0 ps=0.0 m=1 mf=1 nrd=0 nrs=0 sa=0.28 sb=1.19 sd=0 mult=1
.param rdiff='8.900000e+003*sky130_fd_pr__pfet_g5v0d16v0__rdiff_mult'
.param rdiff_tc1=2.500000e-003
.param rdiff_tc2=2.200000e-006
.param sb_cadfixedvalue_pvhv=1.19
* sd intentionally left out for sky130_fd_pr__pfet_g5v0d16v0 devices because poly-poly spacing not uniform in DE FET
xmain1 d1 g s b sky130_fd_pr__pfet_g5v0d16v0__base  w=w l=l ad=0 as=as pd=0 ps=ps nrd=nrd nrs=nrs m=m mult=mult sa=sa sb=sb_cadfixedvalue_pvhv
rldd d d1 '(1/w)*rdiff' tc1 = 'rdiff_tc1' tc2 = 'rdiff_tc2'
dnw1 d b sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn area='ad/2' pj='pd/2'
dnw2 d1 b sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn area='ad/2' pj='pd/2'
.ends sky130_fd_pr__pfet_g5v0d16v0
