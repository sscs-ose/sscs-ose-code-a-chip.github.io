# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  5.110000 BY  4.900000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.842800 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.575000 5.180000 3.855000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.010000 ;
    PORT
      LAYER li1 ;
        RECT 1.915000 0.000000 3.335000 0.685000 ;
        RECT 1.915000 4.215000 3.335000 4.900000 ;
      LAYER mcon ;
        RECT 2.000000 0.095000 3.250000 0.625000 ;
        RECT 2.000000 4.275000 3.250000 4.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.900000 0.000000 3.350000 0.685000 ;
        RECT 1.900000 4.215000 3.350000 4.900000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.045000 5.180000 2.325000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  3.010000 ;
    ANTENNAGATEAREA  1.505000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.045000 0.500000 3.855000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.750000 1.045000 5.045000 3.855000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 1.150000 3.975000 ;
      RECT 0.950000 0.485000 1.280000 0.815000 ;
      RECT 0.950000 0.815000 1.150000 0.925000 ;
      RECT 0.950000 3.975000 1.150000 4.085000 ;
      RECT 0.950000 4.085000 1.280000 4.415000 ;
      RECT 1.760000 0.925000 1.930000 3.975000 ;
      RECT 2.540000 0.925000 2.710000 3.975000 ;
      RECT 3.320000 0.925000 3.490000 3.975000 ;
      RECT 3.970000 0.485000 4.300000 0.815000 ;
      RECT 3.970000 4.085000 4.300000 4.415000 ;
      RECT 4.100000 0.815000 4.300000 0.925000 ;
      RECT 4.100000 0.925000 5.045000 3.975000 ;
      RECT 4.100000 3.975000 4.300000 4.085000 ;
    LAYER mcon ;
      RECT 0.300000 1.105000 0.470000 1.275000 ;
      RECT 0.300000 1.465000 0.470000 1.635000 ;
      RECT 0.300000 1.825000 0.470000 1.995000 ;
      RECT 0.300000 2.185000 0.470000 2.355000 ;
      RECT 0.300000 2.545000 0.470000 2.715000 ;
      RECT 0.300000 2.905000 0.470000 3.075000 ;
      RECT 0.300000 3.265000 0.470000 3.435000 ;
      RECT 0.300000 3.625000 0.470000 3.795000 ;
      RECT 1.760000 1.105000 1.930000 1.275000 ;
      RECT 1.760000 1.465000 1.930000 1.635000 ;
      RECT 1.760000 1.825000 1.930000 1.995000 ;
      RECT 1.760000 2.185000 1.930000 2.355000 ;
      RECT 1.760000 2.545000 1.930000 2.715000 ;
      RECT 1.760000 2.905000 1.930000 3.075000 ;
      RECT 1.760000 3.265000 1.930000 3.435000 ;
      RECT 1.760000 3.625000 1.930000 3.795000 ;
      RECT 2.540000 1.105000 2.710000 1.275000 ;
      RECT 2.540000 1.465000 2.710000 1.635000 ;
      RECT 2.540000 1.825000 2.710000 1.995000 ;
      RECT 2.540000 2.185000 2.710000 2.355000 ;
      RECT 2.540000 2.545000 2.710000 2.715000 ;
      RECT 2.540000 2.905000 2.710000 3.075000 ;
      RECT 2.540000 3.265000 2.710000 3.435000 ;
      RECT 2.540000 3.625000 2.710000 3.795000 ;
      RECT 3.320000 1.105000 3.490000 1.275000 ;
      RECT 3.320000 1.465000 3.490000 1.635000 ;
      RECT 3.320000 1.825000 3.490000 1.995000 ;
      RECT 3.320000 2.185000 3.490000 2.355000 ;
      RECT 3.320000 2.545000 3.490000 2.715000 ;
      RECT 3.320000 2.905000 3.490000 3.075000 ;
      RECT 3.320000 3.265000 3.490000 3.435000 ;
      RECT 3.320000 3.625000 3.490000 3.795000 ;
      RECT 4.780000 1.105000 4.950000 1.275000 ;
      RECT 4.780000 1.465000 4.950000 1.635000 ;
      RECT 4.780000 1.825000 4.950000 1.995000 ;
      RECT 4.780000 2.185000 4.950000 2.355000 ;
      RECT 4.780000 2.545000 4.950000 2.715000 ;
      RECT 4.780000 2.905000 4.950000 3.075000 ;
      RECT 4.780000 3.265000 4.950000 3.435000 ;
      RECT 4.780000 3.625000 4.950000 3.795000 ;
    LAYER met1 ;
      RECT 1.715000 1.045000 1.975000 3.855000 ;
      RECT 2.495000 1.045000 2.755000 3.855000 ;
      RECT 3.275000 1.045000 3.535000 3.855000 ;
    LAYER via ;
      RECT 1.715000 1.075000 1.975000 1.335000 ;
      RECT 1.715000 1.395000 1.975000 1.655000 ;
      RECT 1.715000 1.715000 1.975000 1.975000 ;
      RECT 1.715000 2.035000 1.975000 2.295000 ;
      RECT 2.495000 2.605000 2.755000 2.865000 ;
      RECT 2.495000 2.925000 2.755000 3.185000 ;
      RECT 2.495000 3.245000 2.755000 3.505000 ;
      RECT 2.495000 3.565000 2.755000 3.825000 ;
      RECT 3.275000 1.075000 3.535000 1.335000 ;
      RECT 3.275000 1.395000 3.535000 1.655000 ;
      RECT 3.275000 1.715000 3.535000 1.975000 ;
      RECT 3.275000 2.035000 3.535000 2.295000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50
END LIBRARY
