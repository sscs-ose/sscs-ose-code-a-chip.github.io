* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 40
.param
+ sky130_fd_pr__pfet_01v8_lvt__toxe_mult = 0.9635
+ sky130_fd_pr__pfet_01v8_lvt__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8_lvt__overlap_mult = 0.724
+ sky130_fd_pr__pfet_01v8_lvt__ajunction_mult = 9.3001e-1
+ sky130_fd_pr__pfet_01v8_lvt__pjunction_mult = 9.3439e-1
+ sky130_fd_pr__pfet_01v8_lvt__lint_diff = 1.21275e-8
+ sky130_fd_pr__pfet_01v8_lvt__wint_diff = -2.252e-8
+ sky130_fd_pr__pfet_01v8_lvt__dlc_diff = 2.0382e-8
+ sky130_fd_pr__pfet_01v8_lvt__dwc_diff = -2.252e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 000, W = 1.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_0 = 1.8236e-5
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_0 = 0.057962
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0 = 0.04699
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_0 = 0.1188
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_0 = 0.051281
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 001, W = 1.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_1 = 0.030016
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_1 = 6.3753e-5
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_1 = 0.053089
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1 = 0.062335
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_1 = 0.11351
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 002, W = 1.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_2 = 0.14251
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_2 = 0.034025
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_2 = -2.9718e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_2 = -0.042558
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2 = 0.068905
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 003, W = 1.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_3 = 0.12793
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_3 = 0.033467
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_3 = 5.3522e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_3 = -0.0034386
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3 = 0.060803
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 004, W = 1.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4 = 0.035185
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_4 = -5.7776e-9
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_4 = 0.039388
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_4 = -0.00015853
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4 = 2649.7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_4 = 2.0438e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 005, W = 1.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5 = 0.1099
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_5 = 1.6482e-7
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_5 = 0.036896
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_5 = -0.00012951
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5 = -24859.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_5 = 3.3037e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 006, W = 3.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_6 = 0.19249
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6 = 0.041047
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_6 = 0.04499
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_6 = 0.028443
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_6 = -0.00026304
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_6 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 007, W = 3.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_7 = 0.15046
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7 = 0.033761
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_7 = 0.085016
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_7 = 0.04862
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_7 = -0.00010679
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 008, W = 3.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_8 = 0.13976
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8 = 0.080847
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_8 = 0.067986
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_8 = 0.035894
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_8 = -0.0003169
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 009, W = 3.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_9 = 0.13129
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9 = 0.073616
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_9 = 0.080573
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_9 = 0.03877
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_9 = -0.00030083
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 010, W = 3.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_10 = -0.00028535
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10 = 0.080406
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_10 = 0.03088
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_10 = 0.074414
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_10 = 0.092733
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 011, W = 3.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_11 = -0.00036855
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11 = 6238.9
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11 = 0.040634
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_11 = 0.04248
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_11 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 012, W = 3.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_12 = 0.022657
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_12 = 0.087754
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_12 = -0.00033122
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12 = -13671.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12 = 0.052081
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_12 = -5.7847e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_12 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 013, W = 5.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_13 = 0.034147
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_13 = -0.0039669
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_13 = 0.10427
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_13 = -0.00021283
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13 = 0.06929
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 014, W = 5.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_14 = 0.03164
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_14 = -0.012
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_14 = 0.12605
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_14 = -0.00010143
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14 = 0.044427
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 015, W = 5.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_15 = 0.040581
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_15 = 0.0080084
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_15 = 0.11206
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_15 = -0.00027917
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15 = 0.090708
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 016, W = 5.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_16 = 0.041067
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_16 = 0.039408
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_16 = 0.1007
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_16 = -0.00021219
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16 = 0.078926
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 017, W = 5.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_17 = 0.034165
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_17 = 0.055625
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_17 = 0.097238
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_17 = -0.0002235
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17 = 0.079729
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 018, W = 5.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_18 = 0.035023
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_18 = -0.00012027
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18 = -9547.2
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18 = 0.019246
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 019, W = 5.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_19 = -2.3922e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_19 = 0.02131
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_19 = 0.091925
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_19 = -0.00016727
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19 = -18404.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19 = 0.032189
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 020, W = 7.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_20 = 0.022835
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_20 = 0.10505
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_20 = 0.092125
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_20 = -0.00015806
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20 = 0.042628
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 021, W = 7.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_21 = -0.00015959
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21 = 0.038854
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_21 = 0.040801
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_21 = 0.090482
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_21 = 0.10086
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 022, W = 7.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_22 = 0.16358
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_22 = 0.077614
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_22 = -0.00011519
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22 = 0.04077
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_22 = 1.3e-12
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_22 = 0.044326
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_22 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 023, W = 7.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_23 = 0.035049
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_23 = 0.0040365
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_23 = 0.11133
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_23 = -0.00016106
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23 = 0.072293
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_23 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 024, W = 7.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_24 = 0.032947
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_24 = 0.022112
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_24 = 0.11166
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_24 = -0.00013292
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24 = 0.066105
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 025, W = 7.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_25 = 0.032376
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_25 = -0.00010893
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25 = 2460.8
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25 = -0.004201
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 026, W = 7.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_26 = 0.02304
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_26 = 0.086586
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_26 = -0.00014865
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26 = -7093.1
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26 = 0.030421
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_26 = -3.0509e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 027, W = 0.42, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_27 = 5.4132e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_27 = 4.7258e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_27 = 0.044406
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_27 = 0.00040064
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27 = 0.015981
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 028, W = 0.42, L = 20.0
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_28 = -6.2589e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_28 = 2.1373e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_28 = 0.013052
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_28 = -9.9946e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28 = 0.04864
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 029, W = 0.42, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_29 = 1.1353e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_29 = 2.324e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_29 = 0.023227
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_29 = -3.4446e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29 = 0.075546
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 030, W = 0.42, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_30 = -2.424e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_30 = 2.2494e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_30 = 0.026211
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_30 = -4.4666e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30 = 0.049375
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_30 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 031, W = 0.42, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_31 = 5.9189e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_31 = 2.2715e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_31 = 0.028872
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_31 = -0.00012571
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31 = 0.088628
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 032, W = 0.42, L = 0.35
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_32 = 6.2247e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32 = -5767.1
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32 = 0.11275
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_32 = 0.045505
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 033, W = 0.42, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_33 = -6.6705e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33 = -19424.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33 = 0.059647
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_33 = 1.6932e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_33 = 2.1062e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_33 = 0.026212
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_33 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 034, W = 0.55, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_34 = 0.048415
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_34 = -8.0517e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34 = 0.089735
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_34 = 1.2734e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_34 = 3.9757e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_34 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 035, W = 0.55, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_35 = 0.043931
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_35 = -1.3776e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35 = 0.067319
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_35 = 5.6032e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_35 = 1.9598e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 036, W = 0.55, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_36 = 0.047583
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_36 = -4.5337e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36 = 0.06697
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_36 = 9.857e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_36 = 1.98e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 037, W = 0.55, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_37 = 2.1613e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_37 = 0.034954
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_37 = -8.6545e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37 = 0.057766
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_37 = 5.8275e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 038, W = 0.55, L = 0.35
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_38 = 0.032381
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_38 = 0.00013127
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38 = -394.79
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38 = -0.014067
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 039, W = 0.55, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_39 = 7.5746e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_39 = 3.4088e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_39 = 0.021853
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_39 = 0.00018882
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39 = -21675.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39 = 0.00071188
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_39 = 0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"
