* Contoh PWL sederhana
Vclkin in 0 PWL( 0.0 1.19527884e-08 1e-12 4.32203224e-08 2e-12 4.70966555e-08 4e-12 2.85073125e-08 8e-12 -2.74991319e-08 1.6e-11 -1.24993349e-09 3.2e-11 3.70983458e-08 6.4e-11 -5.80847326e-09
+ 1.28e-10 2.54935826e-08 2.28e-10 1.29570363e-09 3.28e-10 2.07153545e-08 4.28e-10 4.45328005e-09 5.28e-10 1.95803563e-08 6.28e-10 -1.01327143e-08 7.28e-10 5.12884463e-07 8.17641203e-10 -7.53987819e-05
+ 8.87939724e-10 -0.0110687568 9.63955785e-10 0.190862341 1e-09 3.41552034 1.00713579e-09 3.90025356 1.02140738e-09 4.47778749 1.04995055e-09 4.90665375 1.09557449e-09 5.00236731 1.1454732e-09 5.00057418
+ 1.21884515e-09 4.99942076 1.31884515e-09 5.00046968 1.41884515e-09 4.99963881 1.51884515e-09 5.00026755 1.61884515e-09 4.99980393 1.71884515e-09 5.00014112 1.81884515e-09 4.99989828 1.91884515e-09 5.00007243
+ 2.01884515e-09 4.99994809 2.11884515e-09 5.00003679 2.21884515e-09 4.99997367 2.31884515e-09 5.00001861 2.41884515e-09 4.99998667 2.51884515e-09 5.0000094 2.61884515e-09 4.99999325 2.71884515e-09 5.00000474
+ 2.81884515e-09 4.99999657 2.91884515e-09 5.00000238 3.01884515e-09 4.99999825 3.11884515e-09 5.00000119 3.21884515e-09 4.9999991 3.31884515e-09 5.00000059 3.41884515e-09 4.99999953 3.51884515e-09 5.00000028
+ 3.61884515e-09 4.99999975 3.71884515e-09 5.00000013 3.81884515e-09 4.99999986 3.91884515e-09 5.00000005 4.01884515e-09 4.99999991 4.11884515e-09 5.00000001 4.21884515e-09 4.99999994 4.31884515e-09 4.99999999
+ 4.41884515e-09 4.99999996 4.51884515e-09 4.99999998 4.61884515e-09 4.99999996 4.71884515e-09 4.99999998 4.81884515e-09 4.99999997 4.91884515e-09 4.99999997 5.01884515e-09 4.99999997 5.11884515e-09 4.99999997
+ 5.21884515e-09 4.99999997 5.31884515e-09 4.99999997 5.41884515e-09 4.99999997 5.51884515e-09 4.99999997 5.61884515e-09 4.99999997 5.71884515e-09 4.99999997 5.81884515e-09 4.99999997 5.91884515e-09 4.99999997
+ 6.01884515e-09 4.99999997 6.11884515e-09 4.99999997 6.21884515e-09 4.99999997 6.31884515e-09 4.99999997 6.41884515e-09 4.99999997 6.51884515e-09 4.99999997 6.61884515e-09 4.99999997 6.71884515e-09 4.99999997
+ 6.81884515e-09 4.99999997 6.91884515e-09 4.99999997 7.01884515e-09 4.99999997 7.11884515e-09 4.99999997 7.21884515e-09 4.99999997 7.31884515e-09 4.99999997 7.41884515e-09 4.99999997 7.51884515e-09 4.99999997
+ 7.61884515e-09 4.99999997 7.71884515e-09 4.99999997 7.81884515e-09 4.99999997 7.91884515e-09 4.99999997 8.01884515e-09 4.99999997 8.11884515e-09 4.99999997 8.21884515e-09 4.99999997 8.31884515e-09 4.99999997
+ 8.41884515e-09 4.99999997 8.51884515e-09 4.99999997 8.61884515e-09 4.99999997 8.71884515e-09 4.99999997 8.81884515e-09 4.99999997 8.91884515e-09 4.99999997 9.01884515e-09 4.99999997 9.11884515e-09 4.99999997
+ 9.21884515e-09 4.99999997 9.31884515e-09 4.99999997 9.41884515e-09 4.99999997 9.51884515e-09 4.99999997 9.61884515e-09 4.99999997 9.71884515e-09 4.99999997 9.81884515e-09 4.99999997 9.91884515e-09 4.99999997
+ 1.00188451e-08 4.99999997 1.01188451e-08 4.99999997 1.02188451e-08 4.99999997 1.03188451e-08 4.99999997 1.04188451e-08 4.99999997 1.05188451e-08 4.99999997 1.06188451e-08 4.99999997 1.07188451e-08 4.99999997
+ 1.08188451e-08 4.99999997 1.09188451e-08 4.99999997 1.10188451e-08 4.99999997 1.11188451e-08 4.99999997 1.12188451e-08 4.99999997 1.13188451e-08 4.99999997 1.14188451e-08 4.99999997 1.15188451e-08 4.99999997
+ 1.16188451e-08 4.99999997 1.17188451e-08 4.99999997 1.18188451e-08 4.99999997 1.19188451e-08 4.99999997 1.20188451e-08 4.99999997 1.21188451e-08 4.99999997 1.22188451e-08 4.99999997 1.23188451e-08 4.99999997
+ 1.24188451e-08 4.99999997 1.25188451e-08 4.99999997 1.26188451e-08 4.99999997 1.27188451e-08 4.99999997 1.28188451e-08 4.99999997 1.29188451e-08 4.99999997 1.30188451e-08 4.99999997 1.31188451e-08 4.99999997
+ 1.32188451e-08 4.99999997 1.33188451e-08 4.99999997 1.34188451e-08 4.99999997 1.35188451e-08 4.99999997 1.36188451e-08 4.99999997 1.37188451e-08 4.99999997 1.38188451e-08 4.99999997 1.39188451e-08 4.99999997
+ 1.40188451e-08 4.99999997 1.41188451e-08 4.99999997 1.42188451e-08 4.99999997 1.43188451e-08 4.99999997 1.44188451e-08 4.99999997 1.45188451e-08 4.99999997 1.46188451e-08 4.99999997 1.47188451e-08 4.99999997
+ 1.48188451e-08 4.99999997 1.49188451e-08 4.99999997 1.50188451e-08 4.99999997 1.51188451e-08 4.99999997 1.52188451e-08 4.99999997 1.53188451e-08 4.99999997 1.54188451e-08 4.99999997 1.55188451e-08 4.99999997
+ 1.56188451e-08 4.99999997 1.57188451e-08 4.99999997 1.58188451e-08 4.99999997 1.59188451e-08 4.99999997 1.60188451e-08 4.99999997 1.61188451e-08 4.99999997 1.62188451e-08 4.99999997 1.63188451e-08 4.99999997
+ 1.64188451e-08 4.99999997 1.65188451e-08 4.99999997 1.66188451e-08 4.99999997 1.67188451e-08 4.99999997 1.68188451e-08 4.99999997 1.69188451e-08 4.99999997 1.70188451e-08 4.99999997 1.71188451e-08 4.99999997
+ 1.72188451e-08 4.99999997 1.73188451e-08 4.99999997 1.74188451e-08 4.99999997 1.75188451e-08 4.99999997 1.76188451e-08 4.99999997 1.77188451e-08 4.99999997 1.78188451e-08 4.99999997 1.79188451e-08 4.99999997
+ 1.80188451e-08 4.99999997 1.81188451e-08 4.99999997 1.82188451e-08 4.99999997 1.83188451e-08 4.99999997 1.84188451e-08 4.99999997 1.85188451e-08 4.99999997 1.86188451e-08 4.99999997 1.87188451e-08 4.99999997
+ 1.88188451e-08 4.99999997 1.89188451e-08 4.99999997 1.90188451e-08 4.99999997 1.91188451e-08 4.99999997 1.92188451e-08 4.99999997 1.93188451e-08 4.99999997 1.94188451e-08 4.99999997 1.95188451e-08 4.99999997
+ 1.96188451e-08 4.99999997 1.97188451e-08 4.99999997 1.98188451e-08 4.99999997 1.99188451e-08 4.99999997 2e-08 4.99999997 2.001e-08 4.99999997 2.003e-08 4.99999997 2.007e-08 4.99999997
+ 2.01e-08 4.99999997 2.0108e-08 4.99999998 2.0124e-08 4.99999997 2.0156e-08 4.99999996 2.02150599e-08 4.99999999 2.02823902e-08 4.99999997 2.03483061e-08 4.99999995 2.04483061e-08 5.00000001
+ 2.05483061e-08 4.99999993 2.06483061e-08 5.00000003 2.07483061e-08 4.99999991 2.08483061e-08 5.00000004 2.09483061e-08 4.9999999 2.10483061e-08 5.00000004 2.11483061e-08 4.99999991 2.12483061e-08 5.00000003
+ 2.13483061e-08 4.99999992 2.14483061e-08 5.00000001 2.15483061e-08 4.99999994 2.16483061e-08 4.99999999 2.17483061e-08 4.99999996 2.18483061e-08 4.99999998 2.19483061e-08 4.99999997 2.20483061e-08 4.99999997
+ 2.21483061e-08 4.99999998 2.22483061e-08 4.99999997 2.23483061e-08 4.99999998 2.24483061e-08 4.99999996 2.25483061e-08 4.99999998 2.26483061e-08 4.99999996 2.27483061e-08 4.99999998 2.28483061e-08 4.99999996
+ 2.29483061e-08 4.99999998 2.30483061e-08 4.99999996 2.31483061e-08 4.99999998 2.32483061e-08 4.99999997 2.33483061e-08 4.99999998 2.34483061e-08 4.99999997 2.35483061e-08 4.99999998 2.36483061e-08 4.99999997
+ 2.37483061e-08 4.99999998 2.38483061e-08 4.99999997 2.39483061e-08 4.99999998 2.40483061e-08 4.99999997 2.41483061e-08 4.99999998 2.42483061e-08 4.99999997 2.43483061e-08 4.99999997 2.44483061e-08 4.99999997
+ 2.45483061e-08 4.99999997 2.46483061e-08 4.99999997 2.47483061e-08 4.99999997 2.48483061e-08 4.99999997 2.49483061e-08 4.99999997 2.50483061e-08 4.99999997 2.51483061e-08 4.99999997 2.52483061e-08 4.99999997
+ 2.53483061e-08 4.99999997 2.54483061e-08 4.99999997 2.55483061e-08 4.99999997 2.56483061e-08 4.99999997 2.57483061e-08 4.99999997 2.58483061e-08 4.99999997 2.59483061e-08 4.99999997 2.60483061e-08 4.99999997
+ 2.61483061e-08 4.99999997 2.62483061e-08 4.99999997 2.63483061e-08 4.99999997 2.64483061e-08 4.99999997 2.65483061e-08 4.99999997 2.66483061e-08 4.99999997 2.67483061e-08 4.99999997 2.68483061e-08 4.99999997
+ 2.69483061e-08 4.99999997 2.70483061e-08 4.99999997 2.71483061e-08 4.99999997 2.72483061e-08 4.99999997 2.73483061e-08 4.99999997 2.74483061e-08 4.99999997 2.75483061e-08 4.99999997 2.76483061e-08 4.99999997
+ 2.77483061e-08 4.99999997 2.78483061e-08 4.99999997 2.79483061e-08 4.99999997 2.80483061e-08 4.99999997 2.81483061e-08 4.99999997 2.82483061e-08 4.99999997 2.83483061e-08 4.99999997 2.84483061e-08 4.99999997
+ 2.85483061e-08 4.99999997 2.86483061e-08 4.99999997 2.87483061e-08 4.99999997 2.88483061e-08 4.99999997 2.89483061e-08 4.99999997 2.90483061e-08 4.99999997 2.91483061e-08 4.99999997 2.92483061e-08 4.99999997
+ 2.93483061e-08 4.99999997 2.94483061e-08 4.99999997 2.95483061e-08 4.99999997 2.96483061e-08 4.99999997 2.97483061e-08 4.99999997 2.98483061e-08 4.99999997 2.99483061e-08 4.99999997 3.00483061e-08 4.99999997
+ 3.01483061e-08 4.99999997 3.02483061e-08 4.99999997 3.03483061e-08 4.99999997 3.04483061e-08 4.99999997 3.05483061e-08 4.99999997 3.06483061e-08 4.99999997 3.07483061e-08 4.99999997 3.08483061e-08 4.99999997
+ 3.09483061e-08 4.99999997 3.10483061e-08 4.99999997 3.11483061e-08 4.99999997 3.12483061e-08 4.99999997 3.13483061e-08 4.99999997 3.14483061e-08 4.99999997 3.15483061e-08 4.99999997 3.16483061e-08 4.99999997
+ 3.17483061e-08 4.99999997 3.18483061e-08 4.99999997 3.19483061e-08 4.99999997 3.20483061e-08 4.99999997 3.21483061e-08 4.99999997 3.22483061e-08 4.99999997 3.23483061e-08 4.99999997 3.24483061e-08 4.99999997
+ 3.25483061e-08 4.99999997 3.26483061e-08 4.99999997 3.27483061e-08 4.99999997 3.28483061e-08 4.99999997 3.29483061e-08 4.99999997 3.30483061e-08 4.99999997 3.31483061e-08 4.99999997 3.32483061e-08 4.99999997
+ 3.33483061e-08 4.99999997 3.34483061e-08 4.99999997 3.35483061e-08 4.99999997 3.36483061e-08 4.99999997 3.37483061e-08 4.99999997 3.38483061e-08 4.99999997 3.39483061e-08 4.99999997 3.40483061e-08 4.99999997
+ 3.41483061e-08 4.99999997 3.42483061e-08 4.99999997 3.43483061e-08 4.99999997 3.44483061e-08 4.99999997 3.45483061e-08 4.99999997 3.46483061e-08 4.99999997 3.47483061e-08 4.99999997 3.48483061e-08 4.99999997
+ 3.49483061e-08 4.99999997 3.50483061e-08 4.99999997 3.51483061e-08 4.99999997 3.52483061e-08 4.99999997 3.53483061e-08 4.99999997 3.54483061e-08 4.99999997 3.55483061e-08 4.99999997 3.56483061e-08 4.99999997
+ 3.57483061e-08 4.99999997 3.58483061e-08 4.99999997 3.59483061e-08 4.99999997 3.60483061e-08 4.99999997 3.61483061e-08 4.99999997 3.62483061e-08 4.99999997 3.63483061e-08 4.99999997 3.64483061e-08 4.99999997
+ 3.65483061e-08 4.99999997 3.66483061e-08 4.99999997 3.67483061e-08 4.99999997 3.68483061e-08 4.99999997 3.69483061e-08 4.99999997 3.70483061e-08 4.99999997 3.71483061e-08 4.99999997 3.72483061e-08 4.99999997
+ 3.73483061e-08 4.99999997 3.74483061e-08 4.99999997 3.75483061e-08 4.99999997 3.76483061e-08 4.99999997 3.77483061e-08 4.99999997 3.78483061e-08 4.99999997 3.79483061e-08 4.99999997 3.80483061e-08 4.99999997
+ 3.81483061e-08 4.99999997 3.82483061e-08 4.99999997 3.83483061e-08 4.99999997 3.84483061e-08 4.99999997 3.85483061e-08 4.99999997 3.86483061e-08 4.99999997 3.87483061e-08 4.99999997 3.88483061e-08 4.99999997
+ 3.89483061e-08 4.99999997 3.90483061e-08 4.99999997 3.91483061e-08 4.99999997 3.92483061e-08 4.99999997 3.93483061e-08 4.99999997 3.94483061e-08 4.99999997 3.95483061e-08 4.99999997 3.96483061e-08 4.99999997
+ 3.97483061e-08 4.99999997 3.98483061e-08 4.99999997 3.99483061e-08 4.99999997 4.00483061e-08 4.99999997 4.01483061e-08 4.99999997 4.02483061e-08 4.99999997 4.03483061e-08 4.99999997 4.04483061e-08 4.99999997
+ 4.05483061e-08 4.99999997 4.06483061e-08 4.99999997 4.07483061e-08 4.99999997 4.08483061e-08 4.99999997 4.09483061e-08 4.99999997 4.10483061e-08 4.99999997 4.11483061e-08 4.99999997 4.12483061e-08 4.99999997
+ 4.13483061e-08 4.99999997 4.14483061e-08 4.99999997 4.15483061e-08 4.99999997 4.16483061e-08 4.99999997 4.17483061e-08 4.99999997 4.18483061e-08 4.99999997 4.19483061e-08 4.99999997 4.20483061e-08 4.99999997
+ 4.21483061e-08 4.99999997 4.22483061e-08 4.99999997 4.23483061e-08 4.99999997 4.24483061e-08 4.99999997 4.25483061e-08 4.99999997 4.26483061e-08 4.99999997 4.27483061e-08 4.99999997 4.28483061e-08 4.99999997
+ 4.29483061e-08 4.99999997 4.30483061e-08 4.99999997 4.31483061e-08 4.99999997 4.32483061e-08 4.99999997 4.33483061e-08 4.99999997 4.34483061e-08 4.99999997 4.35483061e-08 4.99999997 4.36483061e-08 4.99999997
+ 4.37483061e-08 4.99999997 4.38483061e-08 4.99999997 4.39483061e-08 4.99999997 4.40483061e-08 4.99999997 4.41483061e-08 4.99999997 4.42483061e-08 4.99999997 4.43483061e-08 4.99999997 4.44483061e-08 4.99999997
+ 4.45483061e-08 4.99999997 4.46483061e-08 4.99999997 4.47483061e-08 4.99999997 4.48483061e-08 4.99999997 4.49483061e-08 4.99999997 4.50483061e-08 4.99999997 4.51483061e-08 4.99999997 4.52483061e-08 4.99999997
+ 4.53483061e-08 4.99999997 4.54483061e-08 4.99999997 4.55483061e-08 4.99999997 4.56483061e-08 4.99999997 4.57483061e-08 4.99999997 4.58483061e-08 4.99999997 4.59483061e-08 4.99999997 4.60483061e-08 4.99999997
+ 4.61483061e-08 4.99999997 4.62483061e-08 4.99999997 4.63483061e-08 4.99999997 4.64483061e-08 4.99999997 4.65483061e-08 4.99999997 4.66483061e-08 4.99999997 4.67483061e-08 4.99999997 4.68483061e-08 4.99999997
+ 4.69483061e-08 4.99999997 4.70483061e-08 4.99999997 4.71483061e-08 4.99999997 4.72483061e-08 4.99999997 4.73483061e-08 4.99999997 4.74483061e-08 4.99999997 4.75483061e-08 4.99999997 4.76483061e-08 4.99999997
+ 4.77483061e-08 4.99999997 4.78483061e-08 4.99999997 4.79483061e-08 4.99999997 4.80483061e-08 4.99999997 4.81483061e-08 4.99999997 4.82483061e-08 4.99999997 4.83483061e-08 4.99999997 4.84483061e-08 4.99999997
+ 4.85483061e-08 4.99999997 4.86483061e-08 4.99999997 4.87483061e-08 4.99999997 4.88483061e-08 4.99999997 4.89483061e-08 4.99999997 4.90483061e-08 4.99999997 4.91483061e-08 4.99999997 4.92483061e-08 4.99999997
+ 4.93483061e-08 4.99999997 4.94483061e-08 4.99999997 4.95483061e-08 4.99999997 4.96483061e-08 4.99999997 4.97483061e-08 4.99999997 4.98483061e-08 4.99999997 4.99483061e-08 4.99999997 5.00483061e-08 4.99999997
+ 5.01483061e-08 4.99999997 5.02483061e-08 4.99999997 5.03483061e-08 4.99999997 5.04483061e-08 4.99999997 5.05483061e-08 4.99999997 5.06483061e-08 4.99999997 5.07483061e-08 4.99999997 5.08483061e-08 4.99999997
+ 5.09483061e-08 4.99999997 5.1e-08 4.99999997 5.101e-08 4.99999997 5.103e-08 4.99999998 5.107e-08 4.99999996 5.115e-08 4.99999998 5.125e-08 4.99999997 5.135e-08 4.99999997
+ 5.145e-08 4.99999998 5.155e-08 4.99999996 5.165e-08 4.99999998 5.175e-08 4.99999996 5.185e-08 4.99999999 5.19308282e-08 5.00006476 5.2e-08 4.99916064 5.20086083e-08 4.99761639
+ 5.2025825e-08 4.99311196 5.20602584e-08 5.01027311 5.21061808e-08 5.09906218 5.21500808e-08 4.21229454 5.21980262e-08 0.290284903 5.22553803e-08 -0.0554592023 5.23120186e-08 0.0719468597 5.24042316e-08 -0.0579815953
+ 5.25042316e-08 0.0528904133 5.26042316e-08 -0.0475729854 5.27042316e-08 0.0435757158 5.28042316e-08 -0.0393284178 5.29042316e-08 0.0359989191 5.30042316e-08 -0.0325572549 5.31042316e-08 0.0297863163 5.32042316e-08 -0.0269831353
+ 5.33042316e-08 0.024677895 5.34042316e-08 -0.0223854069 5.35042316e-08 0.0204676265 5.36042316e-08 -0.0185865295 5.37042316e-08 0.0169908361 5.38042316e-08 -0.0154430663 5.39042316e-08 0.0141150741 5.40042316e-08 -0.0128386861
+ 5.41042316e-08 0.0117332242 5.42042316e-08 -0.0106786681 5.43042316e-08 0.00975824024 5.44042316e-08 -0.00888561579 5.45042316e-08 0.00811909449 5.46042316e-08 -0.00739609091 5.47042316e-08 0.00675762723 5.48042316e-08 -0.00615795518
+ 5.49042316e-08 0.00562607399 5.50042316e-08 -0.00512825797 5.51042316e-08 0.00468510952 5.52042316e-08 -0.00427154749 5.53042316e-08 0.00390228875 5.54042316e-08 -0.00355851286 5.55042316e-08 0.00325079606 5.56042316e-08 -0.00296488651
+ 5.57042316e-08 0.002708436 5.58042316e-08 -0.0024705529 5.59042316e-08 0.00225681481 5.60042316e-08 -0.00205882186 5.61042316e-08 0.00188067375 5.62042316e-08 -0.00171583399 5.63042316e-08 0.00156734401 5.64042316e-08 -0.00143007279
+ 5.65042316e-08 0.00130629977 5.66042316e-08 -0.00119196316 5.67042316e-08 0.00108879052 5.68042316e-08 -0.000993540456 5.69042316e-08 0.000907538165 5.70042316e-08 -0.000828177003 5.71042316e-08 0.000756486788 5.72042316e-08 -0.000690355922
+ 5.73042316e-08 0.000630595752 5.74042316e-08 -0.00057548372 5.75042316e-08 0.000525668321 5.76042316e-08 -0.000479734899 5.77042316e-08 0.000438209567 5.78042316e-08 -0.000399922963 5.79042316e-08 0.000365308462 5.80042316e-08 -0.000333393279
+ 5.81042316e-08 0.000304539934 5.82042316e-08 -0.000277934025 5.83042316e-08 0.000253883483 5.84042316e-08 -0.000231702133 5.85042316e-08 0.000211655506 5.86042316e-08 -0.000193161676 5.87042316e-08 0.00017645299 5.88042316e-08 -0.000161032592
+ 5.89042316e-08 0.000147106669 5.90042316e-08 -0.000134248002 5.91042316e-08 0.000122642012 5.92042316e-08 -0.000111918653 5.93042316e-08 0.000102246759 5.94042316e-08 -9.33033252e-05 5.95042316e-08 8.52438625e-05 5.96042316e-08 -7.77841591e-05
+ 5.97042316e-08 7.10689667e-05 5.98042316e-08 -6.48461156e-05 5.99042316e-08 5.92516326e-05 6.00042316e-08 -5.40598536e-05 6.01042316e-08 4.93997007e-05 6.02042316e-08 -4.50674637e-05 6.03042316e-08 4.1186259e-05 6.04042316e-08 -3.75705792e-05
+ 6.05042316e-08 3.43387822e-05 6.06042316e-08 -3.13204669e-05 6.07042316e-08 2.86300808e-05 6.08042316e-08 -2.61097684e-05 6.09042316e-08 2.38707568e-05 6.10042316e-08 -2.17656162e-05 6.11042316e-08 1.99029161e-05 6.12042316e-08 -1.81438953e-05
+ 6.13042316e-08 1.65949269e-05 6.14042316e-08 -1.51244604e-05 6.15042316e-08 1.38370509e-05 6.16042316e-08 -1.26071484e-05 6.17042316e-08 1.15378015e-05 6.18042316e-08 -1.05084548e-05 6.19042316e-08 9.62090752e-06 6.20042316e-08 -8.75876286e-06
+ 6.21042316e-08 8.02278269e-06 6.22042316e-08 -7.30003357e-06 6.23042316e-08 6.69041567e-06 6.24042316e-08 -6.08388026e-06 6.25042316e-08 5.57961126e-06 6.26042316e-08 -5.06996313e-06 6.27042316e-08 4.65352414e-06 6.28042316e-08 -4.22465101e-06
+ 6.29042316e-08 3.88143646e-06 6.30042316e-08 -3.51990563e-06 6.31042316e-08 3.2377388e-06 6.32042316e-08 -2.93235147e-06 6.33042316e-08 2.70108059e-06 6.34042316e-08 -2.44250035e-06 6.35042316e-08 2.25366182e-06 6.36042316e-08 -2.03410493e-06
+ 6.37042316e-08 1.88064262e-06 6.38042316e-08 -1.69361976e-06 6.39042316e-08 1.56965096e-06 6.40042316e-08 -1.40079515e-06 6.41042316e-08 1.32022173e-06 6.42042316e-08 -1.16495133e-06 6.43042316e-08 1.10221056e-06 6.44042316e-08 -9.6884516e-07
+ 6.45042316e-08 9.20524819e-07 6.46042316e-08 -8.05378027e-07 6.47042316e-08 7.69073313e-07 6.48042316e-08 -6.69112959e-07 6.49042316e-08 6.42824092e-07 6.50042316e-08 -5.5552303e-07 6.51042316e-08 5.37583129e-07 6.52042316e-08 -4.60834674e-07
+ 6.53042316e-08 4.49854039e-07 6.54042316e-08 -3.81902022e-07 6.55042316e-08 3.76722702e-07 6.56042316e-08 -3.16103666e-07 6.57042316e-08 3.15760347e-07 6.58042316e-08 -2.61254034e-07 6.59042316e-08 2.64941902e-07 6.60042316e-08 -2.15531327e-07
+ 6.61042316e-08 2.22579744e-07 6.62042316e-08 -1.77426895e-07 6.63042316e-08 1.87286706e-07 6.64042316e-08 -1.45681881e-07 6.65042316e-08 1.57883818e-07 6.66042316e-08 -1.19234761e-07 6.67042316e-08 1.33387831e-07 6.68042316e-08 -9.72011708e-08
+ 6.69042316e-08 1.12979676e-07 6.70042316e-08 -7.88444182e-08 6.71042316e-08 9.5977075e-08 6.72042316e-08 -6.35509314e-08 6.73042316e-08 8.18118485e-08 6.74042316e-08 -5.07711936e-08 6.75042316e-08 6.99714195e-08 6.76042316e-08 -4.01609191e-08
+ 6.77042316e-08 6.01479495e-08 6.78042316e-08 -3.13252177e-08 6.79042316e-08 5.19642415e-08 6.80042316e-08 -2.39641178e-08 6.81042316e-08 4.51463234e-08 6.82042316e-08 -1.78315414e-08 6.83042316e-08 3.94660711e-08 6.84042316e-08 -1.27218748e-08
+ 6.85042316e-08 3.47333458e-08 6.86042316e-08 -8.46503329e-09 6.87042316e-08 3.07907601e-08 6.88042316e-08 -4.9188682e-09 6.89042316e-08 2.75063625e-08 6.90042316e-08 -1.96469058e-09 6.91042316e-08 2.47702336e-08 6.92042316e-08 4.96360592e-10
+ 6.93042316e-08 2.24973263e-08 6.94042316e-08 2.54107269e-09 6.95042316e-08 2.06302864e-08 6.96042316e-08 4.22166857e-09 6.97042316e-08 1.90955815e-08 6.98042316e-08 5.60316635e-09 6.99042316e-08 1.78339741e-08 7.00042316e-08 6.73885944e-09
+ 7.01042316e-08 1.67968134e-08 7.02042316e-08 7.67252992e-09 7.03042316e-08 1.59441272e-08 7.04042316e-08 8.44015105e-09 7.05042316e-08 1.5143766e-08 7.06042316e-08 9.05741654e-09 7.07042316e-08 1.45796351e-08 7.08042316e-08 9.5695612e-09
+ 7.09042316e-08 1.41150197e-08 7.10042316e-08 9.99102767e-09 7.11042316e-08 1.37326954e-08 7.12042316e-08 1.03378474e-08 7.13042316e-08 1.3418081e-08 7.14042316e-08 1.06232494e-08 7.15042316e-08 1.31591765e-08 7.16042316e-08 1.08581189e-08
+ 7.17042316e-08 1.29461085e-08 7.18042316e-08 1.10514114e-08 7.19042316e-08 1.27707539e-08 7.20042316e-08 1.12104946e-08 7.21042316e-08 1.26264306e-08 7.22042316e-08 1.13414295e-08 7.23042316e-08 1.25076402e-08 7.24042316e-08 1.14492033e-08
+ 7.25042316e-08 1.24098599e-08 7.26042316e-08 1.15379184e-08 7.27042316e-08 1.23293677e-08 7.28042316e-08 1.16109512e-08 7.29042316e-08 1.22631022e-08 7.30042316e-08 1.16710779e-08 7.31042316e-08 1.22085441e-08 7.32042316e-08 1.17205841e-08
+ 7.33042316e-08 1.21636207e-08 7.34042316e-08 1.17613498e-08 7.35042316e-08 1.21266268e-08 7.36042316e-08 1.17949218e-08 7.37042316e-08 1.20961591e-08 7.38042316e-08 1.18225734e-08 7.39042316e-08 1.2071063e-08 7.40042316e-08 1.18453512e-08
+ 7.41042316e-08 1.20503885e-08 7.42042316e-08 1.18641169e-08 7.43042316e-08 1.2033354e-08 7.44042316e-08 1.18795805e-08 7.45042316e-08 1.20193162e-08 7.46042316e-08 1.18923249e-08 7.47042316e-08 1.20077459e-08 7.48042316e-08 1.19028301e-08
+ 7.49042316e-08 1.1998207e-08 7.50042316e-08 1.1911492e-08 7.51042316e-08 1.19903412e-08 7.52042316e-08 1.19186351e-08 7.53042316e-08 1.19838536e-08 7.54042316e-08 1.1924528e-08 7.55042316e-08 1.19785007e-08 7.56042316e-08 1.19293902e-08
+ 7.57042316e-08 1.19740839e-08 7.58042316e-08 1.19334033e-08 7.59042316e-08 1.19704374e-08 7.60042316e-08 1.19367169e-08 7.61042316e-08 1.19674258e-08 7.62042316e-08 1.19394544e-08 7.63042316e-08 1.19649375e-08 7.64042316e-08 1.19417163e-08
+ 7.65042316e-08 1.1962881e-08 7.66042316e-08 1.19435867e-08 7.67042316e-08 1.19611798e-08 7.68042316e-08 1.19451338e-08 7.69042316e-08 1.19597724e-08 7.70042316e-08 1.1946414e-08 7.71042316e-08 1.19586075e-08 7.72042316e-08 1.19474741e-08
+ 7.73042316e-08 1.19576425e-08 7.74042316e-08 1.19483529e-08 7.75042316e-08 1.19568423e-08 7.76042316e-08 1.19490814e-08 7.77042316e-08 1.19561787e-08 7.78042316e-08 1.19496862e-08 7.79042316e-08 1.19556277e-08 7.80042316e-08 1.19501884e-08
+ 7.81042316e-08 1.19551702e-08 7.82042316e-08 1.19506057e-08 7.83042316e-08 1.19547894e-08 7.84042316e-08 1.1950953e-08 7.85042316e-08 1.19544723e-08 7.86042316e-08 1.19512423e-08 7.87042316e-08 1.19542082e-08 7.88042316e-08 1.19514836e-08
+ 7.89042316e-08 1.19539879e-08 7.90042316e-08 1.19516851e-08 7.91042316e-08 1.19538036e-08 7.92042316e-08 1.19518535e-08 7.93042316e-08 1.19536496e-08 7.94042316e-08 1.19519949e-08 7.95042316e-08 1.19535202e-08 7.96042316e-08 1.1952113e-08
+ 7.97042316e-08 1.19534117e-08 7.98042316e-08 1.19522124e-08 7.99042316e-08 1.19533209e-08 8.00042316e-08 1.19522957e-08 8.01042316e-08 1.19532438e-08 8.02042316e-08 1.19523665e-08 8.03042316e-08 1.1953179e-08 8.04042316e-08 1.19524259e-08
+ 8.05042316e-08 1.19531247e-08 8.06042316e-08 1.19524759e-08 8.07042316e-08 1.19530783e-08 8.08042316e-08 1.19525188e-08 8.09042316e-08 1.19530389e-08 8.10042316e-08 1.1952555e-08 8.11042316e-08 1.19530056e-08 8.12042316e-08 1.1952586e-08
+ 8.13042316e-08 1.19529771e-08 8.14042316e-08 1.19526124e-08 8.15042316e-08 1.19529523e-08 8.16042316e-08 1.19526352e-08 8.17042316e-08 1.19529313e-08 8.18042316e-08 1.19526544e-08 8.19042316e-08 1.19529137e-08 8.20042316e-08 1.19526709e-08
+ 8.21042316e-08 1.19528983e-08 8.22042316e-08 1.19526853e-08 8.23042316e-08 1.19528848e-08 8.24042316e-08 1.19526976e-08 8.25042316e-08 1.19528734e-08 8.26042316e-08 1.19527083e-08 8.27042316e-08 1.19528634e-08 8.28042316e-08 1.19527175e-08
+ 8.29042316e-08 1.19528546e-08 8.30042316e-08 1.19527257e-08 8.31042316e-08 1.19528473e-08 8.32042316e-08 1.19527327e-08 8.33042316e-08 1.19528406e-08 8.34042316e-08 1.19527392e-08 8.35042316e-08 1.19528347e-08 8.36042316e-08 1.19527446e-08
+ 8.37042316e-08 1.19528298e-08 8.38042316e-08 1.19527492e-08 8.39042316e-08 1.1952825e-08 8.40042316e-08 1.19527536e-08 8.41042316e-08 1.19528211e-08 8.42042316e-08 1.19527572e-08 8.43042316e-08 1.19528178e-08 8.44042316e-08 1.19527606e-08
+ 8.45042316e-08 1.19528146e-08 8.46042316e-08 1.19527634e-08 8.47042316e-08 1.19528118e-08 8.48042316e-08 1.19527659e-08 8.49042316e-08 1.19528095e-08 8.50042316e-08 1.19527683e-08 8.51042316e-08 1.19528072e-08 8.52042316e-08 1.19527702e-08
+ 8.53042316e-08 1.19528053e-08 8.54042316e-08 1.1952772e-08 8.55042316e-08 1.19528037e-08 8.56042316e-08 1.19527737e-08 8.57042316e-08 1.1952802e-08 8.58042316e-08 1.19527752e-08 8.59042316e-08 1.19528006e-08 8.60042316e-08 1.19527765e-08
+ 8.61042316e-08 1.19527997e-08 8.62042316e-08 1.19527775e-08 8.63042316e-08 1.19527986e-08 8.64042316e-08 1.19527785e-08 8.65042316e-08 1.19527975e-08 8.66042316e-08 1.19527796e-08 8.67042316e-08 1.19527964e-08 8.68042316e-08 1.19527805e-08
+ 8.69042316e-08 1.19527956e-08 8.70042316e-08 1.19527813e-08 8.71042316e-08 1.19527947e-08 8.72042316e-08 1.1952782e-08 8.73042316e-08 1.19527943e-08 8.74042316e-08 1.19527827e-08 8.75042316e-08 1.19527936e-08 8.76042316e-08 1.1952783e-08
+ 8.77042316e-08 1.19527933e-08 8.78042316e-08 1.19527836e-08 8.79042316e-08 1.19527929e-08 8.80042316e-08 1.19527841e-08 8.81042316e-08 1.19527925e-08 8.82042316e-08 1.19527844e-08 8.83042316e-08 1.19527919e-08 8.84042316e-08 1.19527848e-08
+ 8.85042316e-08 1.19527918e-08 8.86042316e-08 1.19527851e-08 8.87042316e-08 1.19527915e-08 8.88042316e-08 1.19527855e-08 8.89042316e-08 1.19527911e-08 8.90042316e-08 1.19527858e-08 8.91042316e-08 1.19527907e-08 8.92042316e-08 1.19527862e-08
+ 8.93042316e-08 1.19527902e-08 8.94042316e-08 1.19527863e-08 8.95042316e-08 1.19527903e-08 8.96042316e-08 1.19527865e-08 8.97042316e-08 1.195279e-08 8.98042316e-08 1.19527868e-08 8.99042316e-08 1.19527901e-08 9.00042316e-08 1.19527867e-08
+ 9.01042316e-08 1.19527897e-08 9.02042316e-08 1.1952787e-08 9.03042316e-08 1.19527894e-08 9.04042316e-08 1.19527871e-08 9.05042316e-08 1.19527895e-08 9.06042316e-08 1.19527871e-08 9.07042316e-08 1.19527896e-08 9.08042316e-08 1.19527872e-08
+ 9.09042316e-08 1.19527896e-08 9.10042316e-08 1.19527872e-08 9.11042316e-08 1.19527895e-08 9.12042316e-08 1.19527873e-08 9.13042316e-08 1.19527894e-08 9.14042316e-08 1.19527873e-08 9.15042316e-08 1.19527893e-08 9.16042316e-08 1.19527873e-08
+ 9.17042316e-08 1.19527896e-08 9.18042316e-08 1.19527873e-08 9.19042316e-08 1.19527891e-08 9.20042316e-08 1.19527874e-08 9.21042316e-08 1.19527891e-08 9.22042316e-08 1.19527875e-08 9.23042316e-08 1.19527891e-08 9.24042316e-08 1.19527874e-08
+ 9.25042316e-08 1.19527891e-08 9.26042316e-08 1.19527875e-08 9.27042316e-08 1.19527891e-08 9.28042316e-08 1.19527875e-08 9.29042316e-08 1.19527892e-08 9.30042316e-08 1.19527877e-08 9.31042316e-08 1.1952789e-08 9.32042316e-08 1.19527878e-08
+ 9.33042316e-08 1.19527891e-08 9.34042316e-08 1.19527878e-08 9.35042316e-08 1.1952789e-08 9.36042316e-08 1.19527879e-08 9.37042316e-08 1.1952789e-08 9.38042316e-08 1.19527878e-08 9.39042316e-08 1.19527889e-08 9.40042316e-08 1.19527879e-08
+ 9.41042316e-08 1.19527889e-08 9.42042316e-08 1.19527879e-08 9.43042316e-08 1.19527888e-08 9.44042316e-08 1.1952788e-08 9.45042316e-08 1.19527888e-08 9.46042316e-08 1.1952788e-08 9.47042316e-08 1.19527887e-08 9.48042316e-08 1.19527881e-08
+ 9.49042316e-08 1.19527888e-08 9.50042316e-08 1.19527881e-08 9.51042316e-08 1.19527887e-08 9.52042316e-08 1.19527882e-08 9.53042316e-08 1.19527887e-08 9.54042316e-08 1.19527881e-08 9.55042316e-08 1.19527886e-08 9.56042316e-08 1.19527883e-08
+ 9.57042316e-08 1.19527885e-08 9.58042316e-08 1.19527882e-08 9.59042316e-08 1.19527885e-08 9.60042316e-08 1.19527882e-08 9.61042316e-08 1.19527885e-08 9.62042316e-08 1.19527882e-08 9.63042316e-08 1.19527885e-08 9.64042316e-08 1.19527883e-08
+ 9.65042316e-08 1.19527884e-08 9.66042316e-08 1.19527883e-08 9.67042316e-08 1.19527885e-08 9.68042316e-08 1.19527883e-08 9.69042316e-08 1.19527884e-08 9.70042316e-08 1.19527883e-08 9.71042316e-08 1.19527885e-08 9.72042316e-08 1.19527883e-08
+ 9.73042316e-08 1.19527885e-08 9.74042316e-08 1.19527883e-08 9.75042316e-08 1.19527885e-08 9.76042316e-08 1.19527883e-08 9.77042316e-08 1.19527885e-08 9.78042316e-08 1.19527883e-08 9.79042316e-08 1.19527885e-08 9.80042316e-08 1.19527883e-08
+ 9.81042316e-08 1.19527885e-08 9.82042316e-08 1.19527883e-08 9.83042316e-08 1.19527885e-08 9.84042316e-08 1.19527883e-08 9.85042316e-08 1.19527885e-08 9.86042316e-08 1.19527883e-08 9.87042316e-08 1.19527885e-08 9.88042316e-08 1.19527883e-08
+ 9.89042316e-08 1.19527885e-08 9.90042316e-08 1.19527883e-08 9.91042316e-08 1.19527884e-08 9.92042316e-08 1.19527883e-08 9.93042316e-08 1.19527885e-08 9.94042316e-08 1.19527883e-08 9.95042316e-08 1.19527885e-08 9.96042316e-08 1.19527883e-08
+ 9.97042316e-08 1.19527885e-08 9.98042316e-08 1.19527883e-08 9.99042316e-08 1.19527885e-08 1e-07 1.19527883e-08 1.0001e-07 1.45267509e-08 1.0003e-07 1.23970234e-09 1.0007e-07 2.76375245e-08 1.0015e-07 -4.37848727e-09
+ 1.0025e-07 2.82049085e-08 1.0035e-07 -3.1772773e-09 1.0045e-07 2.52046163e-08 1.0055e-07 2.60784372e-09 1.0065e-07 -4.06484957e-08 1.0075e-07 3.06912285e-06 1.0085e-07 9.51416721e-05 1.00932051e-07 -0.0447831027
+ 1.01e-07 1.97583273 1.01008488e-07 3.09989962 1.01025463e-07 4.14313244 1.01059414e-07 4.88304728 1.0109062e-07 4.97992695 1.0114347e-07 5.00280645 1.01199151e-07 4.99919782 1.01299151e-07 5.00046536
+ 1.01399151e-07 4.99971259 1.01499151e-07 5.00018323 1.01599151e-07 4.99987811 1.01699151e-07 5.00008217 1.01799151e-07 4.99994319 1.01893117e-07 5.00003832 1.01993117e-07 4.99997306 1.02093117e-07 5.00001877
+ 1.02193117e-07 4.99998672 1.02293117e-07 5.00000925 1.02393117e-07 4.99999343 1.02493117e-07 5.00000455 1.02593117e-07 4.99999675 1.02693117e-07 5.00000222 1.02793117e-07 4.9999984 1.02893117e-07 5.00000106
+ 1.02993117e-07 4.99999921 1.03093117e-07 5.0000005 1.03193117e-07 4.99999961 1.03293117e-07 5.00000022 1.03393117e-07 4.9999998 1.03493117e-07 5.00000008 1.03593117e-07 4.9999999 1.03693117e-07 5.00000002
+ 1.03793117e-07 4.99999994 1.03893117e-07 4.99999999 1.03993117e-07 4.99999996 1.04093117e-07 4.99999998 1.04193117e-07 4.99999997 1.04293117e-07 4.99999997 1.04393117e-07 4.99999997 1.04493117e-07 4.99999997
+ 1.04593117e-07 4.99999997 1.04693117e-07 4.99999997 1.04793117e-07 4.99999997 1.04893117e-07 4.99999997 1.04993117e-07 4.99999997 1.05093117e-07 4.99999997 1.05193117e-07 4.99999997 1.05293117e-07 4.99999997
+ 1.05393117e-07 4.99999997 1.05493117e-07 4.99999997 1.05593117e-07 4.99999997 1.05693117e-07 4.99999997 1.05793117e-07 4.99999997 1.05893117e-07 4.99999997 1.05993117e-07 4.99999997 1.06093117e-07 4.99999997
+ 1.06193117e-07 4.99999997 1.06293117e-07 4.99999997 1.06393117e-07 4.99999997 1.06493117e-07 4.99999997 1.06593117e-07 4.99999997 1.06693117e-07 4.99999997 1.06793117e-07 4.99999997 1.06893117e-07 4.99999997
+ 1.06993117e-07 4.99999997 1.07093117e-07 4.99999997 1.07193117e-07 4.99999997 1.07293117e-07 4.99999997 1.07393117e-07 4.99999997 1.07493117e-07 4.99999997 1.07593117e-07 4.99999997 1.07693117e-07 4.99999997
+ 1.07793117e-07 4.99999997 1.07893117e-07 4.99999997 1.07993117e-07 4.99999997 1.08093117e-07 4.99999997 1.08193117e-07 4.99999997 1.08293117e-07 4.99999997 1.08393117e-07 4.99999997 1.08493117e-07 4.99999997
+ 1.08593117e-07 4.99999997 1.08693117e-07 4.99999997 1.08793117e-07 4.99999997 1.08893117e-07 4.99999997 1.08993117e-07 4.99999997 1.09093117e-07 4.99999997 1.09193117e-07 4.99999997 1.09293117e-07 4.99999997
+ 1.09393117e-07 4.99999997 1.09493117e-07 4.99999997 1.09593117e-07 4.99999997 1.09693117e-07 4.99999997 1.09793117e-07 4.99999997 1.09893117e-07 4.99999997 1.09993117e-07 4.99999997 1.10093117e-07 4.99999997
+ 1.10193117e-07 4.99999997 1.10293117e-07 4.99999997 1.10393117e-07 4.99999997 1.10493117e-07 4.99999997 1.10593117e-07 4.99999997 1.10693117e-07 4.99999997 1.10793117e-07 4.99999997 1.10893117e-07 4.99999997
+ 1.10993117e-07 4.99999997 1.11093117e-07 4.99999997 1.11193117e-07 4.99999997 1.11293117e-07 4.99999997 1.11393117e-07 4.99999997 1.11493117e-07 4.99999997 1.11593117e-07 4.99999997 1.11693117e-07 4.99999997
+ 1.11793117e-07 4.99999997 1.11893117e-07 4.99999997 1.11993117e-07 4.99999997 1.12093117e-07 4.99999997 1.12193117e-07 4.99999997 1.12293117e-07 4.99999997 1.12393117e-07 4.99999997 1.12493117e-07 4.99999997
+ 1.12593117e-07 4.99999997 1.12693117e-07 4.99999997 1.12793117e-07 4.99999997 1.12893117e-07 4.99999997 1.12993117e-07 4.99999997 1.13093117e-07 4.99999997 1.13193117e-07 4.99999997 1.13293117e-07 4.99999997
+ 1.13393117e-07 4.99999997 1.13493117e-07 4.99999997 1.13593117e-07 4.99999997 1.13693117e-07 4.99999997 1.13793117e-07 4.99999997 1.13893117e-07 4.99999997 1.13993117e-07 4.99999997 1.14093117e-07 4.99999997
+ 1.14193117e-07 4.99999997 1.14293117e-07 4.99999997 1.14393117e-07 4.99999997 1.14493117e-07 4.99999997 1.14593117e-07 4.99999997 1.14693117e-07 4.99999997 1.14793117e-07 4.99999997 1.14893117e-07 4.99999997
+ 1.14993117e-07 4.99999997 1.15093117e-07 4.99999997 1.15193117e-07 4.99999997 1.15293117e-07 4.99999997 1.15393117e-07 4.99999997 1.15493117e-07 4.99999997 1.15593117e-07 4.99999997 1.15693117e-07 4.99999997
+ 1.15793117e-07 4.99999997 1.15893117e-07 4.99999997 1.15993117e-07 4.99999997 1.16093117e-07 4.99999997 1.16193117e-07 4.99999997 1.16293117e-07 4.99999997 1.16393117e-07 4.99999997 1.16493117e-07 4.99999997
+ 1.16593117e-07 4.99999997 1.16693117e-07 4.99999997 1.16793117e-07 4.99999997 1.16893117e-07 4.99999997 1.16993117e-07 4.99999997 1.17093117e-07 4.99999997 1.17193117e-07 4.99999997 1.17293117e-07 4.99999997
+ 1.17393117e-07 4.99999997 1.17493117e-07 4.99999997 1.17593117e-07 4.99999997 1.17693117e-07 4.99999997 1.17793117e-07 4.99999997 1.17893117e-07 4.99999997 1.17993117e-07 4.99999997 1.18093117e-07 4.99999997
+ 1.18193117e-07 4.99999997 1.18293117e-07 4.99999997 1.18393117e-07 4.99999997 1.18493117e-07 4.99999997 1.18593117e-07 4.99999997 1.18693117e-07 4.99999997 1.18793117e-07 4.99999997 1.18893117e-07 4.99999997
+ 1.18993117e-07 4.99999997 1.19093117e-07 4.99999997 1.19193117e-07 4.99999997 1.19293117e-07 4.99999997 1.19393117e-07 4.99999997 1.19493117e-07 4.99999997 1.19593117e-07 4.99999997 1.19693117e-07 4.99999997
+ 1.19793117e-07 4.99999997 1.19893117e-07 4.99999997 1.19993117e-07 4.99999997 1.20093117e-07 4.99999997 1.20193117e-07 4.99999997 1.20293117e-07 4.99999997 1.20393117e-07 4.99999997 1.20493117e-07 4.99999997
+ 1.20593117e-07 4.99999997 1.20693117e-07 4.99999997 1.20793117e-07 4.99999997 1.20893117e-07 4.99999997 1.20993117e-07 4.99999997 1.21093117e-07 4.99999997 1.21193117e-07 4.99999997 1.21293117e-07 4.99999997
+ 1.21393117e-07 4.99999997 1.21493117e-07 4.99999997 1.21593117e-07 4.99999997 1.21693117e-07 4.99999997 1.21793117e-07 4.99999997 1.21893117e-07 4.99999997 1.21993117e-07 4.99999997 1.22093117e-07 4.99999997
+ 1.22193117e-07 4.99999997 1.22293117e-07 4.99999997 1.22393117e-07 4.99999997 1.22493117e-07 4.99999997 1.22593117e-07 4.99999997 1.22693117e-07 4.99999997 1.22793117e-07 4.99999997 1.22893117e-07 4.99999997
+ 1.22993117e-07 4.99999997 1.23093117e-07 4.99999997 1.23193117e-07 4.99999997 1.23293117e-07 4.99999997 1.23393117e-07 4.99999997 1.23493117e-07 4.99999997 1.23593117e-07 4.99999997 1.23693117e-07 4.99999997
+ 1.23793117e-07 4.99999997 1.23893117e-07 4.99999997 1.23993117e-07 4.99999997 1.24093117e-07 4.99999997 1.24193117e-07 4.99999997 1.24293117e-07 4.99999997 1.24393117e-07 4.99999997 1.24493117e-07 4.99999997
+ 1.24593117e-07 4.99999997 1.24693117e-07 4.99999997 1.24793117e-07 4.99999997 1.24893117e-07 4.99999997 1.24993117e-07 4.99999997 1.25093117e-07 4.99999997 1.25193117e-07 4.99999997 1.25293117e-07 4.99999997
+ 1.25393117e-07 4.99999997 1.25493117e-07 4.99999997 1.25593117e-07 4.99999997 1.25693117e-07 4.99999997 1.25793117e-07 4.99999997 1.25893117e-07 4.99999997 1.25993117e-07 4.99999997 1.26093117e-07 4.99999997
+ 1.26193117e-07 4.99999997 1.26293117e-07 4.99999997 1.26393117e-07 4.99999997 1.26493117e-07 4.99999997 1.26593117e-07 4.99999997 1.26693117e-07 4.99999997 1.26793117e-07 4.99999997 1.26893117e-07 4.99999997
+ 1.26993117e-07 4.99999997 1.27093117e-07 4.99999997 1.27193117e-07 4.99999997 1.27293117e-07 4.99999997 1.27393117e-07 4.99999997 1.27493117e-07 4.99999997 1.27593117e-07 4.99999997 1.27693117e-07 4.99999997
+ 1.27793117e-07 4.99999997 1.27893117e-07 4.99999997 1.27993117e-07 4.99999997 1.28093117e-07 4.99999997 1.28193117e-07 4.99999997 1.28293117e-07 4.99999997 1.28393117e-07 4.99999997 1.28493117e-07 4.99999997
+ 1.28593117e-07 4.99999997 1.28693117e-07 4.99999997 1.28793117e-07 4.99999997 1.28893117e-07 4.99999997 1.28993117e-07 4.99999997 1.29093117e-07 4.99999997 1.29193117e-07 4.99999997 1.29293117e-07 4.99999997
+ 1.29393117e-07 4.99999997 1.29493117e-07 4.99999997 1.29593117e-07 4.99999997 1.29693117e-07 4.99999997 1.29793117e-07 4.99999997 1.29893117e-07 4.99999997 1.29993117e-07 4.99999997 1.30093117e-07 4.99999997
+ 1.30193117e-07 4.99999997 1.30293117e-07 4.99999997 1.30393117e-07 4.99999997 1.30493117e-07 4.99999997 1.30593117e-07 4.99999997 1.30693117e-07 4.99999997 1.30793117e-07 4.99999997 1.30893117e-07 4.99999997
+ 1.30993117e-07 4.99999997 1.31093117e-07 4.99999997 1.31193117e-07 4.99999997 1.31293117e-07 4.99999997 1.31393117e-07 4.99999997 1.31493117e-07 4.99999997 1.31593117e-07 4.99999997 1.31693117e-07 4.99999997
+ 1.31793117e-07 4.99999997 1.31893117e-07 4.99999997 1.31993117e-07 4.99999997 1.32093117e-07 4.99999997 1.32193117e-07 4.99999997 1.32293117e-07 4.99999997 1.32393117e-07 4.99999997 1.32493117e-07 4.99999997
+ 1.32593117e-07 4.99999997 1.32693117e-07 4.99999997 1.32793117e-07 4.99999997 1.32893117e-07 4.99999997 1.32993117e-07 4.99999997 1.33093117e-07 4.99999997 1.33193117e-07 4.99999997 1.33293117e-07 4.99999997
+ 1.33393117e-07 4.99999997 1.33493117e-07 4.99999997 1.33593117e-07 4.99999997 1.33693117e-07 4.99999997 1.33793117e-07 4.99999997 1.33893117e-07 4.99999997 1.33993117e-07 4.99999997 1.34093117e-07 4.99999997
+ 1.34193117e-07 4.99999997 1.34293117e-07 4.99999997 1.34393117e-07 4.99999997 1.34493117e-07 4.99999997 1.34593117e-07 4.99999997 1.34693117e-07 4.99999997 1.34793117e-07 4.99999997 1.34893117e-07 4.99999997
+ 1.34993117e-07 4.99999997 1.35093117e-07 4.99999997 1.35193117e-07 4.99999997 1.35293117e-07 4.99999997 1.35393117e-07 4.99999997 1.35493117e-07 4.99999997 1.35593117e-07 4.99999997 1.35693117e-07 4.99999997
+ 1.35793117e-07 4.99999997 1.35893117e-07 4.99999997 1.35993117e-07 4.99999997 1.36093117e-07 4.99999997 1.36193117e-07 4.99999997 1.36293117e-07 4.99999997 1.36393117e-07 4.99999997 1.36493117e-07 4.99999997
+ 1.36593117e-07 4.99999997 1.36693117e-07 4.99999997 1.36793117e-07 4.99999997 1.36893117e-07 4.99999997 1.36993117e-07 4.99999997 1.37093117e-07 4.99999997 1.37193117e-07 4.99999997 1.37293117e-07 4.99999997
+ 1.37393117e-07 4.99999997 1.37493117e-07 4.99999997 1.37593117e-07 4.99999997 1.37693117e-07 4.99999997 1.37793117e-07 4.99999997 1.37893117e-07 4.99999997 1.37993117e-07 4.99999997 1.38093117e-07 4.99999997
+ 1.38193117e-07 4.99999997 1.38293117e-07 4.99999997 1.38393117e-07 4.99999997 1.38493117e-07 4.99999997 1.38593117e-07 4.99999997 1.38693117e-07 4.99999997 1.38793117e-07 4.99999997 1.38893117e-07 4.99999997
+ 1.38993117e-07 4.99999997 1.39093117e-07 4.99999997 1.39193117e-07 4.99999997 1.39293117e-07 4.99999997 1.39393117e-07 4.99999997 1.39493117e-07 4.99999997 1.39593117e-07 4.99999997 1.39693117e-07 4.99999997
+ 1.39793117e-07 4.99999997 1.39893117e-07 4.99999997 1.39993117e-07 4.99999997 1.40093117e-07 4.99999997 1.40193117e-07 4.99999997 1.40293117e-07 4.99999997 1.40393117e-07 4.99999997 1.40493117e-07 4.99999997
+ 1.40593117e-07 4.99999997 1.40693117e-07 4.99999997 1.40793117e-07 4.99999997 1.40893117e-07 4.99999997 1.40993117e-07 4.99999997 1.41093117e-07 4.99999997 1.41193117e-07 4.99999997 1.41293117e-07 4.99999997
+ 1.41393117e-07 4.99999997 1.41493117e-07 4.99999997 1.41593117e-07 4.99999997 1.41693117e-07 4.99999997 1.41793117e-07 4.99999997 1.41893117e-07 4.99999997 1.41993117e-07 4.99999997 1.42093117e-07 4.99999997
+ 1.42193117e-07 4.99999997 1.42293117e-07 4.99999997 1.42393117e-07 4.99999997 1.42493117e-07 4.99999997 1.42593117e-07 4.99999997 1.42693117e-07 4.99999997 1.42793117e-07 4.99999997 1.42893117e-07 4.99999997
+ 1.42993117e-07 4.99999997 1.43093117e-07 4.99999997 1.43193117e-07 4.99999997 1.43293117e-07 4.99999997 1.43393117e-07 4.99999997 1.43493117e-07 4.99999997 1.43593117e-07 4.99999997 1.43693117e-07 4.99999997
+ 1.43793117e-07 4.99999997 1.43893117e-07 4.99999997 1.43993117e-07 4.99999997 1.44093117e-07 4.99999997 1.44193117e-07 4.99999997 1.44293117e-07 4.99999997 1.44393117e-07 4.99999997 1.44493117e-07 4.99999997
+ 1.44593117e-07 4.99999997 1.44693117e-07 4.99999997 1.44793117e-07 4.99999997 1.44893117e-07 4.99999997 1.44993117e-07 4.99999997 1.45093117e-07 4.99999997 1.45193117e-07 4.99999997 1.45293117e-07 4.99999997
+ 1.45393117e-07 4.99999997 1.45493117e-07 4.99999997 1.45593117e-07 4.99999997 1.45693117e-07 4.99999997 1.45793117e-07 4.99999997 1.45893117e-07 4.99999997 1.45993117e-07 4.99999997 1.46093117e-07 4.99999997
+ 1.46193117e-07 4.99999997 1.46293117e-07 4.99999997 1.46393117e-07 4.99999997 1.46493117e-07 4.99999997 1.46593117e-07 4.99999997 1.46693117e-07 4.99999997 1.46793117e-07 4.99999997 1.46893117e-07 4.99999997
+ 1.46993117e-07 4.99999997 1.47093117e-07 4.99999997 1.47193117e-07 4.99999997 1.47293117e-07 4.99999997 1.47393117e-07 4.99999997 1.47493117e-07 4.99999997 1.47593117e-07 4.99999997 1.47693117e-07 4.99999997
+ 1.47793117e-07 4.99999997 1.47893117e-07 4.99999997 1.47993117e-07 4.99999997 1.48093117e-07 4.99999997 1.48193117e-07 4.99999997 1.48293117e-07 4.99999997 1.48393117e-07 4.99999997 1.48493117e-07 4.99999997
+ 1.48593117e-07 4.99999997 1.48693117e-07 4.99999997 1.48793117e-07 4.99999997 1.48893117e-07 4.99999997 1.48993117e-07 4.99999997 1.49093117e-07 4.99999997 1.49193117e-07 4.99999997 1.49293117e-07 4.99999997
+ 1.49393117e-07 4.99999997 1.49493117e-07 4.99999997 1.49593117e-07 4.99999997 1.49693117e-07 4.99999997 1.49793117e-07 4.99999997 1.49893117e-07 4.99999997 1.49993117e-07 4.99999997 1.50093117e-07 4.99999997
+ 1.50193117e-07 4.99999997 1.50293117e-07 4.99999997 1.50393117e-07 4.99999997 1.50493117e-07 4.99999997 1.50593117e-07 4.99999997 1.50693117e-07 4.99999997 1.50793117e-07 4.99999997 1.50893117e-07 4.99999997
+ 1.50993117e-07 4.99999997 1.51e-07 4.99999997 1.5101e-07 4.99999997 1.5103e-07 4.99999998 1.5107e-07 4.99999996 1.5115e-07 4.99999998 1.5125e-07 4.99999997 1.5135e-07 4.99999997
+ 1.5145e-07 4.99999998 1.5155e-07 4.99999996 1.5165e-07 4.99999998 1.5175e-07 4.99999996 1.5185e-07 4.99999999 1.51930828e-07 5.00006471 1.52e-07 4.99916174 1.52008608e-07 4.99761843
+ 1.52025825e-07 4.99312395 1.52060258e-07 5.01021614 1.52106188e-07 5.09915398 1.52150118e-07 4.21384241 1.5219811e-07 0.290133164 1.52255501e-07 -0.0555601235 1.52312176e-07 0.071992207 1.52404431e-07 -0.0580455459
+ 1.52490774e-07 0.0521266462 1.52590774e-07 -0.046900588 1.52690774e-07 0.042974581 1.52790774e-07 -0.0387934186 1.52890774e-07 0.0355083829 1.52990774e-07 -0.0321185209 1.53090774e-07 0.0293845439 1.53190774e-07 -0.0266224795
+ 1.53290774e-07 0.0243478875 1.53390774e-07 -0.0220883003 1.53490774e-07 0.0201959102 1.53590774e-07 -0.0183413196 1.53690774e-07 0.0167666634 1.53790774e-07 -0.0152403688 1.53890774e-07 0.0139298139 1.53990774e-07 -0.0126709058
+ 1.54090774e-07 0.0115799054 1.54190774e-07 -0.0105396326 1.54290774e-07 0.00963120539 1.54390774e-07 -0.00877029031 1.54490774e-07 0.00801373348 1.54590774e-07 -0.00730035534 1.54690774e-07 0.00667016991 1.54790774e-07 -0.0060784283
+ 1.54890774e-07 0.00555342785 1.54990774e-07 -0.00506215822 1.55090774e-07 0.00462473134 1.55190774e-07 -0.00421658185 1.55290774e-07 0.00385208255 1.55390774e-07 -0.0035127877 1.55490774e-07 0.00320903124 1.55590774e-07 -0.0029268357
+ 1.55690774e-07 0.00267368149 1.55790774e-07 -0.00243887954 1.55890774e-07 0.00222788568 1.55990774e-07 -0.00203245084 1.56090774e-07 0.0018565878 1.56190774e-07 -0.0016938733 1.56290774e-07 0.00154728638 1.56390774e-07 -0.00141178176
+ 1.56490774e-07 0.00128959387 1.56590774e-07 -0.00117672642 1.56690774e-07 0.00107487425 1.56790774e-07 -0.000980846434 1.56890774e-07 0.000895944255 1.56990774e-07 -0.000817600267 1.57090774e-07 0.000746826659 1.57190774e-07 -0.000681542527
+ 1.57290774e-07 0.000622546127 1.57390774e-07 -0.000568139108 1.57490774e-07 0.000518960166 1.57590774e-07 -0.00047361387 1.57690774e-07 0.000432618935 1.57790774e-07 -0.00039482136 1.57890774e-07 0.000360648892 1.57990774e-07 -0.000329141088
+ 1.58090774e-07 0.000300656148 1.58190774e-07 -0.000274389641 1.58290774e-07 0.000250646154 1.58390774e-07 -0.000228747599 1.58490774e-07 0.0002089569 1.58590774e-07 -0.000190698721 1.58690774e-07 0.000174203358 1.58790774e-07 -0.00015897934
+ 1.58890774e-07 0.000145231232 1.58990774e-07 -0.000132536229 1.59090774e-07 0.000121078462 1.59190774e-07 -0.000110491511 1.59290774e-07 0.000100943174 1.59390774e-07 -9.21134357e-05 1.59490774e-07 8.4156973e-05 1.59590774e-07 -7.67920397e-05
+ 1.59690774e-07 7.01627124e-05 1.59790774e-07 -6.40188597e-05 1.59890774e-07 5.84959595e-05 1.59990774e-07 -5.33700348e-05 1.60090774e-07 4.87695597e-05 1.60190774e-07 -4.44922222e-05 1.60290774e-07 4.06607716e-05 1.60390774e-07 -3.70908606e-05
+ 1.60490774e-07 3.39005457e-05 1.60590774e-07 -3.09203885e-05 1.60690774e-07 2.82645887e-05 1.60790774e-07 -2.57760907e-05 1.60890774e-07 2.3565917e-05 1.60990774e-07 -2.14873027e-05 1.61090774e-07 1.96486482e-05 1.61190774e-07 -1.79117455e-05
+ 1.61290774e-07 1.63828276e-05 1.61390774e-07 -1.49308044e-05 1.61490774e-07 1.36601148e-05 1.61590774e-07 -1.24455918e-05 1.61690774e-07 1.1390188e-05 1.61790774e-07 -1.03736667e-05 1.61890774e-07 9.49774736e-06 1.61990774e-07 -8.6462987e-06
+ 1.62090774e-07 7.9200162e-06 1.62190774e-07 -7.20618766e-06 1.62290774e-07 6.60465801e-06 1.62390774e-07 -6.00556286e-06 1.62490774e-07 5.50804017e-06 1.62590774e-07 -5.004598e-06 1.62690774e-07 4.59378634e-06 1.62790774e-07 -4.17008995e-06
+ 1.62890774e-07 3.83156966e-06 1.62990774e-07 -3.47435733e-06 1.63090774e-07 3.19610667e-06 1.63190774e-07 -2.89432215e-06 1.63290774e-07 2.66631855e-06 1.63390774e-07 -2.41074428e-06 1.63490774e-07 2.22463188e-06 1.63590774e-07 -2.00758318e-06
+ 1.63690774e-07 1.85639569e-06 1.63790774e-07 -1.6714659e-06 1.63890774e-07 1.55939899e-06 1.63990774e-07 -1.38082138e-06 1.64090774e-07 1.30227747e-06 1.64190774e-07 -1.14884092e-06 1.64290774e-07 1.08727392e-06 1.64390774e-07 -9.55390911e-07
+ 1.64490774e-07 9.08044283e-07 1.64590774e-07 -7.94134404e-07 1.64690774e-07 7.58642142e-07 1.64790774e-07 -6.59714463e-07 1.64890774e-07 6.34103634e-07 1.64990774e-07 -5.47664793e-07 1.65090774e-07 5.30290583e-07 1.65190774e-07 -4.54262083e-07
+ 1.65290774e-07 4.43753894e-07 1.65390774e-07 -3.764036e-07 1.65490774e-07 3.71618864e-07 1.65590774e-07 -3.1150255e-07 1.65690774e-07 3.11488709e-07 1.65790774e-07 -2.57402481e-07 1.65890774e-07 2.61365518e-07 1.65990774e-07 -2.12307011e-07
+ 1.66090774e-07 2.19586254e-07 1.66190774e-07 -1.74727651e-07 1.66290774e-07 1.84780202e-07 1.66390774e-07 -1.43421281e-07 1.66490774e-07 1.55784186e-07 1.66590774e-07 -1.17340694e-07 1.66690774e-07 1.3162823e-07 1.66790774e-07 -9.56134643e-08
+ 1.66890774e-07 1.11504323e-07 1.66990774e-07 -7.75128519e-08 1.67090774e-07 9.4739428e-08 1.67190774e-07 -6.24336457e-08 1.67290774e-07 8.07731335e-08 1.67390774e-07 -4.98334138e-08 1.67490774e-07 6.90993792e-08 1.67590774e-07 -3.93732592e-08
+ 1.67690774e-07 5.94152844e-08 1.67790774e-07 -3.06632472e-08 1.67890774e-07 5.13482986e-08 1.67990774e-07 -2.34074247e-08 1.68090774e-07 4.46281627e-08 1.68190774e-07 -1.73630594e-08 1.68290774e-07 3.90298631e-08 1.68390774e-07 -1.23273488e-08
+ 1.68490774e-07 3.436586e-08 1.68590774e-07 -8.13252579e-09 1.68690774e-07 3.048091e-08 1.68790774e-07 -4.63838543e-09 1.68890774e-07 2.7244872e-08 1.68990774e-07 -1.72786965e-09 1.69090774e-07 2.45493396e-08 1.69190774e-07 6.96518204e-10
+ 1.69290774e-07 2.23131567e-08 1.69390774e-07 2.70818359e-09 1.69490774e-07 2.0476404e-08 1.69590774e-07 4.36139963e-09 1.69690774e-07 1.89668152e-08 1.69790774e-07 5.720181e-09 1.69890774e-07 1.77260561e-08 1.69990774e-07 6.83700896e-09
+ 1.70090774e-07 1.67062182e-08 1.70190774e-07 7.75499595e-09 1.70290774e-07 1.58679406e-08 1.70390774e-07 8.50956494e-09 1.70490774e-07 1.50799957e-08 1.70590774e-07 9.11601344e-09 1.70690774e-07 1.45257675e-08 1.70790774e-07 9.61910654e-09
+ 1.70890774e-07 1.40694266e-08 1.70990774e-07 1.00330061e-08 1.71090774e-07 1.36940245e-08 1.71190774e-07 1.03734906e-08 1.71290774e-07 1.33852096e-08 1.71390774e-07 1.06535815e-08 1.71490774e-07 1.31311713e-08 1.71590774e-07 1.08839909e-08
+ 1.71690774e-07 1.2922193e-08 1.71790774e-07 1.10735315e-08 1.71890774e-07 1.27502824e-08 1.71990774e-07 1.12294524e-08 1.72090774e-07 1.2608864e-08 1.72190774e-07 1.13577175e-08 1.72290774e-07 1.24925287e-08 1.72390774e-07 1.14632322e-08
+ 1.72490774e-07 1.23968278e-08 1.72590774e-07 1.15500321e-08 1.72690774e-07 1.23181005e-08 1.72790774e-07 1.16214377e-08 1.72890774e-07 1.22533359e-08 1.72990774e-07 1.16801792e-08 1.73090774e-07 1.22000571e-08 1.73190774e-07 1.17285027e-08
+ 1.73290774e-07 1.21562274e-08 1.73390774e-07 1.17682566e-08 1.73490774e-07 1.21201702e-08 1.73590774e-07 1.18009613e-08 1.73690774e-07 1.20905069e-08 1.73790774e-07 1.18278666e-08 1.73890774e-07 1.20661032e-08 1.73990774e-07 1.18500008e-08
+ 1.74090774e-07 1.20460268e-08 1.74190774e-07 1.18682109e-08 1.74290774e-07 1.20295097e-08 1.74390774e-07 1.18831926e-08 1.74490774e-07 1.20159204e-08 1.74590774e-07 1.18955188e-08 1.74690774e-07 1.20047403e-08 1.74790774e-07 1.19056596e-08
+ 1.74890774e-07 1.19955419e-08 1.74990774e-07 1.19140031e-08 1.75090774e-07 1.19879738e-08 1.75190774e-07 1.19208679e-08 1.75290774e-07 1.1981747e-08 1.75390774e-07 1.19265162e-08 1.75490774e-07 1.19766235e-08 1.75590774e-07 1.19311639e-08
+ 1.75690774e-07 1.19724075e-08 1.75790774e-07 1.19349879e-08 1.75890774e-07 1.19689385e-08 1.75990774e-07 1.19381348e-08 1.76090774e-07 1.19660841e-08 1.76190774e-07 1.19407247e-08 1.76290774e-07 1.19637348e-08 1.76390774e-07 1.19428556e-08
+ 1.76490774e-07 1.19618016e-08 1.76590774e-07 1.19446091e-08 1.76690774e-07 1.19602107e-08 1.76790774e-07 1.19460526e-08 1.76890774e-07 1.19589012e-08 1.76990774e-07 1.19472407e-08 1.77090774e-07 1.19578233e-08 1.77190774e-07 1.19482185e-08
+ 1.77290774e-07 1.1956936e-08 1.77390774e-07 1.19490234e-08 1.77490774e-07 1.19562059e-08 1.77590774e-07 1.19496864e-08 1.77690774e-07 1.19556045e-08 1.77790774e-07 1.19502317e-08 1.77890774e-07 1.19551092e-08 1.77990774e-07 1.19506811e-08
+ 1.78090774e-07 1.19547014e-08 1.78190774e-07 1.19510511e-08 1.78290774e-07 1.19543659e-08 1.78390774e-07 1.19513556e-08 1.78490774e-07 1.19540894e-08 1.78590774e-07 1.19516065e-08 1.78690774e-07 1.19538617e-08 1.78790774e-07 1.1951813e-08
+ 1.78890774e-07 1.19536742e-08 1.78990774e-07 1.19519834e-08 1.79090774e-07 1.19535196e-08 1.79190774e-07 1.19521238e-08 1.79290774e-07 1.19533921e-08 1.79390774e-07 1.19522396e-08 1.79490774e-07 1.1953287e-08 1.79590774e-07 1.19523348e-08
+ 1.79690774e-07 1.19532003e-08 1.79790774e-07 1.19524138e-08 1.79890774e-07 1.19531291e-08 1.79990774e-07 1.19524785e-08 1.80090774e-07 1.19530701e-08 1.80190774e-07 1.1952532e-08 1.80290774e-07 1.19530215e-08 1.80390774e-07 1.19525758e-08
+ 1.80490774e-07 1.19529818e-08 1.80590774e-07 1.19526124e-08 1.80690774e-07 1.19529486e-08 1.80790774e-07 1.19526426e-08 1.80890774e-07 1.19529211e-08 1.80990774e-07 1.19526673e-08 1.81090774e-07 1.19528986e-08 1.81190774e-07 1.19526879e-08
+ 1.81290774e-07 1.19528798e-08 1.81390774e-07 1.19527048e-08 1.81490774e-07 1.19528644e-08 1.81590774e-07 1.19527192e-08 1.81690774e-07 1.19528517e-08 1.81790774e-07 1.19527306e-08 1.81890774e-07 1.1952841e-08 1.81990774e-07 1.19527407e-08
+ 1.82090774e-07 1.19528321e-08 1.82190774e-07 1.19527485e-08 1.82290774e-07 1.19528246e-08 1.82390774e-07 1.1952755e-08 1.82490774e-07 1.19528188e-08 1.82590774e-07 1.19527605e-08 1.82690774e-07 1.19528139e-08 1.82790774e-07 1.1952765e-08
+ 1.82890774e-07 1.19528099e-08 1.82990774e-07 1.19527688e-08 1.83090774e-07 1.1952806e-08 1.83190774e-07 1.1952772e-08 1.83290774e-07 1.19528032e-08 1.83390774e-07 1.19527746e-08 1.83490774e-07 1.19528008e-08 1.83590774e-07 1.19527764e-08
+ 1.83690774e-07 1.19527989e-08 1.83790774e-07 1.19527782e-08 1.83890774e-07 1.19527976e-08 1.83990774e-07 1.19527796e-08 1.84090774e-07 1.19527961e-08 1.84190774e-07 1.19527813e-08 1.84290774e-07 1.19527948e-08 1.84390774e-07 1.19527825e-08
+ 1.84490774e-07 1.19527939e-08 1.84590774e-07 1.19527832e-08 1.84690774e-07 1.19527932e-08 1.84790774e-07 1.19527839e-08 1.84890774e-07 1.19527923e-08 1.84990774e-07 1.19527844e-08 1.85090774e-07 1.19527919e-08 1.85190774e-07 1.19527849e-08
+ 1.85290774e-07 1.19527913e-08 1.85390774e-07 1.19527856e-08 1.85490774e-07 1.19527907e-08 1.85590774e-07 1.19527861e-08 1.85690774e-07 1.19527904e-08 1.85790774e-07 1.19527864e-08 1.85890774e-07 1.195279e-08 1.85990774e-07 1.19527868e-08
+ 1.86090774e-07 1.19527899e-08 1.86190774e-07 1.1952787e-08 1.86290774e-07 1.19527897e-08 1.86390774e-07 1.1952787e-08 1.86490774e-07 1.19527893e-08 1.86590774e-07 1.19527872e-08 1.86690774e-07 1.19527894e-08 1.86790774e-07 1.19527873e-08
+ 1.86890774e-07 1.19527893e-08 1.86990774e-07 1.19527874e-08 1.87090774e-07 1.19527892e-08 1.87190774e-07 1.19527875e-08 1.87290774e-07 1.19527892e-08 1.87390774e-07 1.19527875e-08 1.87490774e-07 1.19527892e-08 1.87590774e-07 1.19527876e-08
+ 1.87690774e-07 1.1952789e-08 1.87790774e-07 1.19527877e-08 1.87890774e-07 1.19527891e-08 1.87990774e-07 1.19527877e-08 1.88090774e-07 1.1952789e-08 1.88190774e-07 1.19527878e-08 1.88290774e-07 1.1952789e-08 1.88390774e-07 1.19527879e-08
+ 1.88490774e-07 1.19527888e-08 1.88590774e-07 1.1952788e-08 1.88690774e-07 1.19527889e-08 1.88790774e-07 1.19527879e-08 1.88890774e-07 1.19527888e-08 1.88990774e-07 1.1952788e-08 1.89090774e-07 1.19527888e-08 1.89190774e-07 1.19527881e-08
+ 1.89290774e-07 1.19527888e-08 1.89390774e-07 1.1952788e-08 1.89490774e-07 1.19527887e-08 1.89590774e-07 1.19527882e-08 1.89690774e-07 1.19527887e-08 1.89790774e-07 1.19527881e-08 1.89890774e-07 1.19527886e-08 1.89990774e-07 1.19527882e-08
+ 1.90090774e-07 1.19527887e-08 1.90190774e-07 1.19527881e-08 1.90290774e-07 1.19527886e-08 1.90390774e-07 1.19527882e-08 1.90490774e-07 1.19527886e-08 1.90590774e-07 1.19527883e-08 1.90690774e-07 1.19527885e-08 1.90790774e-07 1.19527881e-08
+ 1.90890774e-07 1.19527887e-08 1.90990774e-07 1.19527882e-08 1.91090774e-07 1.19527886e-08 1.91190774e-07 1.19527881e-08 1.91290774e-07 1.19527886e-08 1.91390774e-07 1.19527882e-08 1.91490774e-07 1.19527886e-08 1.91590774e-07 1.19527882e-08
+ 1.91690774e-07 1.19527885e-08 1.91790774e-07 1.19527882e-08 1.91890774e-07 1.19527885e-08 1.91990774e-07 1.19527883e-08 1.92090774e-07 1.19527884e-08 1.92190774e-07 1.19527883e-08 1.92290774e-07 1.19527885e-08 1.92390774e-07 1.19527883e-08
+ 1.92490774e-07 1.19527884e-08 1.92590774e-07 1.19527883e-08 1.92690774e-07 1.19527884e-08 1.92790774e-07 1.19527883e-08 1.92890774e-07 1.19527884e-08 1.92990774e-07 1.19527883e-08 1.93090774e-07 1.19527884e-08 1.93190774e-07 1.19527883e-08
+ 1.93290774e-07 1.19527884e-08 1.93390774e-07 1.19527883e-08 1.93490774e-07 1.19527884e-08 1.93590774e-07 1.19527883e-08 1.93690774e-07 1.19527884e-08 1.93790774e-07 1.19527883e-08 1.93890774e-07 1.19527884e-08 1.93990774e-07 1.19527883e-08
+ 1.94090774e-07 1.19527884e-08 1.94190774e-07 1.19527883e-08 1.94290774e-07 1.19527884e-08 1.94390774e-07 1.19527883e-08 1.94490774e-07 1.19527884e-08 1.94590774e-07 1.19527883e-08 1.94690774e-07 1.19527884e-08 1.94790774e-07 1.19527883e-08
+ 1.94890774e-07 1.19527884e-08 1.94990774e-07 1.19527883e-08 1.95090774e-07 1.19527884e-08 1.95190774e-07 1.19527883e-08 1.95290774e-07 1.19527884e-08 1.95390774e-07 1.19527883e-08 1.95490774e-07 1.19527884e-08 1.95590774e-07 1.19527883e-08
+ 1.95690774e-07 1.19527884e-08 1.95790774e-07 1.19527883e-08 1.95890774e-07 1.19527884e-08 1.95990774e-07 1.19527883e-08 1.96090774e-07 1.19527884e-08 1.96190774e-07 1.19527883e-08 1.96290774e-07 1.19527884e-08 1.96390774e-07 1.19527883e-08
+ 1.96490774e-07 1.19527884e-08 1.96590774e-07 1.19527883e-08 1.96690774e-07 1.19527884e-08 1.96790774e-07 1.19527883e-08 1.96890774e-07 1.19527884e-08 1.96990774e-07 1.19527883e-08 1.97090774e-07 1.19527884e-08 1.97190774e-07 1.19527883e-08
+ 1.97290774e-07 1.19527884e-08 1.97390774e-07 1.19527883e-08 1.97490774e-07 1.19527884e-08 1.97590774e-07 1.19527883e-08 1.97690774e-07 1.19527884e-08 1.97790774e-07 1.19527883e-08 1.97890774e-07 1.19527884e-08 1.97990774e-07 1.19527883e-08
+ 1.98090774e-07 1.19527884e-08 1.98190774e-07 1.19527883e-08 1.98290774e-07 1.19527884e-08 1.98390774e-07 1.19527883e-08 1.98490774e-07 1.19527884e-08 1.98590774e-07 1.19527883e-08 1.98690774e-07 1.19527884e-08 1.98790774e-07 1.19527883e-08
+ 1.98890774e-07 1.19527884e-08 1.98990774e-07 1.19527883e-08 1.99090774e-07 1.19527884e-08 1.99190774e-07 1.19527883e-08 1.99290774e-07 1.19527884e-08 1.99390774e-07 1.19527883e-08 1.99490774e-07 1.19527884e-08 1.99590774e-07 1.19527883e-08
+ 1.99690774e-07 1.19527884e-08 1.99790774e-07 1.19527883e-08 1.99890774e-07 1.19527884e-08 1.99990774e-07 1.19527883e-08 2e-07 1.19527881e-08 2.0001e-07 1.45272737e-08 2.0003e-07 1.2360668e-09 2.0007e-07 2.76445089e-08
+ 2.0015e-07 -4.38735057e-09 2.0025e-07 2.8215468e-08 2.0035e-07 -3.1892709e-09 2.0045e-07 2.52177597e-08 2.0055e-07 2.59408278e-09 2.0065e-07 -4.06359279e-08 2.0075e-07 3.06902814e-06 2.0085e-07 9.48375612e-05
+ 2.00932239e-07 -0.0448088436 2.01e-07 1.97425329 2.01008502e-07 3.1007477 2.01025505e-07 4.14453646 2.01059511e-07 4.88397722 2.01090728e-07 4.98064226 2.01143656e-07 5.00336705 2.01199398e-07 4.99900033
+ 2.01276452e-07 5.00049859 2.01342062e-07 4.99975148 2.01411951e-07 5.00013732 2.01487979e-07 4.99991579 2.01566956e-07 5.00005277 2.01643585e-07 4.99996651 2.01743585e-07 5.00002357 2.01843585e-07 4.9999831
+ 2.01943585e-07 5.00001203 2.02043585e-07 4.99999123 2.02143585e-07 5.00000632 2.02243585e-07 4.99999529 2.02343585e-07 5.00000343 2.02443585e-07 4.99999737 2.02543585e-07 5.00000193 2.02643585e-07 4.99999847
+ 2.02743585e-07 5.00000113 2.02843585e-07 4.99999907 2.02943585e-07 5.00000068 2.03043585e-07 4.99999941 2.03143585e-07 5.00000042 2.03243585e-07 4.99999961 2.03343585e-07 5.00000026 2.03443585e-07 4.99999974
+ 2.03543585e-07 5.00000017 2.03643585e-07 4.99999981 2.03743585e-07 5.0000001 2.03843585e-07 4.99999986 2.03943585e-07 5.00000006 2.04043585e-07 4.9999999 2.04143585e-07 5.00000003 2.04243585e-07 4.99999992
+ 2.04343585e-07 5.00000001 2.04443585e-07 4.99999994 2.04543585e-07 5.0 2.04643585e-07 4.99999995 2.04743585e-07 4.99999999 2.04843585e-07 4.99999996 2.04943585e-07 4.99999999 2.05043585e-07 4.99999996
+ 2.05143585e-07 4.99999998 2.05243585e-07 4.99999996 2.05343585e-07 4.99999998 2.05443585e-07 4.99999997 2.05543585e-07 4.99999998 2.05643585e-07 4.99999997 2.05743585e-07 4.99999998 2.05843585e-07 4.99999997
+ 2.05943585e-07 4.99999997 2.06043585e-07 4.99999997 2.06143585e-07 4.99999997 2.06243585e-07 4.99999997 2.06343585e-07 4.99999997 2.06443585e-07 4.99999997 2.06543585e-07 4.99999997 2.06643585e-07 4.99999997
+ 2.06743585e-07 4.99999997 2.06843585e-07 4.99999997 2.06943585e-07 4.99999997 2.07043585e-07 4.99999997 2.07143585e-07 4.99999997 2.07243585e-07 4.99999997 2.07343585e-07 4.99999997 2.07443585e-07 4.99999997
+ 2.07543585e-07 4.99999997 2.07643585e-07 4.99999997 2.07743585e-07 4.99999997 2.07843585e-07 4.99999997 2.07943585e-07 4.99999997 2.08043585e-07 4.99999997 2.08143585e-07 4.99999997 2.08243585e-07 4.99999997
+ 2.08343585e-07 4.99999997 2.08443585e-07 4.99999997 2.08543585e-07 4.99999997 2.08643585e-07 4.99999997 2.08743585e-07 4.99999997 2.08843585e-07 4.99999997 2.08943585e-07 4.99999997 2.09043585e-07 4.99999997
+ 2.09143585e-07 4.99999997 2.09243585e-07 4.99999997 2.09343585e-07 4.99999997 2.09443585e-07 4.99999997 2.09543585e-07 4.99999997 2.09643585e-07 4.99999997 2.09743585e-07 4.99999997 2.09843585e-07 4.99999997
+ 2.09943585e-07 4.99999997 2.10043585e-07 4.99999997 2.10143585e-07 4.99999997 2.10243585e-07 4.99999997 2.10343585e-07 4.99999997 2.10443585e-07 4.99999997 2.10543585e-07 4.99999997 2.10643585e-07 4.99999997
+ 2.10743585e-07 4.99999997 2.10843585e-07 4.99999997 2.10943585e-07 4.99999997 2.11043585e-07 4.99999997 2.11143585e-07 4.99999997 2.11243585e-07 4.99999997 2.11343585e-07 4.99999997 2.11443585e-07 4.99999997
+ 2.11543585e-07 4.99999997 2.11643585e-07 4.99999997 2.11743585e-07 4.99999997 2.11843585e-07 4.99999997 2.11943585e-07 4.99999997 2.12043585e-07 4.99999997 2.12143585e-07 4.99999997 2.12243585e-07 4.99999997
+ 2.12343585e-07 4.99999997 2.12443585e-07 4.99999997 2.12543585e-07 4.99999997 2.12643585e-07 4.99999997 2.12743585e-07 4.99999997 2.12843585e-07 4.99999997 2.12943585e-07 4.99999997 2.13043585e-07 4.99999997
+ 2.13143585e-07 4.99999997 2.13243585e-07 4.99999997 2.13343585e-07 4.99999997 2.13443585e-07 4.99999997 2.13543585e-07 4.99999997 2.13643585e-07 4.99999997 2.13743585e-07 4.99999997 2.13843585e-07 4.99999997
+ 2.13943585e-07 4.99999997 2.14043585e-07 4.99999997 2.14143585e-07 4.99999997 2.14243585e-07 4.99999997 2.14343585e-07 4.99999997 2.14443585e-07 4.99999997 2.14543585e-07 4.99999997 2.14643585e-07 4.99999997
+ 2.14743585e-07 4.99999997 2.14843585e-07 4.99999997 2.14943585e-07 4.99999997 2.15043585e-07 4.99999997 2.15143585e-07 4.99999997 2.15243585e-07 4.99999997 2.15343585e-07 4.99999997 2.15443585e-07 4.99999997
+ 2.15543585e-07 4.99999997 2.15643585e-07 4.99999997 2.15743585e-07 4.99999997 2.15843585e-07 4.99999997 2.15943585e-07 4.99999997 2.16043585e-07 4.99999997 2.16143585e-07 4.99999997 2.16243585e-07 4.99999997
+ 2.16343585e-07 4.99999997 2.16443585e-07 4.99999997 2.16543585e-07 4.99999997 2.16643585e-07 4.99999997 2.16743585e-07 4.99999997 2.16843585e-07 4.99999997 2.16943585e-07 4.99999997 2.17043585e-07 4.99999997
+ 2.17143585e-07 4.99999997 2.17243585e-07 4.99999997 2.17343585e-07 4.99999997 2.17443585e-07 4.99999997 2.17543585e-07 4.99999997 2.17643585e-07 4.99999997 2.17743585e-07 4.99999997 2.17843585e-07 4.99999997
+ 2.17943585e-07 4.99999997 2.18043585e-07 4.99999997 2.18143585e-07 4.99999997 2.18243585e-07 4.99999997 2.18343585e-07 4.99999997 2.18443585e-07 4.99999997 2.18543585e-07 4.99999997 2.18643585e-07 4.99999997
+ 2.18743585e-07 4.99999997 2.18843585e-07 4.99999997 2.18943585e-07 4.99999997 2.19043585e-07 4.99999997 2.19143585e-07 4.99999997 2.19243585e-07 4.99999997 2.19343585e-07 4.99999997 2.19443585e-07 4.99999997
+ 2.19543585e-07 4.99999997 2.19643585e-07 4.99999997 2.19743585e-07 4.99999997 2.19843585e-07 4.99999997 2.19943585e-07 4.99999997 2.20043585e-07 4.99999997 2.20143585e-07 4.99999997 2.20243585e-07 4.99999997
+ 2.20343585e-07 4.99999997 2.20443585e-07 4.99999997 2.20543585e-07 4.99999997 2.20643585e-07 4.99999997 2.20743585e-07 4.99999997 2.20843585e-07 4.99999997 2.20943585e-07 4.99999997 2.21043585e-07 4.99999997
+ 2.21143585e-07 4.99999997 2.21243585e-07 4.99999997 2.21343585e-07 4.99999997 2.21443585e-07 4.99999997 2.21543585e-07 4.99999997 2.21643585e-07 4.99999997 2.21743585e-07 4.99999997 2.21843585e-07 4.99999997
+ 2.21943585e-07 4.99999997 2.22043585e-07 4.99999997 2.22143585e-07 4.99999997 2.22243585e-07 4.99999997 2.22343585e-07 4.99999997 2.22443585e-07 4.99999997 2.22543585e-07 4.99999997 2.22643585e-07 4.99999997
+ 2.22743585e-07 4.99999997 2.22843585e-07 4.99999997 2.22943585e-07 4.99999997 2.23043585e-07 4.99999997 2.23143585e-07 4.99999997 2.23243585e-07 4.99999997 2.23343585e-07 4.99999997 2.23443585e-07 4.99999997
+ 2.23543585e-07 4.99999997 2.23643585e-07 4.99999997 2.23743585e-07 4.99999997 2.23843585e-07 4.99999997 2.23943585e-07 4.99999997 2.24043585e-07 4.99999997 2.24143585e-07 4.99999997 2.24243585e-07 4.99999997
+ 2.24343585e-07 4.99999997 2.24443585e-07 4.99999997 2.24543585e-07 4.99999997 2.24643585e-07 4.99999997 2.24743585e-07 4.99999997 2.24843585e-07 4.99999997 2.24943585e-07 4.99999997 2.25043585e-07 4.99999997
+ 2.25143585e-07 4.99999997 2.25243585e-07 4.99999997 2.25343585e-07 4.99999997 2.25443585e-07 4.99999997 2.25543585e-07 4.99999997 2.25643585e-07 4.99999997 2.25743585e-07 4.99999997 2.25843585e-07 4.99999997
+ 2.25943585e-07 4.99999997 2.26043585e-07 4.99999997 2.26143585e-07 4.99999997 2.26243585e-07 4.99999997 2.26343585e-07 4.99999997 2.26443585e-07 4.99999997 2.26543585e-07 4.99999997 2.26643585e-07 4.99999997
+ 2.26743585e-07 4.99999997 2.26843585e-07 4.99999997 2.26943585e-07 4.99999997 2.27043585e-07 4.99999997 2.27143585e-07 4.99999997 2.27243585e-07 4.99999997 2.27343585e-07 4.99999997 2.27443585e-07 4.99999997
+ 2.27543585e-07 4.99999997 2.27643585e-07 4.99999997 2.27743585e-07 4.99999997 2.27843585e-07 4.99999997 2.27943585e-07 4.99999997 2.28043585e-07 4.99999997 2.28143585e-07 4.99999997 2.28243585e-07 4.99999997
+ 2.28343585e-07 4.99999997 2.28443585e-07 4.99999997 2.28543585e-07 4.99999997 2.28643585e-07 4.99999997 2.28743585e-07 4.99999997 2.28843585e-07 4.99999997 2.28943585e-07 4.99999997 2.29043585e-07 4.99999997
+ 2.29143585e-07 4.99999997 2.29243585e-07 4.99999997 2.29343585e-07 4.99999997 2.29443585e-07 4.99999997 2.29543585e-07 4.99999997 2.29643585e-07 4.99999997 2.29743585e-07 4.99999997 2.29843585e-07 4.99999997
+ 2.29943585e-07 4.99999997 2.30043585e-07 4.99999997 2.30143585e-07 4.99999997 2.30243585e-07 4.99999997 2.30343585e-07 4.99999997 2.30443585e-07 4.99999997 2.30543585e-07 4.99999997 2.30643585e-07 4.99999997
+ 2.30743585e-07 4.99999997 2.30843585e-07 4.99999997 2.30943585e-07 4.99999997 2.31043585e-07 4.99999997 2.31143585e-07 4.99999997 2.31243585e-07 4.99999997 2.31343585e-07 4.99999997 2.31443585e-07 4.99999997
+ 2.31543585e-07 4.99999997 2.31643585e-07 4.99999997 2.31743585e-07 4.99999997 2.31843585e-07 4.99999997 2.31943585e-07 4.99999997 2.32043585e-07 4.99999997 2.32143585e-07 4.99999997 2.32243585e-07 4.99999997
+ 2.32343585e-07 4.99999997 2.32443585e-07 4.99999997 2.32543585e-07 4.99999997 2.32643585e-07 4.99999997 2.32743585e-07 4.99999997 2.32843585e-07 4.99999997 2.32943585e-07 4.99999997 2.33043585e-07 4.99999997
+ 2.33143585e-07 4.99999997 2.33243585e-07 4.99999997 2.33343585e-07 4.99999997 2.33443585e-07 4.99999997 2.33543585e-07 4.99999997 2.33643585e-07 4.99999997 2.33743585e-07 4.99999997 2.33843585e-07 4.99999997
+ 2.33943585e-07 4.99999997 2.34043585e-07 4.99999997 2.34143585e-07 4.99999997 2.34243585e-07 4.99999997 2.34343585e-07 4.99999997 2.34443585e-07 4.99999997 2.34543585e-07 4.99999997 2.34643585e-07 4.99999997
+ 2.34743585e-07 4.99999997 2.34843585e-07 4.99999997 2.34943585e-07 4.99999997 2.35043585e-07 4.99999997 2.35143585e-07 4.99999997 2.35243585e-07 4.99999997 2.35343585e-07 4.99999997 2.35443585e-07 4.99999997
+ 2.35543585e-07 4.99999997 2.35643585e-07 4.99999997 2.35743585e-07 4.99999997 2.35843585e-07 4.99999997 2.35943585e-07 4.99999997 2.36043585e-07 4.99999997 2.36143585e-07 4.99999997 2.36243585e-07 4.99999997
+ 2.36343585e-07 4.99999997 2.36443585e-07 4.99999997 2.36543585e-07 4.99999997 2.36643585e-07 4.99999997 2.36743585e-07 4.99999997 2.36843585e-07 4.99999997 2.36943585e-07 4.99999997 2.37043585e-07 4.99999997
+ 2.37143585e-07 4.99999997 2.37243585e-07 4.99999997 2.37343585e-07 4.99999997 2.37443585e-07 4.99999997 2.37543585e-07 4.99999997 2.37643585e-07 4.99999997 2.37743585e-07 4.99999997 2.37843585e-07 4.99999997
+ 2.37943585e-07 4.99999997 2.38043585e-07 4.99999997 2.38143585e-07 4.99999997 2.38243585e-07 4.99999997 2.38343585e-07 4.99999997 2.38443585e-07 4.99999997 2.38543585e-07 4.99999997 2.38643585e-07 4.99999997
+ 2.38743585e-07 4.99999997 2.38843585e-07 4.99999997 2.38943585e-07 4.99999997 2.39043585e-07 4.99999997 2.39143585e-07 4.99999997 2.39243585e-07 4.99999997 2.39343585e-07 4.99999997 2.39443585e-07 4.99999997
+ 2.39543585e-07 4.99999997 2.39643585e-07 4.99999997 2.39743585e-07 4.99999997 2.39843585e-07 4.99999997 2.39943585e-07 4.99999997 2.40043585e-07 4.99999997 2.40143585e-07 4.99999997 2.40243585e-07 4.99999997
+ 2.40343585e-07 4.99999997 2.40443585e-07 4.99999997 2.40543585e-07 4.99999997 2.40643585e-07 4.99999997 2.40743585e-07 4.99999997 2.40843585e-07 4.99999997 2.40943585e-07 4.99999997 2.41043585e-07 4.99999997
+ 2.41143585e-07 4.99999997 2.41243585e-07 4.99999997 2.41343585e-07 4.99999997 2.41443585e-07 4.99999997 2.41543585e-07 4.99999997 2.41643585e-07 4.99999997 2.41743585e-07 4.99999997 2.41843585e-07 4.99999997
+ 2.41943585e-07 4.99999997 2.42043585e-07 4.99999997 2.42143585e-07 4.99999997 2.42243585e-07 4.99999997 2.42343585e-07 4.99999997 2.42443585e-07 4.99999997 2.42543585e-07 4.99999997 2.42643585e-07 4.99999997
+ 2.42743585e-07 4.99999997 2.42843585e-07 4.99999997 2.42943585e-07 4.99999997 2.43043585e-07 4.99999997 2.43143585e-07 4.99999997 2.43243585e-07 4.99999997 2.43343585e-07 4.99999997 2.43443585e-07 4.99999997
+ 2.43543585e-07 4.99999997 2.43643585e-07 4.99999997 2.43743585e-07 4.99999997 2.43843585e-07 4.99999997 2.43943585e-07 4.99999997 2.44043585e-07 4.99999997 2.44143585e-07 4.99999997 2.44243585e-07 4.99999997
+ 2.44343585e-07 4.99999997 2.44443585e-07 4.99999997 2.44543585e-07 4.99999997 2.44643585e-07 4.99999997 2.44743585e-07 4.99999997 2.44843585e-07 4.99999997 2.44943585e-07 4.99999997 2.45043585e-07 4.99999997
+ 2.45143585e-07 4.99999997 2.45243585e-07 4.99999997 2.45343585e-07 4.99999997 2.45443585e-07 4.99999997 2.45543585e-07 4.99999997 2.45643585e-07 4.99999997 2.45743585e-07 4.99999997 2.45843585e-07 4.99999997
+ 2.45943585e-07 4.99999997 2.46043585e-07 4.99999997 2.46143585e-07 4.99999997 2.46243585e-07 4.99999997 2.46343585e-07 4.99999997 2.46443585e-07 4.99999997 2.46543585e-07 4.99999997 2.46643585e-07 4.99999997
+ 2.46743585e-07 4.99999997 2.46843585e-07 4.99999997 2.46943585e-07 4.99999997 2.47043585e-07 4.99999997 2.47143585e-07 4.99999997 2.47243585e-07 4.99999997 2.47343585e-07 4.99999997 2.47443585e-07 4.99999997
+ 2.47543585e-07 4.99999997 2.47643585e-07 4.99999997 2.47743585e-07 4.99999997 2.47843585e-07 4.99999997 2.47943585e-07 4.99999997 2.48043585e-07 4.99999997 2.48143585e-07 4.99999997 2.48243585e-07 4.99999997
+ 2.48343585e-07 4.99999997 2.48443585e-07 4.99999997 2.48543585e-07 4.99999997 2.48643585e-07 4.99999997 2.48743585e-07 4.99999997 2.48843585e-07 4.99999997 2.48943585e-07 4.99999997 2.49043585e-07 4.99999997
+ 2.49143585e-07 4.99999997 2.49243585e-07 4.99999997 2.49343585e-07 4.99999997 2.49443585e-07 4.99999997 2.49543585e-07 4.99999997 2.49643585e-07 4.99999997 2.49743585e-07 4.99999997 2.49843585e-07 4.99999997
+ 2.49943585e-07 4.99999997 2.50043585e-07 4.99999997 2.50143585e-07 4.99999997 2.50243585e-07 4.99999997 2.50343585e-07 4.99999997 2.50443585e-07 4.99999997 2.50543585e-07 4.99999997 2.50643585e-07 4.99999997
+ 2.50743585e-07 4.99999997 2.50843585e-07 4.99999997 2.50943585e-07 4.99999997 2.51e-07 4.99999997 2.5101e-07 4.99999997 2.5103e-07 4.99999998 2.5107e-07 4.99999996 2.5115e-07 4.99999998
+ 2.5125e-07 4.99999997 2.5135e-07 4.99999997 2.5145e-07 4.99999998 2.5155e-07 4.99999996 2.5165e-07 4.99999998 2.5175e-07 4.99999996 2.5185e-07 4.99999999 2.51930828e-07 5.00006476
+ 2.52e-07 4.99916064 2.52008608e-07 4.99761638 2.52025825e-07 4.99311194 2.52060258e-07 5.01027326 2.52106181e-07 5.09906166 2.52150081e-07 4.21228987 2.52198026e-07 0.290284563 2.5225538e-07 -0.0554589573
+ 2.52312019e-07 0.0719466825 2.52404231e-07 -0.0579814231 2.52504231e-07 0.052890252 2.52604231e-07 -0.0475728397 2.52704231e-07 0.0435755801 2.52804231e-07 -0.0393282951 2.52904231e-07 0.0359988053 2.53004231e-07 -0.0325571519
+ 2.53104231e-07 0.029786221 2.53204231e-07 -0.0269830488 2.53304231e-07 0.0246778153 2.53404231e-07 -0.0223853345 2.53504231e-07 0.0204675598 2.53604231e-07 -0.0185864689 2.53704231e-07 0.0169907803 2.53804231e-07 -0.0154430156
+ 2.53904231e-07 0.0141150275 2.54004231e-07 -0.0128386436 2.54104231e-07 0.0117331852 2.54204231e-07 -0.0106786325 2.54304231e-07 0.00975820759 2.54404231e-07 -0.00888558601 2.54504231e-07 0.00811906716 2.54604231e-07 -0.00739606596
+ 2.54704231e-07 0.00675760434 2.54804231e-07 -0.00615793428 2.54904231e-07 0.00562605481 2.55004231e-07 -0.00512824045 2.55104231e-07 0.00468509345 2.55204231e-07 -0.0042715328 2.55304231e-07 0.00390227528 2.55404231e-07 -0.00355850054
+ 2.55504231e-07 0.00325078477 2.55604231e-07 -0.00296487618 2.55704231e-07 0.00270842653 2.55804231e-07 -0.00247054424 2.55904231e-07 0.00225680687 2.56004231e-07 -0.00205881459 2.56104231e-07 0.00188066709 2.56204231e-07 -0.0017158279
+ 2.56304231e-07 0.00156733843 2.56404231e-07 -0.00143006768 2.56504231e-07 0.00130629509 2.56604231e-07 -0.00119195888 2.56704231e-07 0.0010887866 2.56804231e-07 -0.000993536867 2.56904231e-07 0.000907534878 2.57004231e-07 -0.000828173997
+ 2.57104231e-07 0.000756484035 2.57204231e-07 -0.000690353405 2.57304231e-07 0.000630593448 2.57404231e-07 -0.000575481614 2.57504231e-07 0.000525666393 2.57604231e-07 -0.000479733137 2.57704231e-07 0.000438207956 2.57804231e-07 -0.00039992149
+ 2.57904231e-07 0.000365307115 2.58004231e-07 -0.000333392049 2.58104231e-07 0.000304538809 2.58204231e-07 -0.000277932999 2.58304231e-07 0.000253882545 2.58404231e-07 -0.000231701277 2.58504231e-07 0.000211654724 2.58604231e-07 -0.000193160962
+ 2.58704231e-07 0.000176452339 2.58804231e-07 -0.000161031999 2.58904231e-07 0.000147106127 2.59004231e-07 -0.000134247508 2.59104231e-07 0.000122641562 2.59204231e-07 -0.000111918243 2.59304231e-07 0.000102246385 2.59404231e-07 -9.33029846e-05
+ 2.59504231e-07 8.52435523e-05 2.59604231e-07 -7.77838768e-05 2.59704231e-07 7.10687098e-05 2.59804231e-07 -6.4845882e-05 2.59904231e-07 5.925142e-05 2.60004231e-07 -5.40596605e-05 2.60104231e-07 4.93995251e-05 2.60204231e-07 -4.50673043e-05
+ 2.60304231e-07 4.11861142e-05 2.60404231e-07 -3.75704478e-05 2.60504231e-07 3.4338663e-05 2.60604231e-07 -3.13203588e-05 2.60704231e-07 2.86299828e-05 2.60804231e-07 -2.61096797e-05 2.60904231e-07 2.38706765e-05 2.61004231e-07 -2.17655435e-05
+ 2.61104231e-07 1.99028504e-05 2.61204231e-07 -1.81438359e-05 2.61304231e-07 1.65948732e-05 2.61404231e-07 -1.5124412e-05 2.61504231e-07 1.38370073e-05 2.61604231e-07 -1.26071091e-05 2.61704231e-07 1.15377661e-05 2.61804231e-07 -1.0508423e-05
+ 2.61904231e-07 9.62087887e-06 2.62004231e-07 -8.75873714e-06 2.62104231e-07 8.02275961e-06 2.62204231e-07 -7.3000129e-06 2.62304231e-07 6.69039716e-06 2.62404231e-07 -6.08386372e-06 2.62504231e-07 5.5795965e-06 2.62604231e-07 -5.06994997e-06
+ 2.62704231e-07 4.65351243e-06 2.62804231e-07 -4.22464061e-06 2.62904231e-07 3.88142724e-06 2.63004231e-07 -3.51989747e-06 2.63104231e-07 3.2377316e-06 2.63204231e-07 -2.93234513e-06 2.63304231e-07 2.70107501e-06 2.63404231e-07 -2.44249547e-06
+ 2.63504231e-07 2.25365756e-06 2.63604231e-07 -2.03410123e-06 2.63704231e-07 1.88063941e-06 2.63804231e-07 -1.693617e-06 2.63904231e-07 1.56964859e-06 2.64004231e-07 -1.40079315e-06 2.64104231e-07 1.32022001e-06 2.64204231e-07 -1.16494992e-06
+ 2.64304231e-07 1.10220937e-06 2.64404231e-07 -9.68844208e-07 2.64504231e-07 9.20524047e-07 2.64604231e-07 -8.05377434e-07 2.64704231e-07 7.69072859e-07 2.64804231e-07 -6.69112641e-07 2.64904231e-07 6.42823883e-07 2.65004231e-07 -5.55522921e-07
+ 2.65104231e-07 5.37583103e-07 2.65204231e-07 -4.60834721e-07 2.65304231e-07 4.49854148e-07 2.65404231e-07 -3.81902181e-07 2.65504231e-07 3.76722908e-07 2.65604231e-07 -3.16103905e-07 2.65704231e-07 3.15760619e-07 2.65804231e-07 -2.61254327e-07
+ 2.65904231e-07 2.64942218e-07 2.66004231e-07 -2.15531651e-07 2.66104231e-07 2.22580083e-07 2.66204231e-07 -1.77427235e-07 2.66304231e-07 1.87287055e-07 2.66404231e-07 -1.45682225e-07 2.66504231e-07 1.57884166e-07 2.66604231e-07 -1.192351e-07
+ 2.66704231e-07 1.33388171e-07 2.66804231e-07 -9.72014999e-08 2.66904231e-07 1.12980002e-07 2.67004231e-07 -7.8844731e-08 2.67104231e-07 9.59773834e-08 2.67204231e-07 -6.3551226e-08 2.67304231e-07 8.18121369e-08 2.67404231e-07 -5.07714672e-08
+ 2.67504231e-07 6.99716866e-08 2.67604231e-07 -4.01611717e-08 2.67704231e-07 6.01481946e-08 2.67804231e-07 -3.13254487e-08 2.67904231e-07 5.19644652e-08 2.68004231e-07 -2.3964328e-08 2.68104231e-07 4.51465265e-08 2.68204231e-07 -1.78317315e-08
+ 2.68304231e-07 3.94662536e-08 2.68404231e-07 -1.27220454e-08 2.68504231e-07 3.47335097e-08 2.68604231e-07 -8.46518614e-09 2.68704231e-07 3.07909064e-08 2.68804231e-07 -4.91900454e-09 2.68904231e-07 2.75064927e-08 2.69004231e-07 -1.96481095e-09
+ 2.69104231e-07 2.47703487e-08 2.69204231e-07 4.96254232e-10 2.69304231e-07 2.24974266e-08 2.69404231e-07 2.54098009e-09 2.69504231e-07 2.06303728e-08 2.69604231e-07 4.22158872e-09 2.69704231e-07 1.90956558e-08 2.69804231e-07 5.60309771e-09
+ 2.69904231e-07 1.78340379e-08 2.70004231e-07 6.73880085e-09 2.70104231e-07 1.67968681e-08 2.70204231e-07 7.6724801e-09 2.70304231e-07 1.59441737e-08 2.70404231e-07 8.44010861e-09 2.70504231e-07 1.5143805e-08 2.70604231e-07 9.05738082e-09
+ 2.70704231e-07 1.45796679e-08 2.70804231e-07 9.56953133e-09 2.70904231e-07 1.4115047e-08 2.71004231e-07 9.99100275e-09 2.71104231e-07 1.37327179e-08 2.71204231e-07 1.03378271e-08 2.71304231e-07 1.34180993e-08 2.71404231e-07 1.0623233e-08
+ 2.71504231e-07 1.31591912e-08 2.71604231e-07 1.08581061e-08 2.71704231e-07 1.29461198e-08 2.71804231e-07 1.10514014e-08 2.71904231e-07 1.27707626e-08 2.72004231e-07 1.12104871e-08 2.72104231e-07 1.26264374e-08 2.72204231e-07 1.13414238e-08
+ 2.72304231e-07 1.25076452e-08 2.72404231e-07 1.14491993e-08 2.72504231e-07 1.24098631e-08 2.72604231e-07 1.15379162e-08 2.72704231e-07 1.23293693e-08 2.72804231e-07 1.16109499e-08 2.72904231e-07 1.22631029e-08 2.73004231e-07 1.16710779e-08
+ 2.73104231e-07 1.22085438e-08 2.73204231e-07 1.17205853e-08 2.73304231e-07 1.21636195e-08 2.73404231e-07 1.17613514e-08 2.73504231e-07 1.2126625e-08 2.73604231e-07 1.17949243e-08 2.73704231e-07 1.20961568e-08 2.73804231e-07 1.18225761e-08
+ 2.73904231e-07 1.207106e-08 2.74004231e-07 1.18453544e-08 2.74104231e-07 1.2050385e-08 2.74204231e-07 1.18641207e-08 2.74304231e-07 1.20333504e-08 2.74404231e-07 1.18795845e-08 2.74504231e-07 1.20193125e-08 2.74604231e-07 1.18923288e-08
+ 2.74704231e-07 1.2007742e-08 2.74804231e-07 1.19028342e-08 2.74904231e-07 1.19982028e-08 2.75004231e-07 1.1911496e-08 2.75104231e-07 1.19903373e-08 2.75204231e-07 1.1918639e-08 2.75304231e-07 1.19838497e-08 2.75404231e-07 1.19245313e-08
+ 2.75504231e-07 1.19784974e-08 2.75604231e-07 1.19293936e-08 2.75704231e-07 1.19740802e-08 2.75804231e-07 1.19334069e-08 2.75904231e-07 1.19704341e-08 2.76004231e-07 1.19367206e-08 2.76104231e-07 1.19674221e-08 2.76204231e-07 1.19394577e-08
+ 2.76304231e-07 1.1964934e-08 2.76404231e-07 1.19417196e-08 2.76504231e-07 1.19628776e-08 2.76604231e-07 1.19435897e-08 2.76704231e-07 1.1961177e-08 2.76804231e-07 1.19451365e-08 2.76904231e-07 1.19597698e-08 2.77004231e-07 1.19464167e-08
+ 2.77104231e-07 1.19586049e-08 2.77204231e-07 1.19474767e-08 2.77304231e-07 1.19576401e-08 2.77404231e-07 1.19483551e-08 2.77504231e-07 1.195684e-08 2.77604231e-07 1.19490836e-08 2.77704231e-07 1.19561769e-08 2.77804231e-07 1.1949688e-08
+ 2.77904231e-07 1.1955626e-08 2.78004231e-07 1.19501899e-08 2.78104231e-07 1.19551683e-08 2.78204231e-07 1.19506073e-08 2.78304231e-07 1.19547877e-08 2.78404231e-07 1.19509548e-08 2.78504231e-07 1.19544707e-08 2.78604231e-07 1.19512439e-08
+ 2.78704231e-07 1.19542066e-08 2.78804231e-07 1.19514852e-08 2.78904231e-07 1.19539862e-08 2.79004231e-07 1.19516868e-08 2.79104231e-07 1.19538021e-08 2.79204231e-07 1.19518552e-08 2.79304231e-07 1.19536476e-08 2.79404231e-07 1.19519965e-08
+ 2.79504231e-07 1.19535187e-08 2.79604231e-07 1.19521147e-08 2.79704231e-07 1.19534104e-08 2.79804231e-07 1.19522138e-08 2.79904231e-07 1.19533192e-08 2.80004231e-07 1.19522975e-08 2.80104231e-07 1.19532425e-08 2.80204231e-07 1.19523678e-08
+ 2.80304231e-07 1.19531779e-08 2.80404231e-07 1.19524269e-08 2.80504231e-07 1.19531235e-08 2.80604231e-07 1.19524772e-08 2.80704231e-07 1.19530773e-08 2.80804231e-07 1.19525197e-08 2.80904231e-07 1.1953038e-08 2.81004231e-07 1.1952556e-08
+ 2.81104231e-07 1.19530047e-08 2.81204231e-07 1.19525866e-08 2.81304231e-07 1.19529763e-08 2.81404231e-07 1.19526131e-08 2.81504231e-07 1.19529517e-08 2.81604231e-07 1.19526358e-08 2.81704231e-07 1.1952931e-08 2.81804231e-07 1.1952655e-08
+ 2.81904231e-07 1.19529131e-08 2.82004231e-07 1.19526714e-08 2.82104231e-07 1.19528978e-08 2.82204231e-07 1.1952686e-08 2.82304231e-07 1.19528844e-08 2.82404231e-07 1.19526981e-08 2.82504231e-07 1.19528729e-08 2.82604231e-07 1.19527088e-08
+ 2.82704231e-07 1.19528631e-08 2.82804231e-07 1.19527178e-08 2.82904231e-07 1.19528545e-08 2.83004231e-07 1.19527263e-08 2.83104231e-07 1.1952847e-08 2.83204231e-07 1.1952733e-08 2.83304231e-07 1.19528403e-08 2.83404231e-07 1.19527395e-08
+ 2.83504231e-07 1.19528344e-08 2.83604231e-07 1.19527449e-08 2.83704231e-07 1.19528294e-08 2.83804231e-07 1.19527495e-08 2.83904231e-07 1.19528249e-08 2.84004231e-07 1.19527536e-08 2.84104231e-07 1.19528211e-08 2.84204231e-07 1.19527573e-08
+ 2.84304231e-07 1.19528177e-08 2.84404231e-07 1.19527606e-08 2.84504231e-07 1.19528145e-08 2.84604231e-07 1.19527635e-08 2.84704231e-07 1.19528117e-08 2.84804231e-07 1.19527657e-08 2.84904231e-07 1.19528095e-08 2.85004231e-07 1.19527683e-08
+ 2.85104231e-07 1.19528072e-08 2.85204231e-07 1.19527703e-08 2.85304231e-07 1.19528052e-08 2.85404231e-07 1.19527721e-08 2.85504231e-07 1.19528035e-08 2.85604231e-07 1.19527738e-08 2.85704231e-07 1.19528021e-08 2.85804231e-07 1.19527751e-08
+ 2.85904231e-07 1.19528009e-08 2.86004231e-07 1.19527765e-08 2.86104231e-07 1.19527997e-08 2.86204231e-07 1.19527773e-08 2.86304231e-07 1.19527987e-08 2.86404231e-07 1.19527784e-08 2.86504231e-07 1.19527977e-08 2.86604231e-07 1.19527794e-08
+ 2.86704231e-07 1.19527966e-08 2.86804231e-07 1.19527806e-08 2.86904231e-07 1.19527958e-08 2.87004231e-07 1.19527814e-08 2.87104231e-07 1.19527951e-08 2.87204231e-07 1.19527819e-08 2.87304231e-07 1.19527943e-08 2.87404231e-07 1.19527826e-08
+ 2.87504231e-07 1.19527936e-08 2.87604231e-07 1.1952783e-08 2.87704231e-07 1.19527933e-08 2.87804231e-07 1.19527834e-08 2.87904231e-07 1.19527929e-08 2.88004231e-07 1.19527841e-08 2.88104231e-07 1.19527924e-08 2.88204231e-07 1.19527845e-08
+ 2.88304231e-07 1.1952792e-08 2.88404231e-07 1.19527848e-08 2.88504231e-07 1.19527917e-08 2.88604231e-07 1.19527852e-08 2.88704231e-07 1.19527913e-08 2.88804231e-07 1.19527855e-08 2.88904231e-07 1.19527908e-08 2.89004231e-07 1.19527858e-08
+ 2.89104231e-07 1.19527908e-08 2.89204231e-07 1.1952786e-08 2.89304231e-07 1.19527906e-08 2.89404231e-07 1.19527863e-08 2.89504231e-07 1.19527901e-08 2.89604231e-07 1.19527866e-08 2.89704231e-07 1.19527899e-08 2.89804231e-07 1.19527868e-08
+ 2.89904231e-07 1.19527897e-08 2.90004231e-07 1.19527867e-08 2.90104231e-07 1.19527899e-08 2.90204231e-07 1.19527871e-08 2.90304231e-07 1.19527895e-08 2.90404231e-07 1.19527871e-08 2.90504231e-07 1.19527894e-08 2.90604231e-07 1.19527871e-08
+ 2.90704231e-07 1.19527896e-08 2.90804231e-07 1.19527871e-08 2.90904231e-07 1.19527895e-08 2.91004231e-07 1.19527873e-08 2.91104231e-07 1.19527895e-08 2.91204231e-07 1.19527873e-08 2.91304231e-07 1.19527894e-08 2.91404231e-07 1.19527874e-08
+ 2.91504231e-07 1.19527894e-08 2.91604231e-07 1.19527873e-08 2.91704231e-07 1.19527892e-08 2.91804231e-07 1.19527874e-08 2.91904231e-07 1.19527894e-08 2.92004231e-07 1.19527874e-08 2.92104231e-07 1.19527893e-08 2.92204231e-07 1.19527875e-08
+ 2.92304231e-07 1.19527892e-08 2.92404231e-07 1.19527875e-08 2.92504231e-07 1.19527891e-08 2.92604231e-07 1.19527877e-08 2.92704231e-07 1.1952789e-08 2.92804231e-07 1.19527878e-08 2.92904231e-07 1.1952789e-08 2.93004231e-07 1.19527878e-08
+ 2.93104231e-07 1.19527889e-08 2.93204231e-07 1.19527879e-08 2.93304231e-07 1.1952789e-08 2.93404231e-07 1.19527879e-08 2.93504231e-07 1.19527889e-08 2.93604231e-07 1.1952788e-08 2.93704231e-07 1.19527889e-08 2.93804231e-07 1.19527879e-08
+ 2.93904231e-07 1.19527888e-08 2.94004231e-07 1.1952788e-08 2.94104231e-07 1.19527889e-08 2.94204231e-07 1.1952788e-08 2.94304231e-07 1.19527888e-08 2.94404231e-07 1.1952788e-08 2.94504231e-07 1.19527888e-08 2.94604231e-07 1.1952788e-08
+ 2.94704231e-07 1.19527888e-08 2.94804231e-07 1.19527881e-08 2.94904231e-07 1.19527888e-08 2.95004231e-07 1.19527881e-08 2.95104231e-07 1.19527886e-08 2.95204231e-07 1.1952788e-08 2.95304231e-07 1.19527887e-08 2.95404231e-07 1.19527881e-08
+ 2.95504231e-07 1.19527886e-08 2.95604231e-07 1.19527881e-08 2.95704231e-07 1.19527886e-08 2.95804231e-07 1.19527881e-08 2.95904231e-07 1.19527887e-08 2.96004231e-07 1.19527881e-08 2.96104231e-07 1.19527886e-08 2.96204231e-07 1.19527881e-08
+ 2.96304231e-07 1.19527887e-08 2.96404231e-07 1.19527881e-08 2.96504231e-07 1.19527885e-08 2.96604231e-07 1.1952788e-08 2.96704231e-07 1.19527887e-08 2.96804231e-07 1.19527881e-08 2.96904231e-07 1.19527886e-08 2.97004231e-07 1.19527882e-08
+ 2.97104231e-07 1.19527886e-08 2.97204231e-07 1.19527883e-08 2.97304231e-07 1.19527884e-08 2.97404231e-07 1.19527883e-08 2.97504231e-07 1.19527885e-08 2.97604231e-07 1.19527883e-08 2.97704231e-07 1.19527885e-08 2.97804231e-07 1.19527883e-08
+ 2.97904231e-07 1.19527885e-08 2.98004231e-07 1.19527883e-08 2.98104231e-07 1.19527885e-08 2.98204231e-07 1.19527883e-08 2.98304231e-07 1.19527885e-08 2.98404231e-07 1.19527883e-08 2.98504231e-07 1.19527884e-08 2.98604231e-07 1.19527883e-08
+ 2.98704231e-07 1.19527885e-08 2.98804231e-07 1.19527883e-08 2.98904231e-07 1.19527885e-08 2.99004231e-07 1.19527883e-08 2.99104231e-07 1.19527885e-08 2.99204231e-07 1.19527883e-08 2.99304231e-07 1.19527885e-08 2.99404231e-07 1.19527883e-08
+ 2.99504231e-07 1.19527885e-08 2.99604231e-07 1.19527883e-08 2.99704231e-07 1.19527885e-08 2.99804231e-07 1.19527883e-08 2.99904231e-07 1.19527885e-08 3e-07 1.19527882e-08 3.0001e-07 1.45267508e-08 3.0003e-07 1.23970101e-09
+ 3.0007e-07 2.76375266e-08 3.0015e-07 -4.37848929e-09 3.0025e-07 2.82049111e-08 3.0035e-07 -3.17728022e-09 3.0045e-07 2.52046194e-08 3.0055e-07 2.60783994e-09 3.0065e-07 -4.06484911e-08 3.0075e-07 3.06912282e-06
+ 3.0085e-07 9.51416557e-05 3.00931988e-07 -0.0447690188 3.01e-07 1.97565125 3.01008484e-07 3.09900368 3.01025451e-07 4.14251596 3.01059385e-07 4.88272691 3.01090588e-07 4.97988863 3.01143428e-07 5.00280497
+ 3.011991e-07 4.99920014 3.012991e-07 5.00046356 3.013991e-07 4.99971393 3.014991e-07 5.00018225 3.01578678e-07 4.99989094 3.01663998e-07 5.00006899 3.01763998e-07 4.99995201 3.01858547e-07 5.00003258
+ 3.01958547e-07 4.99997704 3.02058547e-07 5.00001602 3.02158547e-07 4.99998864 3.02258547e-07 5.00000791 3.02358547e-07 4.99999437 3.02458547e-07 5.00000389 3.02558547e-07 4.99999721 3.02658547e-07 5.0000019
+ 3.02758547e-07 4.99999862 3.02858547e-07 5.00000091 3.02958547e-07 4.99999932 3.03058547e-07 5.00000042 3.03158547e-07 4.99999966 3.03258547e-07 5.00000018 3.03358547e-07 4.99999983 3.03458547e-07 5.00000007
+ 3.03558547e-07 4.99999991 3.03658547e-07 5.00000001 3.03758547e-07 4.99999995 3.03858547e-07 4.99999999 3.03958547e-07 4.99999996 3.04058547e-07 4.99999998 3.04158547e-07 4.99999997 3.04258547e-07 4.99999997
+ 3.04358547e-07 4.99999997 3.04458547e-07 4.99999997 3.04558547e-07 4.99999997 3.04658547e-07 4.99999997 3.04758547e-07 4.99999997 3.04858547e-07 4.99999997 3.04958547e-07 4.99999997 3.05058547e-07 4.99999997
+ 3.05158547e-07 4.99999997 3.05258547e-07 4.99999997 3.05358547e-07 4.99999997 3.05458547e-07 4.99999997 3.05558547e-07 4.99999997 3.05658547e-07 4.99999997 3.05758547e-07 4.99999997 3.05858547e-07 4.99999997
+ 3.05958547e-07 4.99999997 3.06058547e-07 4.99999997 3.06158547e-07 4.99999997 3.06258547e-07 4.99999997 3.06358547e-07 4.99999997 3.06458547e-07 4.99999997 3.06558547e-07 4.99999997 3.06658547e-07 4.99999997
+ 3.06758547e-07 4.99999997 3.06858547e-07 4.99999997 3.06958547e-07 4.99999997 3.07058547e-07 4.99999997 3.07158547e-07 4.99999997 3.07258547e-07 4.99999997 3.07358547e-07 4.99999997 3.07458547e-07 4.99999997
+ 3.07558547e-07 4.99999997 3.07658547e-07 4.99999997 3.07758547e-07 4.99999997 3.07858547e-07 4.99999997 3.07958547e-07 4.99999997 3.08058547e-07 4.99999997 3.08158547e-07 4.99999997 3.08258547e-07 4.99999997
+ 3.08358547e-07 4.99999997 3.08458547e-07 4.99999997 3.08558547e-07 4.99999997 3.08658547e-07 4.99999997 3.08758547e-07 4.99999997 3.08858547e-07 4.99999997 3.08958547e-07 4.99999997 3.09058547e-07 4.99999997
+ 3.09158547e-07 4.99999997 3.09258547e-07 4.99999997 3.09358547e-07 4.99999997 3.09458547e-07 4.99999997 3.09558547e-07 4.99999997 3.09658547e-07 4.99999997 3.09758547e-07 4.99999997 3.09858547e-07 4.99999997
+ 3.09958547e-07 4.99999997 3.10058547e-07 4.99999997 3.10158547e-07 4.99999997 3.10258547e-07 4.99999997 3.10358547e-07 4.99999997 3.10458547e-07 4.99999997 3.10558547e-07 4.99999997 3.10658547e-07 4.99999997
+ 3.10758547e-07 4.99999997 3.10858547e-07 4.99999997 3.10958547e-07 4.99999997 3.11058547e-07 4.99999997 3.11158547e-07 4.99999997 3.11258547e-07 4.99999997 3.11358547e-07 4.99999997 3.11458547e-07 4.99999997
+ 3.11558547e-07 4.99999997 3.11658547e-07 4.99999997 3.11758547e-07 4.99999997 3.11858547e-07 4.99999997 3.11958547e-07 4.99999997 3.12058547e-07 4.99999997 3.12158547e-07 4.99999997 3.12258547e-07 4.99999997
+ 3.12358547e-07 4.99999997 3.12458547e-07 4.99999997 3.12558547e-07 4.99999997 3.12658547e-07 4.99999997 3.12758547e-07 4.99999997 3.12858547e-07 4.99999997 3.12958547e-07 4.99999997 3.13058547e-07 4.99999997
+ 3.13158547e-07 4.99999997 3.13258547e-07 4.99999997 3.13358547e-07 4.99999997 3.13458547e-07 4.99999997 3.13558547e-07 4.99999997 3.13658547e-07 4.99999997 3.13758547e-07 4.99999997 3.13858547e-07 4.99999997
+ 3.13958547e-07 4.99999997 3.14058547e-07 4.99999997 3.14158547e-07 4.99999997 3.14258547e-07 4.99999997 3.14358547e-07 4.99999997 3.14458547e-07 4.99999997 3.14558547e-07 4.99999997 3.14658547e-07 4.99999997
+ 3.14758547e-07 4.99999997 3.14858547e-07 4.99999997 3.14958547e-07 4.99999997 3.15058547e-07 4.99999997 3.15158547e-07 4.99999997 3.15258547e-07 4.99999997 3.15358547e-07 4.99999997 3.15458547e-07 4.99999997
+ 3.15558547e-07 4.99999997 3.15658547e-07 4.99999997 3.15758547e-07 4.99999997 3.15858547e-07 4.99999997 3.15958547e-07 4.99999997 3.16058547e-07 4.99999997 3.16158547e-07 4.99999997 3.16258547e-07 4.99999997
+ 3.16358547e-07 4.99999997 3.16458547e-07 4.99999997 3.16558547e-07 4.99999997 3.16658547e-07 4.99999997 3.16758547e-07 4.99999997 3.16858547e-07 4.99999997 3.16958547e-07 4.99999997 3.17058547e-07 4.99999997
+ 3.17158547e-07 4.99999997 3.17258547e-07 4.99999997 3.17358547e-07 4.99999997 3.17458547e-07 4.99999997 3.17558547e-07 4.99999997 3.17658547e-07 4.99999997 3.17758547e-07 4.99999997 3.17858547e-07 4.99999997
+ 3.17958547e-07 4.99999997 3.18058547e-07 4.99999997 3.18158547e-07 4.99999997 3.18258547e-07 4.99999997 3.18358547e-07 4.99999997 3.18458547e-07 4.99999997 3.18558547e-07 4.99999997 3.18658547e-07 4.99999997
+ 3.18758547e-07 4.99999997 3.18858547e-07 4.99999997 3.18958547e-07 4.99999997 3.19058547e-07 4.99999997 3.19158547e-07 4.99999997 3.19258547e-07 4.99999997 3.19358547e-07 4.99999997 3.19458547e-07 4.99999997
+ 3.19558547e-07 4.99999997 3.19658547e-07 4.99999997 3.19758547e-07 4.99999997 3.19858547e-07 4.99999997 3.19958547e-07 4.99999997 3.20058547e-07 4.99999997 3.20158547e-07 4.99999997 3.20258547e-07 4.99999997
+ 3.20358547e-07 4.99999997 3.20458547e-07 4.99999997 3.20558547e-07 4.99999997 3.20658547e-07 4.99999997 3.20758547e-07 4.99999997 3.20858547e-07 4.99999997 3.20958547e-07 4.99999997 3.21058547e-07 4.99999997
+ 3.21158547e-07 4.99999997 3.21258547e-07 4.99999997 3.21358547e-07 4.99999997 3.21458547e-07 4.99999997 3.21558547e-07 4.99999997 3.21658547e-07 4.99999997 3.21758547e-07 4.99999997 3.21858547e-07 4.99999997
+ 3.21958547e-07 4.99999997 3.22058547e-07 4.99999997 3.22158547e-07 4.99999997 3.22258547e-07 4.99999997 3.22358547e-07 4.99999997 3.22458547e-07 4.99999997 3.22558547e-07 4.99999997 3.22658547e-07 4.99999997
+ 3.22758547e-07 4.99999997 3.22858547e-07 4.99999997 3.22958547e-07 4.99999997 3.23058547e-07 4.99999997 3.23158547e-07 4.99999997 3.23258547e-07 4.99999997 3.23358547e-07 4.99999997 3.23458547e-07 4.99999997
+ 3.23558547e-07 4.99999997 3.23658547e-07 4.99999997 3.23758547e-07 4.99999997 3.23858547e-07 4.99999997 3.23958547e-07 4.99999997 3.24058547e-07 4.99999997 3.24158547e-07 4.99999997 3.24258547e-07 4.99999997
+ 3.24358547e-07 4.99999997 3.24458547e-07 4.99999997 3.24558547e-07 4.99999997 3.24658547e-07 4.99999997 3.24758547e-07 4.99999997 3.24858547e-07 4.99999997 3.24958547e-07 4.99999997 3.25058547e-07 4.99999997
+ 3.25158547e-07 4.99999997 3.25258547e-07 4.99999997 3.25358547e-07 4.99999997 3.25458547e-07 4.99999997 3.25558547e-07 4.99999997 3.25658547e-07 4.99999997 3.25758547e-07 4.99999997 3.25858547e-07 4.99999997
+ 3.25958547e-07 4.99999997 3.26058547e-07 4.99999997 3.26158547e-07 4.99999997 3.26258547e-07 4.99999997 3.26358547e-07 4.99999997 3.26458547e-07 4.99999997 3.26558547e-07 4.99999997 3.26658547e-07 4.99999997
+ 3.26758547e-07 4.99999997 3.26858547e-07 4.99999997 3.26958547e-07 4.99999997 3.27058547e-07 4.99999997 3.27158547e-07 4.99999997 3.27258547e-07 4.99999997 3.27358547e-07 4.99999997 3.27458547e-07 4.99999997
+ 3.27558547e-07 4.99999997 3.27658547e-07 4.99999997 3.27758547e-07 4.99999997 3.27858547e-07 4.99999997 3.27958547e-07 4.99999997 3.28058547e-07 4.99999997 3.28158547e-07 4.99999997 3.28258547e-07 4.99999997
+ 3.28358547e-07 4.99999997 3.28458547e-07 4.99999997 3.28558547e-07 4.99999997 3.28658547e-07 4.99999997 3.28758547e-07 4.99999997 3.28858547e-07 4.99999997 3.28958547e-07 4.99999997 3.29058547e-07 4.99999997
+ 3.29158547e-07 4.99999997 3.29258547e-07 4.99999997 3.29358547e-07 4.99999997 3.29458547e-07 4.99999997 3.29558547e-07 4.99999997 3.29658547e-07 4.99999997 3.29758547e-07 4.99999997 3.29858547e-07 4.99999997
+ 3.29958547e-07 4.99999997 3.30058547e-07 4.99999997 3.30158547e-07 4.99999997 3.30258547e-07 4.99999997 3.30358547e-07 4.99999997 3.30458547e-07 4.99999997 3.30558547e-07 4.99999997 3.30658547e-07 4.99999997
+ 3.30758547e-07 4.99999997 3.30858547e-07 4.99999997 3.30958547e-07 4.99999997 3.31058547e-07 4.99999997 3.31158547e-07 4.99999997 3.31258547e-07 4.99999997 3.31358547e-07 4.99999997 3.31458547e-07 4.99999997
+ 3.31558547e-07 4.99999997 3.31658547e-07 4.99999997 3.31758547e-07 4.99999997 3.31858547e-07 4.99999997 3.31958547e-07 4.99999997 3.32058547e-07 4.99999997 3.32158547e-07 4.99999997 3.32258547e-07 4.99999997
+ 3.32358547e-07 4.99999997 3.32458547e-07 4.99999997 3.32558547e-07 4.99999997 3.32658547e-07 4.99999997 3.32758547e-07 4.99999997 3.32858547e-07 4.99999997 3.32958547e-07 4.99999997 3.33058547e-07 4.99999997
+ 3.33158547e-07 4.99999997 3.33258547e-07 4.99999997 3.33358547e-07 4.99999997 3.33458547e-07 4.99999997 3.33558547e-07 4.99999997 3.33658547e-07 4.99999997 3.33758547e-07 4.99999997 3.33858547e-07 4.99999997
+ 3.33958547e-07 4.99999997 3.34058547e-07 4.99999997 3.34158547e-07 4.99999997 3.34258547e-07 4.99999997 3.34358547e-07 4.99999997 3.34458547e-07 4.99999997 3.34558547e-07 4.99999997 3.34658547e-07 4.99999997
+ 3.34758547e-07 4.99999997 3.34858547e-07 4.99999997 3.34958547e-07 4.99999997 3.35058547e-07 4.99999997 3.35158547e-07 4.99999997 3.35258547e-07 4.99999997 3.35358547e-07 4.99999997 3.35458547e-07 4.99999997
+ 3.35558547e-07 4.99999997 3.35658547e-07 4.99999997 3.35758547e-07 4.99999997 3.35858547e-07 4.99999997 3.35958547e-07 4.99999997 3.36058547e-07 4.99999997 3.36158547e-07 4.99999997 3.36258547e-07 4.99999997
+ 3.36358547e-07 4.99999997 3.36458547e-07 4.99999997 3.36558547e-07 4.99999997 3.36658547e-07 4.99999997 3.36758547e-07 4.99999997 3.36858547e-07 4.99999997 3.36958547e-07 4.99999997 3.37058547e-07 4.99999997
+ 3.37158547e-07 4.99999997 3.37258547e-07 4.99999997 3.37358547e-07 4.99999997 3.37458547e-07 4.99999997 3.37558547e-07 4.99999997 3.37658547e-07 4.99999997 3.37758547e-07 4.99999997 3.37858547e-07 4.99999997
+ 3.37958547e-07 4.99999997 3.38058547e-07 4.99999997 3.38158547e-07 4.99999997 3.38258547e-07 4.99999997 3.38358547e-07 4.99999997 3.38458547e-07 4.99999997 3.38558547e-07 4.99999997 3.38658547e-07 4.99999997
+ 3.38758547e-07 4.99999997 3.38858547e-07 4.99999997 3.38958547e-07 4.99999997 3.39058547e-07 4.99999997 3.39158547e-07 4.99999997 3.39258547e-07 4.99999997 3.39358547e-07 4.99999997 3.39458547e-07 4.99999997
+ 3.39558547e-07 4.99999997 3.39658547e-07 4.99999997 3.39758547e-07 4.99999997 3.39858547e-07 4.99999997 3.39958547e-07 4.99999997 3.40058547e-07 4.99999997 3.40158547e-07 4.99999997 3.40258547e-07 4.99999997
+ 3.40358547e-07 4.99999997 3.40458547e-07 4.99999997 3.40558547e-07 4.99999997 3.40658547e-07 4.99999997 3.40758547e-07 4.99999997 3.40858547e-07 4.99999997 3.40958547e-07 4.99999997 3.41058547e-07 4.99999997
+ 3.41158547e-07 4.99999997 3.41258547e-07 4.99999997 3.41358547e-07 4.99999997 3.41458547e-07 4.99999997 3.41558547e-07 4.99999997 3.41658547e-07 4.99999997 3.41758547e-07 4.99999997 3.41858547e-07 4.99999997
+ 3.41958547e-07 4.99999997 3.42058547e-07 4.99999997 3.42158547e-07 4.99999997 3.42258547e-07 4.99999997 3.42358547e-07 4.99999997 3.42458547e-07 4.99999997 3.42558547e-07 4.99999997 3.42658547e-07 4.99999997
+ 3.42758547e-07 4.99999997 3.42858547e-07 4.99999997 3.42958547e-07 4.99999997 3.43058547e-07 4.99999997 3.43158547e-07 4.99999997 3.43258547e-07 4.99999997 3.43358547e-07 4.99999997 3.43458547e-07 4.99999997
+ 3.43558547e-07 4.99999997 3.43658547e-07 4.99999997 3.43758547e-07 4.99999997 3.43858547e-07 4.99999997 3.43958547e-07 4.99999997 3.44058547e-07 4.99999997 3.44158547e-07 4.99999997 3.44258547e-07 4.99999997
+ 3.44358547e-07 4.99999997 3.44458547e-07 4.99999997 3.44558547e-07 4.99999997 3.44658547e-07 4.99999997 3.44758547e-07 4.99999997 3.44858547e-07 4.99999997 3.44958547e-07 4.99999997 3.45058547e-07 4.99999997
+ 3.45158547e-07 4.99999997 3.45258547e-07 4.99999997 3.45358547e-07 4.99999997 3.45458547e-07 4.99999997 3.45558547e-07 4.99999997 3.45658547e-07 4.99999997 3.45758547e-07 4.99999997 3.45858547e-07 4.99999997
+ 3.45958547e-07 4.99999997 3.46058547e-07 4.99999997 3.46158547e-07 4.99999997 3.46258547e-07 4.99999997 3.46358547e-07 4.99999997 3.46458547e-07 4.99999997 3.46558547e-07 4.99999997 3.46658547e-07 4.99999997
+ 3.46758547e-07 4.99999997 3.46858547e-07 4.99999997 3.46958547e-07 4.99999997 3.47058547e-07 4.99999997 3.47158547e-07 4.99999997 3.47258547e-07 4.99999997 3.47358547e-07 4.99999997 3.47458547e-07 4.99999997
+ 3.47558547e-07 4.99999997 3.47658547e-07 4.99999997 3.47758547e-07 4.99999997 3.47858547e-07 4.99999997 3.47958547e-07 4.99999997 3.48058547e-07 4.99999997 3.48158547e-07 4.99999997 3.48258547e-07 4.99999997
+ 3.48358547e-07 4.99999997 3.48458547e-07 4.99999997 3.48558547e-07 4.99999997 3.48658547e-07 4.99999997 3.48758547e-07 4.99999997 3.48858547e-07 4.99999997 3.48958547e-07 4.99999997 3.49058547e-07 4.99999997
+ 3.49158547e-07 4.99999997 3.49258547e-07 4.99999997 3.49358547e-07 4.99999997 3.49458547e-07 4.99999997 3.49558547e-07 4.99999997 3.49658547e-07 4.99999997 3.49758547e-07 4.99999997 3.49858547e-07 4.99999997
+ 3.49958547e-07 4.99999997 3.50058547e-07 4.99999997 3.50158547e-07 4.99999997 3.50258547e-07 4.99999997 3.50358547e-07 4.99999997 3.50458547e-07 4.99999997 3.50558547e-07 4.99999997 3.50658547e-07 4.99999997
+ 3.50758547e-07 4.99999997 3.50858547e-07 4.99999997 3.50958547e-07 4.99999997 3.51e-07 4.99999997 3.5101e-07 4.99999997 3.5103e-07 4.99999998 3.5107e-07 4.99999996 3.5115e-07 4.99999998
+ 3.5125e-07 4.99999997 3.5135e-07 4.99999997 3.5145e-07 4.99999998 3.5155e-07 4.99999996 3.5165e-07 4.99999998 3.5175e-07 4.99999996 3.5185e-07 4.99999999 3.51930828e-07 5.00006471
+ 3.52e-07 4.99916173 3.52008608e-07 4.99761842 3.52025825e-07 4.99312391 3.52060258e-07 5.01021642 3.52106188e-07 5.09915302 3.52150118e-07 4.2138351 3.5219811e-07 0.290132927 3.522555e-07 -0.055559802
+ 3.52312176e-07 0.0719919946 3.52404431e-07 -0.0580528341 3.52490759e-07 0.0521271683 3.52590759e-07 -0.0468986726 3.52690759e-07 0.0429726694 3.52790759e-07 -0.0387916891 3.52890759e-07 0.0355067968 3.52990759e-07 -0.0321238152
+ 3.53090759e-07 0.0293826519 3.53190759e-07 -0.0266208089 3.53290759e-07 0.0243463628 3.53390759e-07 -0.0220869282 3.53490759e-07 0.0201946558 3.53590759e-07 -0.018340188 3.53690759e-07 0.0167656294 3.53790759e-07 -0.0152394344
+ 3.53890759e-07 0.0139289603 3.53990759e-07 -0.0126701333 3.54090759e-07 0.0115791999 3.54190759e-07 -0.0105389933 3.54290759e-07 0.00963062169 3.54390759e-07 -0.00876976083 3.54490759e-07 0.00801325014 3.54590759e-07 -0.00729991652
+ 3.54690759e-07 0.00666976939 3.54790759e-07 -0.00607806441 3.54890759e-07 0.00555309574 3.54990759e-07 -0.00506185631 3.55090759e-07 0.00462445582 3.55190759e-07 -0.00421633125 3.55290759e-07 0.00385185386 3.55390759e-07 -0.00351257961
+ 3.55490759e-07 0.00320884134 3.55590759e-07 -0.00292666284 3.55690759e-07 0.00267352374 3.55790759e-07 -0.00243873589 3.55890759e-07 0.00222775459 3.55990759e-07 -0.00203233144 3.56090759e-07 0.00185647883 3.56190759e-07 -0.00169377401
+ 3.56290759e-07 0.00154719576 3.56390759e-07 -0.00141169917 3.56490759e-07 0.00128951848 3.56590759e-07 -0.00117744179 3.56690759e-07 0.00107519826 3.56790759e-07 -0.000980224982 3.56890759e-07 0.000896201859 3.56990759e-07 -0.000816256475
+ 3.57090759e-07 0.000747091622 3.57190759e-07 -0.000679905625 3.57290759e-07 0.000622853518 3.57390759e-07 -0.000568158092 3.57490759e-07 0.000518950145 3.57590759e-07 -0.000473602727 3.57690759e-07 0.000432609181 3.57790759e-07 -0.000394813042
+ 3.57890759e-07 0.000360641794 3.57990759e-07 -0.00032913503 3.58090759e-07 0.000300650957 3.58190759e-07 -0.000274385188 3.58290759e-07 0.000250642317 3.58390759e-07 -0.000227597045 3.58490759e-07 0.000209143757 3.58590759e-07 -0.000189777838
+ 3.58690759e-07 0.000174428486 3.58790759e-07 -0.000158243287 3.58890759e-07 0.000146480534 3.58990759e-07 -0.000131798715 3.59090759e-07 0.000122072762 3.59190759e-07 -0.000109833166 3.59290759e-07 0.000101741072 3.59390759e-07 -9.15328229e-05
+ 3.59490759e-07 8.4798664e-05 3.59590759e-07 -7.62841394e-05 3.59690759e-07 7.06796878e-05 3.59790759e-07 -6.3577359e-05 3.59890759e-07 5.89130619e-05 3.59990759e-07 -5.29881514e-05 3.60090759e-07 4.91064763e-05 3.60190759e-07 -4.41632069e-05
+ 3.60290759e-07 4.09331671e-05 3.60390759e-07 -3.68082931e-05 3.60490759e-07 3.41209287e-05 3.60590759e-07 -3.06783363e-05 3.60690759e-07 2.84429787e-05 3.60790759e-07 -2.55691818e-05 3.60890759e-07 2.37103609e-05 3.60990759e-07 -2.13107424e-05
+ 3.61090759e-07 1.97656238e-05 3.61190759e-07 -1.77613005e-05 3.61290759e-07 1.64775595e-05 3.61390759e-07 -1.48027673e-05 3.61490759e-07 1.37368234e-05 3.61590759e-07 -1.23367368e-05 3.61690759e-07 1.14522874e-05 3.61790759e-07 -1.02812005e-05
+ 3.61890759e-07 9.54800221e-06 3.61990759e-07 -8.56781254e-06 3.62090759e-07 7.96066694e-06 3.62190759e-07 -7.13961088e-06 3.62290759e-07 6.63752161e-06 3.62390759e-07 -5.94912011e-06 3.62490759e-07 5.5345908e-06 3.62590759e-07 -4.95677035e-06
+ 3.62690759e-07 4.61522039e-06 3.62790759e-07 -4.1295802e-06 3.62890759e-07 3.84885826e-06 3.62990759e-07 -3.44005922e-06 3.63090759e-07 3.21003811e-06 3.63190759e-07 -2.86529346e-06 3.63290759e-07 2.67753269e-06 3.63390759e-07 -2.38618332e-06
+ 3.63490759e-07 2.23364797e-06 3.63590759e-07 -1.98680848e-06 3.63690759e-07 1.86363501e-06 3.63790759e-07 -1.65389859e-06 3.63890759e-07 1.55519979e-06 3.63990759e-07 -1.37639223e-06 3.64090759e-07 1.29809458e-06 3.64190759e-07 -1.14506907e-06
+ 3.64290759e-07 1.08377708e-06 3.64390759e-07 -9.52243233e-07 3.64490759e-07 9.05126584e-07 3.64590759e-07 -7.91507923e-07 3.64690759e-07 7.56207395e-07 3.64790759e-07 -6.57522578e-07 3.64890759e-07 6.32071612e-07 3.64990759e-07 -5.4583533e-07
+ 3.65090759e-07 5.28594424e-07 3.65190759e-07 -4.52734886e-07 3.65290759e-07 4.42337866e-07 3.65390759e-07 -3.7512853e-07 3.65490759e-07 3.70436519e-07 3.65590759e-07 -3.10437819e-07 3.65690759e-07 3.10501328e-07 3.65790759e-07 -2.56513247e-07
+ 3.65890759e-07 2.60540816e-07 3.65990759e-07 -2.11564428e-07 3.66090759e-07 2.18897721e-07 3.66190759e-07 -1.74107636e-07 3.66290759e-07 1.84205258e-07 3.66390759e-07 -1.42903498e-07 3.66490759e-07 1.55303991e-07 3.66590759e-07 -1.16908189e-07
+ 3.66690759e-07 1.31227074e-07 3.66790759e-07 -9.52521049e-08 3.66890759e-07 1.11169114e-07 3.66990759e-07 -7.72108563e-08 3.67090759e-07 9.44592506e-08 3.67190759e-07 -6.21811994e-08 3.67290759e-07 8.05388985e-08 3.67390759e-07 -4.96223675e-08
+ 3.67490759e-07 6.89035346e-08 3.67590759e-07 -3.91967472e-08 3.67690759e-07 5.92514597e-08 3.67790759e-07 -3.05155714e-08 3.67890759e-07 5.12112143e-08 3.67990759e-07 -2.32838318e-08 3.68090759e-07 4.45134132e-08 3.68190759e-07 -1.72595827e-08
+ 3.68290759e-07 3.8933772e-08 3.68390759e-07 -1.22406799e-08 3.68490759e-07 3.42853601e-08 3.68590759e-07 -8.05990238e-09 3.68690759e-07 3.04134395e-08 3.68790759e-07 -4.57750141e-09 3.68890759e-07 2.7188293e-08 3.68990759e-07 -1.67680012e-09
+ 3.69090759e-07 2.45018676e-08 3.69190759e-07 7.39380085e-10 3.69290759e-07 2.22738644e-08 3.69390759e-07 2.74369891e-09 3.69490759e-07 2.04438306e-08 3.69590759e-07 4.39085479e-09 3.69690759e-07 1.89397881e-08 3.69790759e-07 5.74463174e-09
+ 3.69890759e-07 1.77036105e-08 3.69990759e-07 6.85732479e-09 3.70090759e-07 1.66875589e-08 3.70190759e-07 7.77189357e-09 3.70290759e-07 1.58524127e-08 3.70390759e-07 8.52363466e-09 3.70490759e-07 1.50671433e-08 3.70590759e-07 9.12775389e-09
+ 3.70690759e-07 1.45150393e-08 3.70790759e-07 9.62891189e-09 3.70890759e-07 1.40604611e-08 3.70990759e-07 1.00412063e-08 3.71090759e-07 1.36865216e-08 3.71190759e-07 1.03803583e-08 3.71290759e-07 1.33789217e-08 3.71390759e-07 1.06593409e-08
+ 3.71490759e-07 1.31258936e-08 3.71590759e-07 1.08888287e-08 3.71690759e-07 1.29177563e-08 3.71790759e-07 1.10776014e-08 3.71890759e-07 1.27465467e-08 3.71990759e-07 1.12328827e-08 3.72090759e-07 1.26057125e-08 3.72190759e-07 1.13606134e-08
+ 3.72290759e-07 1.24898661e-08 3.72390759e-07 1.14656818e-08 3.72490759e-07 1.23945733e-08 3.72590759e-07 1.15521083e-08 3.72690759e-07 1.23161877e-08 3.72790759e-07 1.1623201e-08 3.72890759e-07 1.22517099e-08 3.72990759e-07 1.16816798e-08
+ 3.73090759e-07 1.2198672e-08 3.73190759e-07 1.17297825e-08 3.73290759e-07 1.21550447e-08 3.73390759e-07 1.17693508e-08 3.73490759e-07 1.2119158e-08 3.73590759e-07 1.18018984e-08 3.73690759e-07 1.20896388e-08 3.73790759e-07 1.18286712e-08
+ 3.73890759e-07 1.20653571e-08 3.73990759e-07 1.18506933e-08 3.74090759e-07 1.20453839e-08 3.74190759e-07 1.18688085e-08 3.74290759e-07 1.20289544e-08 3.74390759e-07 1.18837093e-08 3.74490759e-07 1.20154398e-08 3.74590759e-07 1.18959663e-08
+ 3.74690759e-07 1.20043232e-08 3.74790759e-07 1.19060486e-08 3.74890759e-07 1.19951792e-08 3.74990759e-07 1.19143418e-08 3.75090759e-07 1.19876575e-08 3.75190759e-07 1.19211636e-08 3.75290759e-07 1.19814705e-08 3.75390759e-07 1.19267746e-08
+ 3.75490759e-07 1.19763813e-08 3.75590759e-07 1.19313906e-08 3.75690759e-07 1.19721951e-08 3.75790759e-07 1.19351871e-08 3.75890759e-07 1.1968752e-08 3.75990759e-07 1.19383102e-08 3.76090759e-07 1.19659191e-08 3.76190759e-07 1.19408792e-08
+ 3.76290759e-07 1.19635896e-08 3.76390759e-07 1.19429921e-08 3.76490759e-07 1.1961673e-08 3.76590759e-07 1.19447303e-08 3.76690759e-07 1.19600962e-08 3.76790759e-07 1.19461604e-08 3.76890759e-07 1.19587998e-08 3.76990759e-07 1.19473367e-08
+ 3.77090759e-07 1.19577328e-08 3.77190759e-07 1.19483037e-08 3.77290759e-07 1.19568556e-08 3.77390759e-07 1.19490997e-08 3.77490759e-07 1.19561338e-08 3.77590759e-07 1.1949754e-08 3.77690759e-07 1.19555401e-08 3.77790759e-07 1.19502923e-08
+ 3.77890759e-07 1.19550519e-08 3.77990759e-07 1.19507352e-08 3.78090759e-07 1.19546502e-08 3.78190759e-07 1.19510997e-08 3.78290759e-07 1.195432e-08 3.78390759e-07 1.19513993e-08 3.78490759e-07 1.19540481e-08 3.78590759e-07 1.19516457e-08
+ 3.78690759e-07 1.19538247e-08 3.78790759e-07 1.19518484e-08 3.78890759e-07 1.19536403e-08 3.78990759e-07 1.19520154e-08 3.79090759e-07 1.19534893e-08 3.79190759e-07 1.19521525e-08 3.79290759e-07 1.1953365e-08 3.79390759e-07 1.19522656e-08
+ 3.79490759e-07 1.19532626e-08 3.79590759e-07 1.19523582e-08 3.79690759e-07 1.19531783e-08 3.79790759e-07 1.19524344e-08 3.79890759e-07 1.19531096e-08 3.79990759e-07 1.19524973e-08 3.80090759e-07 1.19530524e-08 3.80190759e-07 1.19525491e-08
+ 3.80290759e-07 1.19530054e-08 3.80390759e-07 1.19525915e-08 3.80490759e-07 1.1952967e-08 3.80590759e-07 1.19526265e-08 3.80690759e-07 1.19529349e-08 3.80790759e-07 1.19526556e-08 3.80890759e-07 1.19529092e-08 3.80990759e-07 1.19526788e-08
+ 3.81090759e-07 1.19528875e-08 3.81190759e-07 1.19526982e-08 3.81290759e-07 1.19528699e-08 3.81390759e-07 1.19527144e-08 3.81490759e-07 1.19528554e-08 3.81590759e-07 1.19527274e-08 3.81690759e-07 1.19528434e-08 3.81790759e-07 1.19527383e-08
+ 3.81890759e-07 1.19528339e-08 3.81990759e-07 1.19527474e-08 3.82090759e-07 1.19528254e-08 3.82190759e-07 1.19527547e-08 3.82290759e-07 1.19528189e-08 3.82390759e-07 1.19527609e-08 3.82490759e-07 1.19528134e-08 3.82590759e-07 1.19527653e-08
+ 3.82690759e-07 1.19528089e-08 3.82790759e-07 1.19527697e-08 3.82890759e-07 1.19528051e-08 3.82990759e-07 1.19527729e-08 3.83090759e-07 1.19528021e-08 3.83190759e-07 1.19527757e-08 3.83290759e-07 1.19527996e-08 3.83390759e-07 1.19527782e-08
+ 3.83490759e-07 1.19527974e-08 3.83590759e-07 1.19527797e-08 3.83690759e-07 1.19527961e-08 3.83790759e-07 1.19527815e-08 3.83890759e-07 1.19527945e-08 3.83990759e-07 1.19527826e-08 3.84090759e-07 1.19527933e-08 3.84190759e-07 1.19527837e-08
+ 3.84290759e-07 1.19527925e-08 3.84390759e-07 1.19527844e-08 3.84490759e-07 1.1952792e-08 3.84590759e-07 1.1952785e-08 3.84690759e-07 1.19527912e-08 3.84790759e-07 1.19527855e-08 3.84890759e-07 1.19527909e-08 3.84990759e-07 1.19527858e-08
+ 3.85090759e-07 1.19527904e-08 3.85190759e-07 1.19527864e-08 3.85290759e-07 1.195279e-08 3.85390759e-07 1.19527868e-08 3.85490759e-07 1.19527897e-08 3.85590759e-07 1.1952787e-08 3.85690759e-07 1.19527895e-08 3.85790759e-07 1.19527871e-08
+ 3.85890759e-07 1.19527893e-08 3.85990759e-07 1.19527872e-08 3.86090759e-07 1.19527893e-08 3.86190759e-07 1.19527872e-08 3.86290759e-07 1.19527895e-08 3.86390759e-07 1.19527873e-08 3.86490759e-07 1.1952789e-08 3.86590759e-07 1.19527875e-08
+ 3.86690759e-07 1.1952789e-08 3.86790759e-07 1.19527878e-08 3.86890759e-07 1.19527889e-08 3.86990759e-07 1.19527879e-08 3.87090759e-07 1.19527889e-08 3.87190759e-07 1.19527879e-08 3.87290759e-07 1.19527887e-08 3.87390759e-07 1.1952788e-08
+ 3.87490759e-07 1.19527887e-08 3.87590759e-07 1.19527881e-08 3.87690759e-07 1.19527886e-08 3.87790759e-07 1.19527882e-08 3.87890759e-07 1.19527885e-08 3.87990759e-07 1.19527883e-08 3.88090759e-07 1.19527884e-08 3.88190759e-07 1.19527883e-08
+ 3.88290759e-07 1.19527885e-08 3.88390759e-07 1.19527883e-08 3.88490759e-07 1.19527885e-08 3.88590759e-07 1.19527883e-08 3.88690759e-07 1.19527885e-08 3.88790759e-07 1.19527883e-08 3.88890759e-07 1.19527885e-08 3.88990759e-07 1.19527883e-08
+ 3.89090759e-07 1.19527885e-08 3.89190759e-07 1.19527883e-08 3.89290759e-07 1.19527885e-08 3.89390759e-07 1.19527883e-08 3.89490759e-07 1.19527885e-08 3.89590759e-07 1.19527883e-08 3.89690759e-07 1.19527885e-08 3.89790759e-07 1.19527883e-08
+ 3.89890759e-07 1.19527885e-08 3.89990759e-07 1.19527883e-08 3.90090759e-07 1.19527885e-08 3.90190759e-07 1.19527883e-08 3.90290759e-07 1.19527885e-08 3.90390759e-07 1.19527883e-08 3.90490759e-07 1.19527885e-08 3.90590759e-07 1.19527883e-08
+ 3.90690759e-07 1.19527885e-08 3.90790759e-07 1.19527883e-08 3.90890759e-07 1.19527885e-08 3.90990759e-07 1.19527883e-08 3.91090759e-07 1.19527885e-08 3.91190759e-07 1.19527883e-08 3.91290759e-07 1.19527885e-08 3.91390759e-07 1.19527883e-08
+ 3.91490759e-07 1.19527885e-08 3.91590759e-07 1.19527883e-08 3.91690759e-07 1.19527885e-08 3.91790759e-07 1.19527883e-08 3.91890759e-07 1.19527885e-08 3.91990759e-07 1.19527883e-08 3.92090759e-07 1.19527885e-08 3.92190759e-07 1.19527883e-08
+ 3.92290759e-07 1.19527885e-08 3.92390759e-07 1.19527883e-08 3.92490759e-07 1.19527885e-08 3.92590759e-07 1.19527883e-08 3.92690759e-07 1.19527885e-08 3.92790759e-07 1.19527883e-08 3.92890759e-07 1.19527885e-08 3.92990759e-07 1.19527883e-08
+ 3.93090759e-07 1.19527885e-08 3.93190759e-07 1.19527883e-08 3.93290759e-07 1.19527885e-08 3.93390759e-07 1.19527883e-08 3.93490759e-07 1.19527885e-08 3.93590759e-07 1.19527883e-08 3.93690759e-07 1.19527885e-08 3.93790759e-07 1.19527883e-08
+ 3.93890759e-07 1.19527885e-08 3.93990759e-07 1.19527883e-08 3.94090759e-07 1.19527885e-08 3.94190759e-07 1.19527883e-08 3.94290759e-07 1.19527885e-08 3.94390759e-07 1.19527883e-08 3.94490759e-07 1.19527885e-08 3.94590759e-07 1.19527883e-08
+ 3.94690759e-07 1.19527885e-08 3.94790759e-07 1.19527883e-08 3.94890759e-07 1.19527885e-08 3.94990759e-07 1.19527883e-08 3.95090759e-07 1.19527885e-08 3.95190759e-07 1.19527883e-08 3.95290759e-07 1.19527885e-08 3.95390759e-07 1.19527883e-08
+ 3.95490759e-07 1.19527885e-08 3.95590759e-07 1.19527883e-08 3.95690759e-07 1.19527885e-08 3.95790759e-07 1.19527883e-08 3.95890759e-07 1.19527885e-08 3.95990759e-07 1.19527883e-08 3.96090759e-07 1.19527885e-08 3.96190759e-07 1.19527883e-08
+ 3.96290759e-07 1.19527885e-08 3.96390759e-07 1.19527883e-08 3.96490759e-07 1.19527885e-08 3.96590759e-07 1.19527883e-08 3.96690759e-07 1.19527885e-08 3.96790759e-07 1.19527883e-08 3.96890759e-07 1.19527885e-08 3.96990759e-07 1.19527883e-08
+ 3.97090759e-07 1.19527885e-08 3.97190759e-07 1.19527883e-08 3.97290759e-07 1.19527885e-08 3.97390759e-07 1.19527883e-08 3.97490759e-07 1.19527885e-08 3.97590759e-07 1.19527883e-08 3.97690759e-07 1.19527885e-08 3.97790759e-07 1.19527883e-08
+ 3.97890759e-07 1.19527885e-08 3.97990759e-07 1.19527883e-08 3.98090759e-07 1.19527885e-08 3.98190759e-07 1.19527883e-08 3.98290759e-07 1.19527885e-08 3.98390759e-07 1.19527883e-08 3.98490759e-07 1.19527885e-08 3.98590759e-07 1.19527883e-08
+ 3.98690759e-07 1.19527885e-08 3.98790759e-07 1.19527883e-08 3.98890759e-07 1.19527885e-08 3.98990759e-07 1.19527883e-08 3.99090759e-07 1.19527885e-08 3.99190759e-07 1.19527883e-08 3.99290759e-07 1.19527885e-08 3.99390759e-07 1.19527883e-08
+ 3.99490759e-07 1.19527885e-08 3.99590759e-07 1.19527883e-08 3.99690759e-07 1.19527885e-08 3.99790759e-07 1.19527883e-08 3.99890759e-07 1.19527885e-08 3.99990759e-07 1.19527883e-08 4e-07 1.19527885e-08 4.0001e-07 1.45272737e-08
+ 4.0003e-07 1.23606536e-09 4.0007e-07 2.76445116e-08 4.0015e-07 -4.38735384e-09 4.0025e-07 2.82154727e-08 4.0035e-07 -3.18927745e-09 4.0045e-07 2.52177678e-08 4.0055e-07 2.59407285e-09 4.0065e-07 -4.06359154e-08
+ 4.0075e-07 3.06902779e-06 4.0085e-07 9.4837652e-05 4.00931913e-07 -0.0447404595 4.01e-07 1.97335451 4.01008477e-07 3.09581876 4.01025432e-07 4.14108237 4.01059342e-07 4.88215046 4.01090545e-07 4.98042869
+ 4.01143412e-07 5.00336525 4.01199108e-07 4.99901157 4.01266691e-07 5.00044073 4.01329415e-07 4.99978464 4.01394829e-07 5.00011532 4.01464618e-07 4.99993177 4.01533535e-07 5.00004011 4.01610366e-07 4.99997429
+ 4.01709241e-07 5.00001814 4.01809241e-07 4.99998689 4.01909241e-07 5.00000939 4.02009241e-07 4.99999309 4.02109241e-07 5.000005 4.02209241e-07 4.99999625 4.02309241e-07 5.00000274 4.02409241e-07 4.99999789
+ 4.02509241e-07 5.00000154 4.02609241e-07 4.99999877 4.02709241e-07 5.00000089 4.02809241e-07 4.99999926 4.02909241e-07 5.00000052 4.03009241e-07 4.99999954 4.03109241e-07 5.00000031 4.03209241e-07 4.9999997
+ 4.03309241e-07 5.00000019 4.03409241e-07 4.9999998 4.03509241e-07 5.00000011 4.03609241e-07 4.99999986 4.03709241e-07 5.00000006 4.03809241e-07 4.9999999 4.03909241e-07 5.00000003 4.04009241e-07 4.99999992
+ 4.04109241e-07 5.00000001 4.04209241e-07 4.99999994 4.04309241e-07 5.0 4.04409241e-07 4.99999995 4.04509241e-07 4.99999999 4.04609241e-07 4.99999996 4.04709241e-07 4.99999999 4.04809241e-07 4.99999996
+ 4.04909241e-07 4.99999998 4.05009241e-07 4.99999996 4.05109241e-07 4.99999998 4.05209241e-07 4.99999997 4.05309241e-07 4.99999998 4.05409241e-07 4.99999997 4.05509241e-07 4.99999998 4.05609241e-07 4.99999997
+ 4.05709241e-07 4.99999997 4.05809241e-07 4.99999997 4.05909241e-07 4.99999997 4.06009241e-07 4.99999997 4.06109241e-07 4.99999997 4.06209241e-07 4.99999997 4.06309241e-07 4.99999997 4.06409241e-07 4.99999997
+ 4.06509241e-07 4.99999997 4.06609241e-07 4.99999997 4.06709241e-07 4.99999997 4.06809241e-07 4.99999997 4.06909241e-07 4.99999997 4.07009241e-07 4.99999997 4.07109241e-07 4.99999997 4.07209241e-07 4.99999997
+ 4.07309241e-07 4.99999997 4.07409241e-07 4.99999997 4.07509241e-07 4.99999997 4.07609241e-07 4.99999997 4.07709241e-07 4.99999997 4.07809241e-07 4.99999997 4.07909241e-07 4.99999997 4.08009241e-07 4.99999997
+ 4.08109241e-07 4.99999997 4.08209241e-07 4.99999997 4.08309241e-07 4.99999997 4.08409241e-07 4.99999997 4.08509241e-07 4.99999997 4.08609241e-07 4.99999997 4.08709241e-07 4.99999997 4.08809241e-07 4.99999997
+ 4.08909241e-07 4.99999997 4.09009241e-07 4.99999997 4.09109241e-07 4.99999997 4.09209241e-07 4.99999997 4.09309241e-07 4.99999997 4.09409241e-07 4.99999997 4.09509241e-07 4.99999997 4.09609241e-07 4.99999997
+ 4.09709241e-07 4.99999997 4.09809241e-07 4.99999997 4.09909241e-07 4.99999997 4.10009241e-07 4.99999997 4.10109241e-07 4.99999997 4.10209241e-07 4.99999997 4.10309241e-07 4.99999997 4.10409241e-07 4.99999997
+ 4.10509241e-07 4.99999997 4.10609241e-07 4.99999997 4.10709241e-07 4.99999997 4.10809241e-07 4.99999997 4.10909241e-07 4.99999997 4.11009241e-07 4.99999997 4.11109241e-07 4.99999997 4.11209241e-07 4.99999997
+ 4.11309241e-07 4.99999997 4.11409241e-07 4.99999997 4.11509241e-07 4.99999997 4.11609241e-07 4.99999997 4.11709241e-07 4.99999997 4.11809241e-07 4.99999997 4.11909241e-07 4.99999997 4.12009241e-07 4.99999997
+ 4.12109241e-07 4.99999997 4.12209241e-07 4.99999997 4.12309241e-07 4.99999997 4.12409241e-07 4.99999997 4.12509241e-07 4.99999997 4.12609241e-07 4.99999997 4.12709241e-07 4.99999997 4.12809241e-07 4.99999997
+ 4.12909241e-07 4.99999997 4.13009241e-07 4.99999997 4.13109241e-07 4.99999997 4.13209241e-07 4.99999997 4.13309241e-07 4.99999997 4.13409241e-07 4.99999997 4.13509241e-07 4.99999997 4.13609241e-07 4.99999997
+ 4.13709241e-07 4.99999997 4.13809241e-07 4.99999997 4.13909241e-07 4.99999997 4.14009241e-07 4.99999997 4.14109241e-07 4.99999997 4.14209241e-07 4.99999997 4.14309241e-07 4.99999997 4.14409241e-07 4.99999997
+ 4.14509241e-07 4.99999997 4.14609241e-07 4.99999997 4.14709241e-07 4.99999997 4.14809241e-07 4.99999997 4.14909241e-07 4.99999997 4.15009241e-07 4.99999997 4.15109241e-07 4.99999997 4.15209241e-07 4.99999997
+ 4.15309241e-07 4.99999997 4.15409241e-07 4.99999997 4.15509241e-07 4.99999997 4.15609241e-07 4.99999997 4.15709241e-07 4.99999997 4.15809241e-07 4.99999997 4.15909241e-07 4.99999997 4.16009241e-07 4.99999997
+ 4.16109241e-07 4.99999997 4.16209241e-07 4.99999997 4.16309241e-07 4.99999997 4.16409241e-07 4.99999997 4.16509241e-07 4.99999997 4.16609241e-07 4.99999997 4.16709241e-07 4.99999997 4.16809241e-07 4.99999997
+ 4.16909241e-07 4.99999997 4.17009241e-07 4.99999997 4.17109241e-07 4.99999997 4.17209241e-07 4.99999997 4.17309241e-07 4.99999997 4.17409241e-07 4.99999997 4.17509241e-07 4.99999997 4.17609241e-07 4.99999997
+ 4.17709241e-07 4.99999997 4.17809241e-07 4.99999997 4.17909241e-07 4.99999997 4.18009241e-07 4.99999997 4.18109241e-07 4.99999997 4.18209241e-07 4.99999997 4.18309241e-07 4.99999997 4.18409241e-07 4.99999997
+ 4.18509241e-07 4.99999997 4.18609241e-07 4.99999997 4.18709241e-07 4.99999997 4.18809241e-07 4.99999997 4.18909241e-07 4.99999997 4.19009241e-07 4.99999997 4.19109241e-07 4.99999997 4.19209241e-07 4.99999997
+ 4.19309241e-07 4.99999997 4.19409241e-07 4.99999997 4.19509241e-07 4.99999997 4.19609241e-07 4.99999997 4.19709241e-07 4.99999997 4.19809241e-07 4.99999997 4.19909241e-07 4.99999997 4.20009241e-07 4.99999997
+ 4.20109241e-07 4.99999997 4.20209241e-07 4.99999997 4.20309241e-07 4.99999997 4.20409241e-07 4.99999997 4.20509241e-07 4.99999997 4.20609241e-07 4.99999997 4.20709241e-07 4.99999997 4.20809241e-07 4.99999997
+ 4.20909241e-07 4.99999997 4.21009241e-07 4.99999997 4.21109241e-07 4.99999997 4.21209241e-07 4.99999997 4.21309241e-07 4.99999997 4.21409241e-07 4.99999997 4.21509241e-07 4.99999997 4.21609241e-07 4.99999997
+ 4.21709241e-07 4.99999997 4.21809241e-07 4.99999997 4.21909241e-07 4.99999997 4.22009241e-07 4.99999997 4.22109241e-07 4.99999997 4.22209241e-07 4.99999997 4.22309241e-07 4.99999997 4.22409241e-07 4.99999997
+ 4.22509241e-07 4.99999997 4.22609241e-07 4.99999997 4.22709241e-07 4.99999997 4.22809241e-07 4.99999997 4.22909241e-07 4.99999997 4.23009241e-07 4.99999997 4.23109241e-07 4.99999997 4.23209241e-07 4.99999997
+ 4.23309241e-07 4.99999997 4.23409241e-07 4.99999997 4.23509241e-07 4.99999997 4.23609241e-07 4.99999997 4.23709241e-07 4.99999997 4.23809241e-07 4.99999997 4.23909241e-07 4.99999997 4.24009241e-07 4.99999997
+ 4.24109241e-07 4.99999997 4.24209241e-07 4.99999997 4.24309241e-07 4.99999997 4.24409241e-07 4.99999997 4.24509241e-07 4.99999997 4.24609241e-07 4.99999997 4.24709241e-07 4.99999997 4.24809241e-07 4.99999997
+ 4.24909241e-07 4.99999997 4.25009241e-07 4.99999997 4.25109241e-07 4.99999997 4.25209241e-07 4.99999997 4.25309241e-07 4.99999997 4.25409241e-07 4.99999997 4.25509241e-07 4.99999997 4.25609241e-07 4.99999997
+ 4.25709241e-07 4.99999997 4.25809241e-07 4.99999997 4.25909241e-07 4.99999997 4.26009241e-07 4.99999997 4.26109241e-07 4.99999997 4.26209241e-07 4.99999997 4.26309241e-07 4.99999997 4.26409241e-07 4.99999997
+ 4.26509241e-07 4.99999997 4.26609241e-07 4.99999997 4.26709241e-07 4.99999997 4.26809241e-07 4.99999997 4.26909241e-07 4.99999997 4.27009241e-07 4.99999997 4.27109241e-07 4.99999997 4.27209241e-07 4.99999997
+ 4.27309241e-07 4.99999997 4.27409241e-07 4.99999997 4.27509241e-07 4.99999997 4.27609241e-07 4.99999997 4.27709241e-07 4.99999997 4.27809241e-07 4.99999997 4.27909241e-07 4.99999997 4.28009241e-07 4.99999997
+ 4.28109241e-07 4.99999997 4.28209241e-07 4.99999997 4.28309241e-07 4.99999997 4.28409241e-07 4.99999997 4.28509241e-07 4.99999997 4.28609241e-07 4.99999997 4.28709241e-07 4.99999997 4.28809241e-07 4.99999997
+ 4.28909241e-07 4.99999997 4.29009241e-07 4.99999997 4.29109241e-07 4.99999997 4.29209241e-07 4.99999997 4.29309241e-07 4.99999997 4.29409241e-07 4.99999997 4.29509241e-07 4.99999997 4.29609241e-07 4.99999997
+ 4.29709241e-07 4.99999997 4.29809241e-07 4.99999997 4.29909241e-07 4.99999997 4.30009241e-07 4.99999997 4.30109241e-07 4.99999997 4.30209241e-07 4.99999997 4.30309241e-07 4.99999997 4.30409241e-07 4.99999997
+ 4.30509241e-07 4.99999997 4.30609241e-07 4.99999997 4.30709241e-07 4.99999997 4.30809241e-07 4.99999997 4.30909241e-07 4.99999997 4.31009241e-07 4.99999997 4.31109241e-07 4.99999997 4.31209241e-07 4.99999997
+ 4.31309241e-07 4.99999997 4.31409241e-07 4.99999997 4.31509241e-07 4.99999997 4.31609241e-07 4.99999997 4.31709241e-07 4.99999997 4.31809241e-07 4.99999997 4.31909241e-07 4.99999997 4.32009241e-07 4.99999997
+ 4.32109241e-07 4.99999997 4.32209241e-07 4.99999997 4.32309241e-07 4.99999997 4.32409241e-07 4.99999997 4.32509241e-07 4.99999997 4.32609241e-07 4.99999997 4.32709241e-07 4.99999997 4.32809241e-07 4.99999997
+ 4.32909241e-07 4.99999997 4.33009241e-07 4.99999997 4.33109241e-07 4.99999997 4.33209241e-07 4.99999997 4.33309241e-07 4.99999997 4.33409241e-07 4.99999997 4.33509241e-07 4.99999997 4.33609241e-07 4.99999997
+ 4.33709241e-07 4.99999997 4.33809241e-07 4.99999997 4.33909241e-07 4.99999997 4.34009241e-07 4.99999997 4.34109241e-07 4.99999997 4.34209241e-07 4.99999997 4.34309241e-07 4.99999997 4.34409241e-07 4.99999997
+ 4.34509241e-07 4.99999997 4.34609241e-07 4.99999997 4.34709241e-07 4.99999997 4.34809241e-07 4.99999997 4.34909241e-07 4.99999997 4.35009241e-07 4.99999997 4.35109241e-07 4.99999997 4.35209241e-07 4.99999997
+ 4.35309241e-07 4.99999997 4.35409241e-07 4.99999997 4.35509241e-07 4.99999997 4.35609241e-07 4.99999997 4.35709241e-07 4.99999997 4.35809241e-07 4.99999997 4.35909241e-07 4.99999997 4.36009241e-07 4.99999997
+ 4.36109241e-07 4.99999997 4.36209241e-07 4.99999997 4.36309241e-07 4.99999997 4.36409241e-07 4.99999997 4.36509241e-07 4.99999997 4.36609241e-07 4.99999997 4.36709241e-07 4.99999997 4.36809241e-07 4.99999997
+ 4.36909241e-07 4.99999997 4.37009241e-07 4.99999997 4.37109241e-07 4.99999997 4.37209241e-07 4.99999997 4.37309241e-07 4.99999997 4.37409241e-07 4.99999997 4.37509241e-07 4.99999997 4.37609241e-07 4.99999997
+ 4.37709241e-07 4.99999997 4.37809241e-07 4.99999997 4.37909241e-07 4.99999997 4.38009241e-07 4.99999997 4.38109241e-07 4.99999997 4.38209241e-07 4.99999997 4.38309241e-07 4.99999997 4.38409241e-07 4.99999997
+ 4.38509241e-07 4.99999997 4.38609241e-07 4.99999997 4.38709241e-07 4.99999997 4.38809241e-07 4.99999997 4.38909241e-07 4.99999997 4.39009241e-07 4.99999997 4.39109241e-07 4.99999997 4.39209241e-07 4.99999997
+ 4.39309241e-07 4.99999997 4.39409241e-07 4.99999997 4.39509241e-07 4.99999997 4.39609241e-07 4.99999997 4.39709241e-07 4.99999997 4.39809241e-07 4.99999997 4.39909241e-07 4.99999997 4.40009241e-07 4.99999997
+ 4.40109241e-07 4.99999997 4.40209241e-07 4.99999997 4.40309241e-07 4.99999997 4.40409241e-07 4.99999997 4.40509241e-07 4.99999997 4.40609241e-07 4.99999997 4.40709241e-07 4.99999997 4.40809241e-07 4.99999997
+ 4.40909241e-07 4.99999997 4.41009241e-07 4.99999997 4.41109241e-07 4.99999997 4.41209241e-07 4.99999997 4.41309241e-07 4.99999997 4.41409241e-07 4.99999997 4.41509241e-07 4.99999997 4.41609241e-07 4.99999997
+ 4.41709241e-07 4.99999997 4.41809241e-07 4.99999997 4.41909241e-07 4.99999997 4.42009241e-07 4.99999997 4.42109241e-07 4.99999997 4.42209241e-07 4.99999997 4.42309241e-07 4.99999997 4.42409241e-07 4.99999997
+ 4.42509241e-07 4.99999997 4.42609241e-07 4.99999997 4.42709241e-07 4.99999997 4.42809241e-07 4.99999997 4.42909241e-07 4.99999997 4.43009241e-07 4.99999997 4.43109241e-07 4.99999997 4.43209241e-07 4.99999997
+ 4.43309241e-07 4.99999997 4.43409241e-07 4.99999997 4.43509241e-07 4.99999997 4.43609241e-07 4.99999997 4.43709241e-07 4.99999997 4.43809241e-07 4.99999997 4.43909241e-07 4.99999997 4.44009241e-07 4.99999997
+ 4.44109241e-07 4.99999997 4.44209241e-07 4.99999997 4.44309241e-07 4.99999997 4.44409241e-07 4.99999997 4.44509241e-07 4.99999997 4.44609241e-07 4.99999997 4.44709241e-07 4.99999997 4.44809241e-07 4.99999997
+ 4.44909241e-07 4.99999997 4.45009241e-07 4.99999997 4.45109241e-07 4.99999997 4.45209241e-07 4.99999997 4.45309241e-07 4.99999997 4.45409241e-07 4.99999997 4.45509241e-07 4.99999997 4.45609241e-07 4.99999997
+ 4.45709241e-07 4.99999997 4.45809241e-07 4.99999997 4.45909241e-07 4.99999997 4.46009241e-07 4.99999997 4.46109241e-07 4.99999997 4.46209241e-07 4.99999997 4.46309241e-07 4.99999997 4.46409241e-07 4.99999997
+ 4.46509241e-07 4.99999997 4.46609241e-07 4.99999997 4.46709241e-07 4.99999997 4.46809241e-07 4.99999997 4.46909241e-07 4.99999997 4.47009241e-07 4.99999997 4.47109241e-07 4.99999997 4.47209241e-07 4.99999997
+ 4.47309241e-07 4.99999997 4.47409241e-07 4.99999997 4.47509241e-07 4.99999997 4.47609241e-07 4.99999997 4.47709241e-07 4.99999997 4.47809241e-07 4.99999997 4.47909241e-07 4.99999997 4.48009241e-07 4.99999997
+ 4.48109241e-07 4.99999997 4.48209241e-07 4.99999997 4.48309241e-07 4.99999997 4.48409241e-07 4.99999997 4.48509241e-07 4.99999997 4.48609241e-07 4.99999997 4.48709241e-07 4.99999997 4.48809241e-07 4.99999997
+ 4.48909241e-07 4.99999997 4.49009241e-07 4.99999997 4.49109241e-07 4.99999997 4.49209241e-07 4.99999997 4.49309241e-07 4.99999997 4.49409241e-07 4.99999997 4.49509241e-07 4.99999997 4.49609241e-07 4.99999997
+ 4.49709241e-07 4.99999997 4.49809241e-07 4.99999997 4.49909241e-07 4.99999997 4.50009241e-07 4.99999997 4.50109241e-07 4.99999997 4.50209241e-07 4.99999997 4.50309241e-07 4.99999997 4.50409241e-07 4.99999997
+ 4.50509241e-07 4.99999997 4.50609241e-07 4.99999997 4.50709241e-07 4.99999997 4.50809241e-07 4.99999997 4.50909241e-07 4.99999997 4.51e-07 4.99999997 4.5101e-07 4.99999997 4.5103e-07 4.99999998
+ 4.5107e-07 4.99999996 4.5115e-07 4.99999998 4.5125e-07 4.99999997 4.5135e-07 4.99999997 4.5145e-07 4.99999998 4.5155e-07 4.99999996 4.5165e-07 4.99999998 4.5175e-07 4.99999996
+ 4.5185e-07 4.99999999 4.51930828e-07 5.00006476 4.52e-07 4.99916064 4.52008608e-07 4.99761639 4.52025825e-07 4.99311196 4.52060258e-07 5.01027311 4.52106181e-07 5.09906218 4.52150081e-07 4.21229454
+ 4.52198026e-07 0.290284903 4.5225538e-07 -0.0554592023 4.52312019e-07 0.0719468597 4.52404232e-07 -0.0579815953 4.52504232e-07 0.0528904133 4.52604232e-07 -0.0475729854 4.52704232e-07 0.0435757158 4.52804232e-07 -0.0393284178
+ 4.52904232e-07 0.0359989191 4.53004232e-07 -0.0325572549 4.53104232e-07 0.0297863163 4.53204232e-07 -0.0269831353 4.53304232e-07 0.024677895 4.53404232e-07 -0.0223854069 4.53504232e-07 0.0204676265 4.53604232e-07 -0.0185865295
+ 4.53704232e-07 0.0169908361 4.53804232e-07 -0.0154430663 4.53904232e-07 0.0141150741 4.54004232e-07 -0.0128386861 4.54104232e-07 0.0117332242 4.54204232e-07 -0.0106786681 4.54304232e-07 0.00975824024 4.54404232e-07 -0.00888561579
+ 4.54504232e-07 0.00811909449 4.54604232e-07 -0.00739609091 4.54704232e-07 0.00675762723 4.54804232e-07 -0.00615795518 4.54904232e-07 0.00562607399 4.55004232e-07 -0.00512825797 4.55104232e-07 0.00468510952 4.55204232e-07 -0.00427154749
+ 4.55304232e-07 0.00390228875 4.55404232e-07 -0.00355851286 4.55504232e-07 0.00325079606 4.55604232e-07 -0.00296488651 4.55704232e-07 0.002708436 4.55804232e-07 -0.0024705529 4.55904232e-07 0.00225681481 4.56004232e-07 -0.00205882186
+ 4.56104232e-07 0.00188067375 4.56204232e-07 -0.00171583399 4.56304232e-07 0.00156734401 4.56404232e-07 -0.00143007279 4.56504232e-07 0.00130629977 4.56604232e-07 -0.00119196316 4.56704232e-07 0.00108879052 4.56804232e-07 -0.000993540456
+ 4.56904232e-07 0.000907538165 4.57004232e-07 -0.000828177003 4.57104232e-07 0.000756486787 4.57204232e-07 -0.000690355922 4.57304232e-07 0.000630595752 4.57404232e-07 -0.00057548372 4.57504232e-07 0.00052566832 4.57604232e-07 -0.000479734899
+ 4.57704232e-07 0.000438209567 4.57804232e-07 -0.000399922963 4.57904232e-07 0.000365308462 4.58004232e-07 -0.000333393279 4.58104232e-07 0.000304539933 4.58204232e-07 -0.000277934025 4.58304232e-07 0.000253883483 4.58404232e-07 -0.000231702133
+ 4.58504232e-07 0.000211655506 4.58604232e-07 -0.000193161676 4.58704232e-07 0.00017645299 4.58804232e-07 -0.000161032592 4.58904232e-07 0.000147106668 4.59004232e-07 -0.000134248002 4.59104232e-07 0.000122642012 4.59204232e-07 -0.000111918653
+ 4.59304232e-07 0.000102246759 4.59404232e-07 -9.33033251e-05 4.59504232e-07 8.52438625e-05 4.59604232e-07 -7.7784159e-05 4.59704232e-07 7.10689667e-05 4.59804232e-07 -6.48461156e-05 4.59904232e-07 5.92516325e-05 4.60004232e-07 -5.40598536e-05
+ 4.60104232e-07 4.93997006e-05 4.60204232e-07 -4.50674637e-05 4.60304232e-07 4.11862589e-05 4.60404232e-07 -3.75705791e-05 4.60504232e-07 3.43387821e-05 4.60604232e-07 -3.13204668e-05 4.60704232e-07 2.86300807e-05 4.60804232e-07 -2.61097683e-05
+ 4.60904232e-07 2.38707567e-05 4.61004232e-07 -2.17656161e-05 4.61104232e-07 1.9902916e-05 4.61204232e-07 -1.81438953e-05 4.61304232e-07 1.65949268e-05 4.61404232e-07 -1.51244604e-05 4.61504232e-07 1.38370509e-05 4.61604232e-07 -1.26071484e-05
+ 4.61704232e-07 1.15378015e-05 4.61804232e-07 -1.05084548e-05 4.61904232e-07 9.62090748e-06 4.62004232e-07 -8.75876282e-06 4.62104232e-07 8.02278265e-06 4.62204232e-07 -7.30003353e-06 4.62304232e-07 6.69041563e-06 4.62404232e-07 -6.08388022e-06
+ 4.62504232e-07 5.57961123e-06 4.62604232e-07 -5.0699631e-06 4.62704232e-07 4.65352411e-06 4.62804232e-07 -4.22465098e-06 4.62904232e-07 3.88143644e-06 4.63004232e-07 -3.5199056e-06 4.63104232e-07 3.23773878e-06 4.63204232e-07 -2.93235145e-06
+ 4.63304232e-07 2.70108056e-06 4.63404232e-07 -2.44250033e-06 4.63504232e-07 2.2536618e-06 4.63604232e-07 -2.03410491e-06 4.63704232e-07 1.88064259e-06 4.63804232e-07 -1.69361974e-06 4.63904232e-07 1.56965094e-06 4.64004232e-07 -1.40079513e-06
+ 4.64104232e-07 1.32022171e-06 4.64204232e-07 -1.16495131e-06 4.64304232e-07 1.10221054e-06 4.64404232e-07 -9.68845144e-07 4.64504232e-07 9.20524804e-07 4.64604232e-07 -8.05378012e-07 4.64704232e-07 7.69073298e-07 4.64804232e-07 -6.69112945e-07
+ 4.64904232e-07 6.42824079e-07 4.65004232e-07 -5.55523017e-07 4.65104232e-07 5.37583116e-07 4.65204232e-07 -4.60834662e-07 4.65304232e-07 4.49854028e-07 4.65404232e-07 -3.81902011e-07 4.65504232e-07 3.76722691e-07 4.65604232e-07 -3.16103656e-07
+ 4.65704232e-07 3.15760337e-07 4.65804232e-07 -2.61254025e-07 4.65904232e-07 2.64941894e-07 4.66004232e-07 -2.15531318e-07 4.66104232e-07 2.22579736e-07 4.66204232e-07 -1.77426887e-07 4.66304232e-07 1.87286699e-07 4.66404232e-07 -1.45681874e-07
+ 4.66504232e-07 1.57883812e-07 4.66604232e-07 -1.19234754e-07 4.66704232e-07 1.33387825e-07 4.66804232e-07 -9.7201165e-08 4.66904232e-07 1.1297967e-07 4.67004232e-07 -7.88444124e-08 4.67104232e-07 9.59770696e-08 4.67204232e-07 -6.35509264e-08
+ 4.67304232e-07 8.18118435e-08 4.67404232e-07 -5.07711887e-08 4.67504232e-07 6.9971415e-08 4.67604232e-07 -4.0160915e-08 4.67704232e-07 6.01479454e-08 4.67804232e-07 -3.1325214e-08 4.67904232e-07 5.19642376e-08 4.68004232e-07 -2.39641145e-08
+ 4.68104232e-07 4.51463201e-08 4.68204232e-07 -1.78315383e-08 4.68304232e-07 3.94660681e-08 4.68404232e-07 -1.2721872e-08 4.68504232e-07 3.47333433e-08 4.68604232e-07 -8.46503093e-09 4.68704232e-07 3.07907578e-08 4.68804232e-07 -4.91886631e-09
+ 4.68904232e-07 2.75063602e-08 4.69004232e-07 -1.9646888e-09 4.69104232e-07 2.47702317e-08 4.69204232e-07 4.96362479e-10 4.69304232e-07 2.24973244e-08 4.69404232e-07 2.54107449e-09 4.69504232e-07 2.06302845e-08 4.69604232e-07 4.22167032e-09
+ 4.69704232e-07 1.90955796e-08 4.69804232e-07 5.6031679e-09 4.69904232e-07 1.78339728e-08 4.70004232e-07 6.73886061e-09 4.70104232e-07 1.67968122e-08 4.70204232e-07 7.67253117e-09 4.70304232e-07 1.59441263e-08 4.70404232e-07 8.44015202e-09
+ 4.70504232e-07 1.51437649e-08 4.70604232e-07 9.05741745e-09 4.70704232e-07 1.4579634e-08 4.70804232e-07 9.56956203e-09 4.70904232e-07 1.41150189e-08 4.71004232e-07 9.99102859e-09 4.71104232e-07 1.37326945e-08 4.71204232e-07 1.03378478e-08
+ 4.71304232e-07 1.34180805e-08 4.71404232e-07 1.062325e-08 4.71504232e-07 1.3159176e-08 4.71604232e-07 1.08581194e-08 4.71704232e-07 1.29461077e-08 4.71804232e-07 1.1051412e-08 4.71904232e-07 1.27707533e-08 4.72004232e-07 1.12104949e-08
+ 4.72104232e-07 1.262643e-08 4.72204232e-07 1.134143e-08 4.72304232e-07 1.25076398e-08 4.72404232e-07 1.14492033e-08 4.72504232e-07 1.24098596e-08 4.72604232e-07 1.15379188e-08 4.72704232e-07 1.23293677e-08 4.72804232e-07 1.1610951e-08
+ 4.72904232e-07 1.2263102e-08 4.73004232e-07 1.16710782e-08 4.73104232e-07 1.22085438e-08 4.73204232e-07 1.17205845e-08 4.73304232e-07 1.21636204e-08 4.73404232e-07 1.17613501e-08 4.73504232e-07 1.21266266e-08 4.73604232e-07 1.17949225e-08
+ 4.73704232e-07 1.2096159e-08 4.73804232e-07 1.18225736e-08 4.73904232e-07 1.20710629e-08 4.74004232e-07 1.18453513e-08 4.74104232e-07 1.20503886e-08 4.74204232e-07 1.1864117e-08 4.74304232e-07 1.20333541e-08 4.74404232e-07 1.18795807e-08
+ 4.74504232e-07 1.20193162e-08 4.74604232e-07 1.18923249e-08 4.74704232e-07 1.20077457e-08 4.74804232e-07 1.19028301e-08 4.74904232e-07 1.1998207e-08 4.75004232e-07 1.19114919e-08 4.75104232e-07 1.19903414e-08 4.75204232e-07 1.1918635e-08
+ 4.75304232e-07 1.19838537e-08 4.75404232e-07 1.19245278e-08 4.75504232e-07 1.19785012e-08 4.75604232e-07 1.192939e-08 4.75704232e-07 1.19740841e-08 4.75804232e-07 1.19334031e-08 4.75904232e-07 1.19704371e-08 4.76004232e-07 1.19367171e-08
+ 4.76104232e-07 1.19674258e-08 4.76204232e-07 1.19394543e-08 4.76304232e-07 1.19649374e-08 4.76404232e-07 1.19417164e-08 4.76504232e-07 1.19628805e-08 4.76604232e-07 1.19435865e-08 4.76704232e-07 1.196118e-08 4.76804232e-07 1.19451336e-08
+ 4.76904232e-07 1.19597726e-08 4.77004232e-07 1.19464138e-08 4.77104232e-07 1.19586077e-08 4.77204232e-07 1.19474739e-08 4.77304232e-07 1.19576427e-08 4.77404232e-07 1.19483529e-08 4.77504232e-07 1.19568424e-08 4.77604232e-07 1.19490813e-08
+ 4.77704232e-07 1.19561788e-08 4.77804232e-07 1.19496862e-08 4.77904232e-07 1.19556277e-08 4.78004232e-07 1.19501884e-08 4.78104232e-07 1.19551702e-08 4.78204232e-07 1.19506057e-08 4.78304232e-07 1.19547894e-08 4.78404232e-07 1.1950953e-08
+ 4.78504232e-07 1.19544725e-08 4.78604232e-07 1.19512423e-08 4.78704232e-07 1.19542082e-08 4.78804232e-07 1.19514837e-08 4.78904232e-07 1.19539876e-08 4.79004232e-07 1.19516851e-08 4.79104232e-07 1.19538035e-08 4.79204232e-07 1.19518536e-08
+ 4.79304232e-07 1.19536495e-08 4.79404232e-07 1.19519948e-08 4.79504232e-07 1.19535202e-08 4.79604232e-07 1.1952113e-08 4.79704232e-07 1.19534118e-08 4.79804232e-07 1.19522125e-08 4.79904232e-07 1.19533208e-08 4.80004232e-07 1.19522958e-08
+ 4.80104232e-07 1.19532439e-08 4.80204232e-07 1.19523663e-08 4.80304232e-07 1.19531791e-08 4.80404232e-07 1.19524258e-08 4.80504232e-07 1.19531248e-08 4.80604232e-07 1.19524758e-08 4.80704232e-07 1.19530783e-08 4.80804232e-07 1.19525187e-08
+ 4.80904232e-07 1.19530391e-08 4.81004232e-07 1.19525552e-08 4.81104232e-07 1.19530055e-08 4.81204232e-07 1.1952586e-08 4.81304232e-07 1.1952977e-08 4.81404232e-07 1.19526125e-08 4.81504232e-07 1.19529524e-08 4.81604232e-07 1.1952635e-08
+ 4.81704232e-07 1.19529315e-08 4.81804232e-07 1.19526543e-08 4.81904232e-07 1.19529137e-08 4.82004232e-07 1.19526708e-08 4.82104232e-07 1.19528984e-08 4.82204232e-07 1.19526852e-08 4.82304232e-07 1.1952885e-08 4.82404232e-07 1.19526976e-08
+ 4.82504232e-07 1.19528736e-08 4.82604232e-07 1.19527083e-08 4.82704232e-07 1.19528635e-08 4.82804232e-07 1.19527175e-08 4.82904232e-07 1.19528548e-08 4.83004232e-07 1.19527256e-08 4.83104232e-07 1.19528473e-08 4.83204232e-07 1.19527328e-08
+ 4.83304232e-07 1.19528407e-08 4.83404232e-07 1.19527389e-08 4.83504232e-07 1.19528349e-08 4.83604232e-07 1.19527445e-08 4.83704232e-07 1.19528298e-08 4.83804232e-07 1.19527492e-08 4.83904232e-07 1.19528253e-08 4.84004232e-07 1.19527536e-08
+ 4.84104232e-07 1.19528211e-08 4.84204232e-07 1.19527571e-08 4.84304232e-07 1.19528178e-08 4.84404232e-07 1.19527602e-08 4.84504232e-07 1.19528147e-08 4.84604232e-07 1.19527633e-08 4.84704232e-07 1.19528119e-08 4.84804232e-07 1.19527657e-08
+ 4.84904232e-07 1.19528096e-08 4.85004232e-07 1.19527682e-08 4.85104232e-07 1.19528074e-08 4.85204232e-07 1.195277e-08 4.85304232e-07 1.19528055e-08 4.85404232e-07 1.19527721e-08 4.85504232e-07 1.19528036e-08 4.85604232e-07 1.19527737e-08
+ 4.85704232e-07 1.19528021e-08 4.85804232e-07 1.19527753e-08 4.85904232e-07 1.19528009e-08 4.86004232e-07 1.19527765e-08 4.86104232e-07 1.19527997e-08 4.86204232e-07 1.19527773e-08 4.86304232e-07 1.19527987e-08 4.86404232e-07 1.19527784e-08
+ 4.86504232e-07 1.19527976e-08 4.86604232e-07 1.19527795e-08 4.86704232e-07 1.19527965e-08 4.86804232e-07 1.19527806e-08 4.86904232e-07 1.19527958e-08 4.87004232e-07 1.19527815e-08 4.87104232e-07 1.19527949e-08 4.87204232e-07 1.1952782e-08
+ 4.87304232e-07 1.19527943e-08 4.87404232e-07 1.19527827e-08 4.87504232e-07 1.19527936e-08 4.87604232e-07 1.1952783e-08 4.87704232e-07 1.19527934e-08 4.87804232e-07 1.19527834e-08 4.87904232e-07 1.19527929e-08 4.88004232e-07 1.19527841e-08
+ 4.88104232e-07 1.19527923e-08 4.88204232e-07 1.19527846e-08 4.88304232e-07 1.19527918e-08 4.88404232e-07 1.19527848e-08 4.88504232e-07 1.19527917e-08 4.88604232e-07 1.19527852e-08 4.88704232e-07 1.19527915e-08 4.88804232e-07 1.19527855e-08
+ 4.88904232e-07 1.19527911e-08 4.89004232e-07 1.19527857e-08 4.89104232e-07 1.19527907e-08 4.89204232e-07 1.19527859e-08 4.89304232e-07 1.19527907e-08 4.89404232e-07 1.19527863e-08 4.89504232e-07 1.19527904e-08 4.89604232e-07 1.19527866e-08
+ 4.89704232e-07 1.19527898e-08 4.89804232e-07 1.19527868e-08 4.89904232e-07 1.19527897e-08 4.90004232e-07 1.19527869e-08 4.90104232e-07 1.19527897e-08 4.90204232e-07 1.19527868e-08 4.90304232e-07 1.19527899e-08 4.90404232e-07 1.1952787e-08
+ 4.90504232e-07 1.19527897e-08 4.90604232e-07 1.1952787e-08 4.90704232e-07 1.19527898e-08 4.90804232e-07 1.1952787e-08 4.90904232e-07 1.19527898e-08 4.91004232e-07 1.1952787e-08 4.91104232e-07 1.19527894e-08 4.91204232e-07 1.19527871e-08
+ 4.91304232e-07 1.19527895e-08 4.91404232e-07 1.19527871e-08 4.91504232e-07 1.19527893e-08 4.91604232e-07 1.19527872e-08 4.91704232e-07 1.19527897e-08 4.91804232e-07 1.19527872e-08 4.91904232e-07 1.19527895e-08 4.92004232e-07 1.19527873e-08
+ 4.92104232e-07 1.19527893e-08 4.92204232e-07 1.19527873e-08 4.92304232e-07 1.19527895e-08 4.92404232e-07 1.19527873e-08 4.92504232e-07 1.19527894e-08 4.92604232e-07 1.19527874e-08 4.92704232e-07 1.19527892e-08 4.92804232e-07 1.19527876e-08
+ 4.92904232e-07 1.19527893e-08 4.93004232e-07 1.19527876e-08 4.93104232e-07 1.1952789e-08 4.93204232e-07 1.19527878e-08 4.93304232e-07 1.19527891e-08 4.93404232e-07 1.19527878e-08 4.93504232e-07 1.1952789e-08 4.93604232e-07 1.19527878e-08
+ 4.93704232e-07 1.1952789e-08 4.93804232e-07 1.19527878e-08 4.93904232e-07 1.19527889e-08 4.94004232e-07 1.19527879e-08 4.94104232e-07 1.1952789e-08 4.94204232e-07 1.19527879e-08 4.94304232e-07 1.19527889e-08 4.94404232e-07 1.19527879e-08
+ 4.94504232e-07 1.1952789e-08 4.94604232e-07 1.19527879e-08 4.94704232e-07 1.19527888e-08 4.94804232e-07 1.1952788e-08 4.94904232e-07 1.19527887e-08 4.95004232e-07 1.19527881e-08 4.95104232e-07 1.19527886e-08 4.95204232e-07 1.19527882e-08
+ 4.95304232e-07 1.19527885e-08 4.95404232e-07 1.19527882e-08 4.95504232e-07 1.19527886e-08 4.95604232e-07 1.19527883e-08 4.95704232e-07 1.19527884e-08 4.95804232e-07 1.19527883e-08 4.95904232e-07 1.19527885e-08 4.96004232e-07 1.19527883e-08
+ 4.96104232e-07 1.19527884e-08 4.96204232e-07 1.19527883e-08 4.96304232e-07 1.19527885e-08 4.96404232e-07 1.19527883e-08 4.96504232e-07 1.19527884e-08 4.96604232e-07 1.19527883e-08 4.96704232e-07 1.19527884e-08 4.96804232e-07 1.19527883e-08
+ 4.96904232e-07 1.19527884e-08 4.97004232e-07 1.19527883e-08 4.97104232e-07 1.19527885e-08 4.97204232e-07 1.19527883e-08 4.97304232e-07 1.19527884e-08 4.97404232e-07 1.19527883e-08 4.97504232e-07 1.19527884e-08 4.97604232e-07 1.19527883e-08
+ 4.97704232e-07 1.19527884e-08 4.97804232e-07 1.19527883e-08 4.97904232e-07 1.19527884e-08 4.98004232e-07 1.19527883e-08 4.98104232e-07 1.19527884e-08 4.98204232e-07 1.19527883e-08 4.98304232e-07 1.19527884e-08 4.98404232e-07 1.19527883e-08
+ 4.98504232e-07 1.19527884e-08 4.98604232e-07 1.19527883e-08 4.98704232e-07 1.19527884e-08 4.98804232e-07 1.19527883e-08 4.98904232e-07 1.19527885e-08 4.99004232e-07 1.19527883e-08 4.99104232e-07 1.19527884e-08 4.99204232e-07 1.19527883e-08
+ 4.99304232e-07 1.19527884e-08 4.99404232e-07 1.19527883e-08 4.99504232e-07 1.19527884e-08 4.99604232e-07 1.19527883e-08 4.99704232e-07 1.19527884e-08 4.99804232e-07 1.19527883e-08 4.99904232e-07 1.19527884e-08 5e-07 1.19527884e-08
+ 5.0001e-07 1.45267509e-08 5.0003e-07 1.23970223e-09 5.0007e-07 2.7637525e-08 5.0015e-07 -4.37848716e-09 5.0025e-07 2.82049084e-08 5.0035e-07 -3.17727716e-09 5.0045e-07 2.52046159e-08 5.0055e-07 2.60784397e-09
+ 5.0065e-07 -4.06484961e-08 5.0075e-07 3.06912285e-06 5.0085e-07 9.51416721e-05 5.00932051e-07 -0.0447831027 5.01e-07 1.97583273 5.01008488e-07 3.09989962 5.01025463e-07 4.14313244 5.01059414e-07 4.88304728
+ 5.0109062e-07 4.97992695 5.0114347e-07 5.00280645 5.01199151e-07 4.99919782 5.01299151e-07 5.00046536 5.01399151e-07 4.99971259 5.01499151e-07 5.00018323 5.01599151e-07 4.99987811 5.01699151e-07 5.00008217
+ 5.01799151e-07 4.99994319 5.01893327e-07 5.00003835 5.01993327e-07 4.99997304 5.02093327e-07 5.00001879 5.02193327e-07 4.99998671 5.02293327e-07 5.00000926 5.02393327e-07 4.99999342 5.02493327e-07 5.00000455
+ 5.02593327e-07 4.99999675 5.02693327e-07 5.00000222 5.02793327e-07 4.9999984 5.02893327e-07 5.00000107 5.02993327e-07 4.99999921 5.03093327e-07 5.0000005 5.03193327e-07 4.99999961 5.03293327e-07 5.00000022
+ 5.03393327e-07 4.9999998 5.03493327e-07 5.00000008 5.03593327e-07 4.9999999 5.03693327e-07 5.00000002 5.03793327e-07 4.99999994 5.03893327e-07 4.99999999 5.03993327e-07 4.99999996 5.04093327e-07 4.99999998
+ 5.04193327e-07 4.99999997 5.04293327e-07 4.99999997 5.04393327e-07 4.99999997 5.04493327e-07 4.99999997 5.04593327e-07 4.99999997 5.04693327e-07 4.99999997 5.04793327e-07 4.99999997 5.04893327e-07 4.99999997
+ 5.04993327e-07 4.99999997 5.05093327e-07 4.99999997 5.05193327e-07 4.99999997 5.05293327e-07 4.99999997 5.05393327e-07 4.99999997 5.05493327e-07 4.99999997 5.05593327e-07 4.99999997 5.05693327e-07 4.99999997
+ 5.05793327e-07 4.99999997 5.05893327e-07 4.99999997 5.05993327e-07 4.99999997 5.06093327e-07 4.99999997 5.06193327e-07 4.99999997 5.06293327e-07 4.99999997 5.06393327e-07 4.99999997 5.06493327e-07 4.99999997
+ 5.06593327e-07 4.99999997 5.06693327e-07 4.99999997 5.06793327e-07 4.99999997 5.06893327e-07 4.99999997 5.06993327e-07 4.99999997 5.07093327e-07 4.99999997 5.07193327e-07 4.99999997 5.07293327e-07 4.99999997
+ 5.07393327e-07 4.99999997 5.07493327e-07 4.99999997 5.07593327e-07 4.99999997 5.07693327e-07 4.99999997 5.07793327e-07 4.99999997 5.07893327e-07 4.99999997 5.07993327e-07 4.99999997 5.08093327e-07 4.99999997
+ 5.08193327e-07 4.99999997 5.08293327e-07 4.99999997 5.08393327e-07 4.99999997 5.08493327e-07 4.99999997 5.08593327e-07 4.99999997 5.08693327e-07 4.99999997 5.08793327e-07 4.99999997 5.08893327e-07 4.99999997
+ 5.08993327e-07 4.99999997 5.09093327e-07 4.99999997 5.09193327e-07 4.99999997 5.09293327e-07 4.99999997 5.09393327e-07 4.99999997 5.09493327e-07 4.99999997 5.09593327e-07 4.99999997 5.09693327e-07 4.99999997
+ 5.09793327e-07 4.99999997 5.09893327e-07 4.99999997 5.09993327e-07 4.99999997 5.10093327e-07 4.99999997 5.10193327e-07 4.99999997 5.10293327e-07 4.99999997 5.10393327e-07 4.99999997 5.10493327e-07 4.99999997
+ 5.10593327e-07 4.99999997 5.10693327e-07 4.99999997 5.10793327e-07 4.99999997 5.10893327e-07 4.99999997 5.10993327e-07 4.99999997 5.11093327e-07 4.99999997 5.11193327e-07 4.99999997 5.11293327e-07 4.99999997
+ 5.11393327e-07 4.99999997 5.11493327e-07 4.99999997 5.11593327e-07 4.99999997 5.11693327e-07 4.99999997 5.11793327e-07 4.99999997 5.11893327e-07 4.99999997 5.11993327e-07 4.99999997 5.12093327e-07 4.99999997
+ 5.12193327e-07 4.99999997 5.12293327e-07 4.99999997 5.12393327e-07 4.99999997 5.12493327e-07 4.99999997 5.12593327e-07 4.99999997 5.12693327e-07 4.99999997 5.12793327e-07 4.99999997 5.12893327e-07 4.99999997
+ 5.12993327e-07 4.99999997 5.13093327e-07 4.99999997 5.13193327e-07 4.99999997 5.13293327e-07 4.99999997 5.13393327e-07 4.99999997 5.13493327e-07 4.99999997 5.13593327e-07 4.99999997 5.13693327e-07 4.99999997
+ 5.13793327e-07 4.99999997 5.13893327e-07 4.99999997 5.13993327e-07 4.99999997 5.14093327e-07 4.99999997 5.14193327e-07 4.99999997 5.14293327e-07 4.99999997 5.14393327e-07 4.99999997 5.14493327e-07 4.99999997
+ 5.14593327e-07 4.99999997 5.14693327e-07 4.99999997 5.14793327e-07 4.99999997 5.14893327e-07 4.99999997 5.14993327e-07 4.99999997 5.15093327e-07 4.99999997 5.15193327e-07 4.99999997 5.15293327e-07 4.99999997
+ 5.15393327e-07 4.99999997 5.15493327e-07 4.99999997 5.15593327e-07 4.99999997 5.15693327e-07 4.99999997 5.15793327e-07 4.99999997 5.15893327e-07 4.99999997 5.15993327e-07 4.99999997 5.16093327e-07 4.99999997
+ 5.16193327e-07 4.99999997 5.16293327e-07 4.99999997 5.16393327e-07 4.99999997 5.16493327e-07 4.99999997 5.16593327e-07 4.99999997 5.16693327e-07 4.99999997 5.16793327e-07 4.99999997 5.16893327e-07 4.99999997
+ 5.16993327e-07 4.99999997 5.17093327e-07 4.99999997 5.17193327e-07 4.99999997 5.17293327e-07 4.99999997 5.17393327e-07 4.99999997 5.17493327e-07 4.99999997 5.17593327e-07 4.99999997 5.17693327e-07 4.99999997
+ 5.17793327e-07 4.99999997 5.17893327e-07 4.99999997 5.17993327e-07 4.99999997 5.18093327e-07 4.99999997 5.18193327e-07 4.99999997 5.18293327e-07 4.99999997 5.18393327e-07 4.99999997 5.18493327e-07 4.99999997
+ 5.18593327e-07 4.99999997 5.18693327e-07 4.99999997 5.18793327e-07 4.99999997 5.18893327e-07 4.99999997 5.18993327e-07 4.99999997 5.19093327e-07 4.99999997 5.19193327e-07 4.99999997 5.19293327e-07 4.99999997
+ 5.19393327e-07 4.99999997 5.19493327e-07 4.99999997 5.19593327e-07 4.99999997 5.19693327e-07 4.99999997 5.19793327e-07 4.99999997 5.19893327e-07 4.99999997 5.19993327e-07 4.99999997 5.20093327e-07 4.99999997
+ 5.20193327e-07 4.99999997 5.20293327e-07 4.99999997 5.20393327e-07 4.99999997 5.20493327e-07 4.99999997 5.20593327e-07 4.99999997 5.20693327e-07 4.99999997 5.20793327e-07 4.99999997 5.20893327e-07 4.99999997
+ 5.20993327e-07 4.99999997 5.21093327e-07 4.99999997 5.21193327e-07 4.99999997 5.21293327e-07 4.99999997 5.21393327e-07 4.99999997 5.21493327e-07 4.99999997 5.21593327e-07 4.99999997 5.21693327e-07 4.99999997
+ 5.21793327e-07 4.99999997 5.21893327e-07 4.99999997 5.21993327e-07 4.99999997 5.22093327e-07 4.99999997 5.22193327e-07 4.99999997 5.22293327e-07 4.99999997 5.22393327e-07 4.99999997 5.22493327e-07 4.99999997
+ 5.22593327e-07 4.99999997 5.22693327e-07 4.99999997 5.22793327e-07 4.99999997 5.22893327e-07 4.99999997 5.22993327e-07 4.99999997 5.23093327e-07 4.99999997 5.23193327e-07 4.99999997 5.23293327e-07 4.99999997
+ 5.23393327e-07 4.99999997 5.23493327e-07 4.99999997 5.23593327e-07 4.99999997 5.23693327e-07 4.99999997 5.23793327e-07 4.99999997 5.23893327e-07 4.99999997 5.23993327e-07 4.99999997 5.24093327e-07 4.99999997
+ 5.24193327e-07 4.99999997 5.24293327e-07 4.99999997 5.24393327e-07 4.99999997 5.24493327e-07 4.99999997 5.24593327e-07 4.99999997 5.24693327e-07 4.99999997 5.24793327e-07 4.99999997 5.24893327e-07 4.99999997
+ 5.24993327e-07 4.99999997 5.25093327e-07 4.99999997 5.25193327e-07 4.99999997 5.25293327e-07 4.99999997 5.25393327e-07 4.99999997 5.25493327e-07 4.99999997 5.25593327e-07 4.99999997 5.25693327e-07 4.99999997
+ 5.25793327e-07 4.99999997 5.25893327e-07 4.99999997 5.25993327e-07 4.99999997 5.26093327e-07 4.99999997 5.26193327e-07 4.99999997 5.26293327e-07 4.99999997 5.26393327e-07 4.99999997 5.26493327e-07 4.99999997
+ 5.26593327e-07 4.99999997 5.26693327e-07 4.99999997 5.26793327e-07 4.99999997 5.26893327e-07 4.99999997 5.26993327e-07 4.99999997 5.27093327e-07 4.99999997 5.27193327e-07 4.99999997 5.27293327e-07 4.99999997
+ 5.27393327e-07 4.99999997 5.27493327e-07 4.99999997 5.27593327e-07 4.99999997 5.27693327e-07 4.99999997 5.27793327e-07 4.99999997 5.27893327e-07 4.99999997 5.27993327e-07 4.99999997 5.28093327e-07 4.99999997
+ 5.28193327e-07 4.99999997 5.28293327e-07 4.99999997 5.28393327e-07 4.99999997 5.28493327e-07 4.99999997 5.28593327e-07 4.99999997 5.28693327e-07 4.99999997 5.28793327e-07 4.99999997 5.28893327e-07 4.99999997
+ 5.28993327e-07 4.99999997 5.29093327e-07 4.99999997 5.29193327e-07 4.99999997 5.29293327e-07 4.99999997 5.29393327e-07 4.99999997 5.29493327e-07 4.99999997 5.29593327e-07 4.99999997 5.29693327e-07 4.99999997
+ 5.29793327e-07 4.99999997 5.29893327e-07 4.99999997 5.29993327e-07 4.99999997 5.30093327e-07 4.99999997 5.30193327e-07 4.99999997 5.30293327e-07 4.99999997 5.30393327e-07 4.99999997 5.30493327e-07 4.99999997
+ 5.30593327e-07 4.99999997 5.30693327e-07 4.99999997 5.30793327e-07 4.99999997 5.30893327e-07 4.99999997 5.30993327e-07 4.99999997 5.31093327e-07 4.99999997 5.31193327e-07 4.99999997 5.31293327e-07 4.99999997
+ 5.31393327e-07 4.99999997 5.31493327e-07 4.99999997 5.31593327e-07 4.99999997 5.31693327e-07 4.99999997 5.31793327e-07 4.99999997 5.31893327e-07 4.99999997 5.31993327e-07 4.99999997 5.32093327e-07 4.99999997
+ 5.32193327e-07 4.99999997 5.32293327e-07 4.99999997 5.32393327e-07 4.99999997 5.32493327e-07 4.99999997 5.32593327e-07 4.99999997 5.32693327e-07 4.99999997 5.32793327e-07 4.99999997 5.32893327e-07 4.99999997
+ 5.32993327e-07 4.99999997 5.33093327e-07 4.99999997 5.33193327e-07 4.99999997 5.33293327e-07 4.99999997 5.33393327e-07 4.99999997 5.33493327e-07 4.99999997 5.33593327e-07 4.99999997 5.33693327e-07 4.99999997
+ 5.33793327e-07 4.99999997 5.33893327e-07 4.99999997 5.33993327e-07 4.99999997 5.34093327e-07 4.99999997 5.34193327e-07 4.99999997 5.34293327e-07 4.99999997 5.34393327e-07 4.99999997 5.34493327e-07 4.99999997
+ 5.34593327e-07 4.99999997 5.34693327e-07 4.99999997 5.34793327e-07 4.99999997 5.34893327e-07 4.99999997 5.34993327e-07 4.99999997 5.35093327e-07 4.99999997 5.35193327e-07 4.99999997 5.35293327e-07 4.99999997
+ 5.35393327e-07 4.99999997 5.35493327e-07 4.99999997 5.35593327e-07 4.99999997 5.35693327e-07 4.99999997 5.35793327e-07 4.99999997 5.35893327e-07 4.99999997 5.35993327e-07 4.99999997 5.36093327e-07 4.99999997
+ 5.36193327e-07 4.99999997 5.36293327e-07 4.99999997 5.36393327e-07 4.99999997 5.36493327e-07 4.99999997 5.36593327e-07 4.99999997 5.36693327e-07 4.99999997 5.36793327e-07 4.99999997 5.36893327e-07 4.99999997
+ 5.36993327e-07 4.99999997 5.37093327e-07 4.99999997 5.37193327e-07 4.99999997 5.37293327e-07 4.99999997 5.37393327e-07 4.99999997 5.37493327e-07 4.99999997 5.37593327e-07 4.99999997 5.37693327e-07 4.99999997
+ 5.37793327e-07 4.99999997 5.37893327e-07 4.99999997 5.37993327e-07 4.99999997 5.38093327e-07 4.99999997 5.38193327e-07 4.99999997 5.38293327e-07 4.99999997 5.38393327e-07 4.99999997 5.38493327e-07 4.99999997
+ 5.38593327e-07 4.99999997 5.38693327e-07 4.99999997 5.38793327e-07 4.99999997 5.38893327e-07 4.99999997 5.38993327e-07 4.99999997 5.39093327e-07 4.99999997 5.39193327e-07 4.99999997 5.39293327e-07 4.99999997
+ 5.39393327e-07 4.99999997 5.39493327e-07 4.99999997 5.39593327e-07 4.99999997 5.39693327e-07 4.99999997 5.39793327e-07 4.99999997 5.39893327e-07 4.99999997 5.39993327e-07 4.99999997 5.40093327e-07 4.99999997
+ 5.40193327e-07 4.99999997 5.40293327e-07 4.99999997 5.40393327e-07 4.99999997 5.40493327e-07 4.99999997 5.40593327e-07 4.99999997 5.40693327e-07 4.99999997 5.40793327e-07 4.99999997 5.40893327e-07 4.99999997
+ 5.40993327e-07 4.99999997 5.41093327e-07 4.99999997 5.41193327e-07 4.99999997 5.41293327e-07 4.99999997 5.41393327e-07 4.99999997 5.41493327e-07 4.99999997 5.41593327e-07 4.99999997 5.41693327e-07 4.99999997
+ 5.41793327e-07 4.99999997 5.41893327e-07 4.99999997 5.41993327e-07 4.99999997 5.42093327e-07 4.99999997 5.42193327e-07 4.99999997 5.42293327e-07 4.99999997 5.42393327e-07 4.99999997 5.42493327e-07 4.99999997
+ 5.42593327e-07 4.99999997 5.42693327e-07 4.99999997 5.42793327e-07 4.99999997 5.42893327e-07 4.99999997 5.42993327e-07 4.99999997 5.43093327e-07 4.99999997 5.43193327e-07 4.99999997 5.43293327e-07 4.99999997
+ 5.43393327e-07 4.99999997 5.43493327e-07 4.99999997 5.43593327e-07 4.99999997 5.43693327e-07 4.99999997 5.43793327e-07 4.99999997 5.43893327e-07 4.99999997 5.43993327e-07 4.99999997 5.44093327e-07 4.99999997
+ 5.44193327e-07 4.99999997 5.44293327e-07 4.99999997 5.44393327e-07 4.99999997 5.44493327e-07 4.99999997 5.44593327e-07 4.99999997 5.44693327e-07 4.99999997 5.44793327e-07 4.99999997 5.44893327e-07 4.99999997
+ 5.44993327e-07 4.99999997 5.45093327e-07 4.99999997 5.45193327e-07 4.99999997 5.45293327e-07 4.99999997 5.45393327e-07 4.99999997 5.45493327e-07 4.99999997 5.45593327e-07 4.99999997 5.45693327e-07 4.99999997
+ 5.45793327e-07 4.99999997 5.45893327e-07 4.99999997 5.45993327e-07 4.99999997 5.46093327e-07 4.99999997 5.46193327e-07 4.99999997 5.46293327e-07 4.99999997 5.46393327e-07 4.99999997 5.46493327e-07 4.99999997
+ 5.46593327e-07 4.99999997 5.46693327e-07 4.99999997 5.46793327e-07 4.99999997 5.46893327e-07 4.99999997 5.46993327e-07 4.99999997 5.47093327e-07 4.99999997 5.47193327e-07 4.99999997 5.47293327e-07 4.99999997
+ 5.47393327e-07 4.99999997 5.47493327e-07 4.99999997 5.47593327e-07 4.99999997 5.47693327e-07 4.99999997 5.47793327e-07 4.99999997 5.47893327e-07 4.99999997 5.47993327e-07 4.99999997 5.48093327e-07 4.99999997
+ 5.48193327e-07 4.99999997 5.48293327e-07 4.99999997 5.48393327e-07 4.99999997 5.48493327e-07 4.99999997 5.48593327e-07 4.99999997 5.48693327e-07 4.99999997 5.48793327e-07 4.99999997 5.48893327e-07 4.99999997
+ 5.48993327e-07 4.99999997 5.49093327e-07 4.99999997 5.49193327e-07 4.99999997 5.49293327e-07 4.99999997 5.49393327e-07 4.99999997 5.49493327e-07 4.99999997 5.49593327e-07 4.99999997 5.49693327e-07 4.99999997
+ 5.49793327e-07 4.99999997 5.49893327e-07 4.99999997 5.49993327e-07 4.99999997 5.50093327e-07 4.99999997 5.50193327e-07 4.99999997 5.50293327e-07 4.99999997 5.50393327e-07 4.99999997 5.50493327e-07 4.99999997
+ 5.50593327e-07 4.99999997 5.50693327e-07 4.99999997 5.50793327e-07 4.99999997 5.50893327e-07 4.99999997 5.50993327e-07 4.99999997 5.51e-07 4.99999997 5.5101e-07 4.99999997 5.5103e-07 4.99999998
+ 5.5107e-07 4.99999996 5.5115e-07 4.99999998 5.5125e-07 4.99999997 5.5135e-07 4.99999997 5.5145e-07 4.99999998 5.5155e-07 4.99999996 5.5165e-07 4.99999998 5.5175e-07 4.99999996
+ 5.5185e-07 4.99999999 5.51930828e-07 5.00006471 5.52e-07 4.99916174 5.52008608e-07 4.99761843 5.52025825e-07 4.99312395 5.52060258e-07 5.01021614 5.52106188e-07 5.09915398 5.52150118e-07 4.21384241
+ 5.5219811e-07 0.290133164 5.52255501e-07 -0.0555601235 5.52312176e-07 0.071992207 5.52404431e-07 -0.0580455459 5.52490774e-07 0.0521266462 5.52590774e-07 -0.046900588 5.52690774e-07 0.042974581 5.52790774e-07 -0.0387934186
+ 5.52890774e-07 0.0355083829 5.52990774e-07 -0.0321185209 5.53090774e-07 0.0293845439 5.53190774e-07 -0.0266224795 5.53290774e-07 0.0243478875 5.53390774e-07 -0.0220883003 5.53490774e-07 0.0201959102 5.53590774e-07 -0.0183413196
+ 5.53690774e-07 0.0167666634 5.53790774e-07 -0.0152403688 5.53890774e-07 0.0139298139 5.53990774e-07 -0.0126709058 5.54090774e-07 0.0115799054 5.54190774e-07 -0.0105396326 5.54290774e-07 0.00963120539 5.54390774e-07 -0.00877029031
+ 5.54490774e-07 0.00801373348 5.54590774e-07 -0.00730035533 5.54690774e-07 0.00667016991 5.54790774e-07 -0.0060784283 5.54890774e-07 0.00555342785 5.54990774e-07 -0.00506215822 5.55090774e-07 0.00462473134 5.55190774e-07 -0.00421658185
+ 5.55290774e-07 0.00385208255 5.55390774e-07 -0.0035127877 5.55490774e-07 0.00320903124 5.55590774e-07 -0.0029268357 5.55690774e-07 0.00267368149 5.55790774e-07 -0.00243887954 5.55890774e-07 0.00222788568 5.55990774e-07 -0.00203245084
+ 5.56090774e-07 0.0018565878 5.56190774e-07 -0.0016938733 5.56290774e-07 0.00154728638 5.56390774e-07 -0.00141178176 5.56490774e-07 0.00128959387 5.56590774e-07 -0.00117672642 5.56690774e-07 0.00107487425 5.56790774e-07 -0.000980846434
+ 5.56890774e-07 0.000895944254 5.56990774e-07 -0.000817600267 5.57090774e-07 0.000746826659 5.57190774e-07 -0.000681542527 5.57290774e-07 0.000622546127 5.57390774e-07 -0.000568139108 5.57490774e-07 0.000518960166 5.57590774e-07 -0.00047361387
+ 5.57690774e-07 0.000432618935 5.57790774e-07 -0.00039482136 5.57890774e-07 0.000360648892 5.57990774e-07 -0.000329141088 5.58090774e-07 0.000300656148 5.58190774e-07 -0.000274389641 5.58290774e-07 0.000250646154 5.58390774e-07 -0.000228747599
+ 5.58490774e-07 0.0002089569 5.58590774e-07 -0.000190698721 5.58690774e-07 0.000174203358 5.58790774e-07 -0.00015897934 5.58890774e-07 0.000145231232 5.58990774e-07 -0.000132536229 5.59090774e-07 0.000121078462 5.59190774e-07 -0.000110491511
+ 5.59290774e-07 0.000100943174 5.59390774e-07 -9.21134357e-05 5.59490774e-07 8.4156973e-05 5.59590774e-07 -7.67920397e-05 5.59690774e-07 7.01627124e-05 5.59790774e-07 -6.40188597e-05 5.59890774e-07 5.84959595e-05 5.59990774e-07 -5.33700348e-05
+ 5.60090774e-07 4.87695597e-05 5.60190774e-07 -4.44922222e-05 5.60290774e-07 4.06607716e-05 5.60390774e-07 -3.70908606e-05 5.60490774e-07 3.39005457e-05 5.60590774e-07 -3.09203885e-05 5.60690774e-07 2.82645887e-05 5.60790774e-07 -2.57760907e-05
+ 5.60890774e-07 2.3565917e-05 5.60990774e-07 -2.14873027e-05 5.61090774e-07 1.96486482e-05 5.61190774e-07 -1.79117455e-05 5.61290774e-07 1.63828276e-05 5.61390774e-07 -1.49308044e-05 5.61490774e-07 1.36601148e-05 5.61590774e-07 -1.24455918e-05
+ 5.61690774e-07 1.1390188e-05 5.61790774e-07 -1.03736667e-05 5.61890774e-07 9.49774736e-06 5.61990774e-07 -8.6462987e-06 5.62090774e-07 7.9200162e-06 5.62190774e-07 -7.20618766e-06 5.62290774e-07 6.60465801e-06 5.62390774e-07 -6.00556286e-06
+ 5.62490774e-07 5.50804017e-06 5.62590774e-07 -5.004598e-06 5.62690774e-07 4.59378634e-06 5.62790774e-07 -4.17008995e-06 5.62890774e-07 3.83156966e-06 5.62990774e-07 -3.47435733e-06 5.63090774e-07 3.19610667e-06 5.63190774e-07 -2.89432215e-06
+ 5.63290774e-07 2.66631855e-06 5.63390774e-07 -2.41074428e-06 5.63490774e-07 2.22463188e-06 5.63590774e-07 -2.00758319e-06 5.63690774e-07 1.85639569e-06 5.63790774e-07 -1.6714659e-06 5.63890774e-07 1.55939899e-06 5.63990774e-07 -1.38082138e-06
+ 5.64090774e-07 1.30227747e-06 5.64190774e-07 -1.14884092e-06 5.64290774e-07 1.08727392e-06 5.64390774e-07 -9.55390912e-07 5.64490774e-07 9.08044284e-07 5.64590774e-07 -7.94134405e-07 5.64690774e-07 7.58642143e-07 5.64790774e-07 -6.59714464e-07
+ 5.64890774e-07 6.34103635e-07 5.64990774e-07 -5.47664794e-07 5.65090774e-07 5.30290584e-07 5.65190774e-07 -4.54262083e-07 5.65290774e-07 4.43753895e-07 5.65390774e-07 -3.76403601e-07 5.65490774e-07 3.71618865e-07 5.65590774e-07 -3.11502551e-07
+ 5.65690774e-07 3.11488709e-07 5.65790774e-07 -2.57402481e-07 5.65890774e-07 2.61365519e-07 5.65990774e-07 -2.12307012e-07 5.66090774e-07 2.19586255e-07 5.66190774e-07 -1.74727651e-07 5.66290774e-07 1.84780202e-07 5.66390774e-07 -1.43421282e-07
+ 5.66490774e-07 1.55784187e-07 5.66590774e-07 -1.17340694e-07 5.66690774e-07 1.3162823e-07 5.66790774e-07 -9.56134645e-08 5.66890774e-07 1.11504324e-07 5.66990774e-07 -7.7512852e-08 5.67090774e-07 9.47394286e-08 5.67190774e-07 -6.2433646e-08
+ 5.67290774e-07 8.0773134e-08 5.67390774e-07 -4.98334141e-08 5.67490774e-07 6.90993794e-08 5.67590774e-07 -3.93732595e-08 5.67690774e-07 5.94152848e-08 5.67790774e-07 -3.06632475e-08 5.67890774e-07 5.13482988e-08 5.67990774e-07 -2.34074253e-08
+ 5.68090774e-07 4.4628163e-08 5.68190774e-07 -1.73630594e-08 5.68290774e-07 3.90298633e-08 5.68390774e-07 -1.23273488e-08 5.68490774e-07 3.43658604e-08 5.68590774e-07 -8.13252615e-09 5.68690774e-07 3.04809101e-08 5.68790774e-07 -4.63838568e-09
+ 5.68890774e-07 2.72448722e-08 5.68990774e-07 -1.72786987e-09 5.69090774e-07 2.45493397e-08 5.69190774e-07 6.96517788e-10 5.69290774e-07 2.23131569e-08 5.69390774e-07 2.70818365e-09 5.69490774e-07 2.04764042e-08 5.69590774e-07 4.36139963e-09
+ 5.69690774e-07 1.89668153e-08 5.69790774e-07 5.72018083e-09 5.69890774e-07 1.77260564e-08 5.69990774e-07 6.83700865e-09 5.70090774e-07 1.67062181e-08 5.70190774e-07 7.75499581e-09 5.70290774e-07 1.58679406e-08 5.70390774e-07 8.50956489e-09
+ 5.70490774e-07 1.50799959e-08 5.70590774e-07 9.11601342e-09 5.70690774e-07 1.45257672e-08 5.70790774e-07 9.61910654e-09 5.70890774e-07 1.40694267e-08 5.70990774e-07 1.00330061e-08 5.71090774e-07 1.36940245e-08 5.71190774e-07 1.03734907e-08
+ 5.71290774e-07 1.33852095e-08 5.71390774e-07 1.06535818e-08 5.71490774e-07 1.31311713e-08 5.71590774e-07 1.08839911e-08 5.71690774e-07 1.2922193e-08 5.71790774e-07 1.10735315e-08 5.71890774e-07 1.27502821e-08 5.71990774e-07 1.12294523e-08
+ 5.72090774e-07 1.26088636e-08 5.72190774e-07 1.13577175e-08 5.72290774e-07 1.24925286e-08 5.72390774e-07 1.14632323e-08 5.72490774e-07 1.23968277e-08 5.72590774e-07 1.15500322e-08 5.72690774e-07 1.23181004e-08 5.72790774e-07 1.16214377e-08
+ 5.72890774e-07 1.22533358e-08 5.72990774e-07 1.16801792e-08 5.73090774e-07 1.2200057e-08 5.73190774e-07 1.1728503e-08 5.73290774e-07 1.21562273e-08 5.73390774e-07 1.17682569e-08 5.73490774e-07 1.212017e-08 5.73590774e-07 1.18009615e-08
+ 5.73690774e-07 1.20905067e-08 5.73790774e-07 1.18278664e-08 5.73890774e-07 1.20661031e-08 5.73990774e-07 1.1850001e-08 5.74090774e-07 1.20460267e-08 5.74190774e-07 1.18682111e-08 5.74290774e-07 1.20295097e-08 5.74390774e-07 1.18831928e-08
+ 5.74490774e-07 1.20159206e-08 5.74590774e-07 1.18955186e-08 5.74690774e-07 1.20047404e-08 5.74790774e-07 1.19056593e-08 5.74890774e-07 1.19955423e-08 5.74990774e-07 1.1914003e-08 5.75090774e-07 1.19879739e-08 5.75190774e-07 1.19208679e-08
+ 5.75290774e-07 1.1981747e-08 5.75390774e-07 1.19265162e-08 5.75490774e-07 1.19766236e-08 5.75590774e-07 1.19311639e-08 5.75690774e-07 1.19724075e-08 5.75790774e-07 1.1934988e-08 5.75890774e-07 1.19689385e-08 5.75990774e-07 1.19381348e-08
+ 5.76090774e-07 1.1966084e-08 5.76190774e-07 1.19407247e-08 5.76290774e-07 1.19637345e-08 5.76390774e-07 1.19428558e-08 5.76490774e-07 1.19618012e-08 5.76590774e-07 1.19446095e-08 5.76690774e-07 1.19602105e-08 5.76790774e-07 1.19460527e-08
+ 5.76890774e-07 1.19589011e-08 5.76990774e-07 1.19472407e-08 5.77090774e-07 1.19578232e-08 5.77190774e-07 1.19482186e-08 5.77290774e-07 1.19569361e-08 5.77390774e-07 1.19490235e-08 5.77490774e-07 1.19562055e-08 5.77590774e-07 1.19496864e-08
+ 5.77690774e-07 1.19556043e-08 5.77790774e-07 1.19502318e-08 5.77890774e-07 1.19551091e-08 5.77990774e-07 1.19506812e-08 5.78090774e-07 1.19547013e-08 5.78190774e-07 1.19510512e-08 5.78290774e-07 1.19543659e-08 5.78390774e-07 1.19513556e-08
+ 5.78490774e-07 1.19540895e-08 5.78590774e-07 1.19516065e-08 5.78690774e-07 1.19538618e-08 5.78790774e-07 1.19518133e-08 5.78890774e-07 1.19536744e-08 5.78990774e-07 1.19519833e-08 5.79090774e-07 1.19535197e-08 5.79190774e-07 1.19521236e-08
+ 5.79290774e-07 1.19533923e-08 5.79390774e-07 1.19522393e-08 5.79490774e-07 1.19532873e-08 5.79590774e-07 1.19523345e-08 5.79690774e-07 1.19532005e-08 5.79790774e-07 1.19524136e-08 5.79890774e-07 1.19531291e-08 5.79990774e-07 1.19524783e-08
+ 5.80090774e-07 1.19530705e-08 5.80190774e-07 1.19525317e-08 5.80290774e-07 1.19530218e-08 5.80390774e-07 1.19525758e-08 5.80490774e-07 1.19529818e-08 5.80590774e-07 1.19526123e-08 5.80690774e-07 1.19529487e-08 5.80790774e-07 1.19526425e-08
+ 5.80890774e-07 1.19529213e-08 5.80990774e-07 1.19526671e-08 5.81090774e-07 1.19528987e-08 5.81190774e-07 1.19526877e-08 5.81290774e-07 1.19528798e-08 5.81390774e-07 1.19527051e-08 5.81490774e-07 1.19528645e-08 5.81590774e-07 1.19527188e-08
+ 5.81690774e-07 1.19528517e-08 5.81790774e-07 1.19527306e-08 5.81890774e-07 1.1952841e-08 5.81990774e-07 1.19527402e-08 5.82090774e-07 1.19528323e-08 5.82190774e-07 1.19527482e-08 5.82290774e-07 1.19528252e-08 5.82390774e-07 1.19527549e-08
+ 5.82490774e-07 1.19528191e-08 5.82590774e-07 1.19527603e-08 5.82690774e-07 1.19528143e-08 5.82790774e-07 1.19527648e-08 5.82890774e-07 1.19528102e-08 5.82990774e-07 1.19527686e-08 5.83090774e-07 1.19528064e-08 5.83190774e-07 1.19527718e-08
+ 5.83290774e-07 1.19528035e-08 5.83390774e-07 1.19527743e-08 5.83490774e-07 1.1952801e-08 5.83590774e-07 1.19527766e-08 5.83690774e-07 1.19527989e-08 5.83790774e-07 1.19527785e-08 5.83890774e-07 1.19527976e-08 5.83990774e-07 1.19527798e-08
+ 5.84090774e-07 1.19527963e-08 5.84190774e-07 1.19527812e-08 5.84290774e-07 1.19527949e-08 5.84390774e-07 1.19527823e-08 5.84490774e-07 1.19527937e-08 5.84590774e-07 1.1952783e-08 5.84690774e-07 1.19527931e-08 5.84790774e-07 1.1952784e-08
+ 5.84890774e-07 1.19527925e-08 5.84990774e-07 1.19527845e-08 5.85090774e-07 1.19527918e-08 5.85190774e-07 1.19527851e-08 5.85290774e-07 1.19527913e-08 5.85390774e-07 1.19527856e-08 5.85490774e-07 1.19527907e-08 5.85590774e-07 1.19527861e-08
+ 5.85690774e-07 1.19527904e-08 5.85790774e-07 1.19527865e-08 5.85890774e-07 1.19527903e-08 5.85990774e-07 1.19527867e-08 5.86090774e-07 1.19527897e-08 5.86190774e-07 1.1952787e-08 5.86290774e-07 1.19527898e-08 5.86390774e-07 1.19527871e-08
+ 5.86490774e-07 1.19527897e-08 5.86590774e-07 1.19527872e-08 5.86690774e-07 1.19527894e-08 5.86790774e-07 1.19527871e-08 5.86890774e-07 1.19527897e-08 5.86990774e-07 1.19527872e-08 5.87090774e-07 1.19527891e-08 5.87190774e-07 1.19527873e-08
+ 5.87290774e-07 1.19527894e-08 5.87390774e-07 1.19527874e-08 5.87490774e-07 1.1952789e-08 5.87590774e-07 1.19527875e-08 5.87690774e-07 1.1952789e-08 5.87790774e-07 1.19527877e-08 5.87890774e-07 1.19527891e-08 5.87990774e-07 1.19527877e-08
+ 5.88090774e-07 1.19527891e-08 5.88190774e-07 1.19527877e-08 5.88290774e-07 1.19527891e-08 5.88390774e-07 1.19527878e-08 5.88490774e-07 1.1952789e-08 5.88590774e-07 1.19527879e-08 5.88690774e-07 1.1952789e-08 5.88790774e-07 1.19527878e-08
+ 5.88890774e-07 1.19527888e-08 5.88990774e-07 1.19527878e-08 5.89090774e-07 1.1952789e-08 5.89190774e-07 1.19527879e-08 5.89290774e-07 1.19527889e-08 5.89390774e-07 1.1952788e-08 5.89490774e-07 1.19527889e-08 5.89590774e-07 1.19527879e-08
+ 5.89690774e-07 1.19527888e-08 5.89790774e-07 1.1952788e-08 5.89890774e-07 1.19527889e-08 5.89990774e-07 1.19527879e-08 5.90090774e-07 1.19527889e-08 5.90190774e-07 1.1952788e-08 5.90290774e-07 1.19527888e-08 5.90390774e-07 1.1952788e-08
+ 5.90490774e-07 1.19527887e-08 5.90590774e-07 1.19527881e-08 5.90690774e-07 1.19527888e-08 5.90790774e-07 1.19527881e-08 5.90890774e-07 1.19527887e-08 5.90990774e-07 1.19527882e-08 5.91090774e-07 1.19527886e-08 5.91190774e-07 1.19527882e-08
+ 5.91290774e-07 1.19527885e-08 5.91390774e-07 1.19527882e-08 5.91490774e-07 1.19527885e-08 5.91590774e-07 1.19527882e-08 5.91690774e-07 1.19527885e-08 5.91790774e-07 1.19527883e-08 5.91890774e-07 1.19527884e-08 5.91990774e-07 1.19527883e-08
+ 5.92090774e-07 1.19527885e-08 5.92190774e-07 1.19527883e-08 5.92290774e-07 1.19527884e-08 5.92390774e-07 1.19527883e-08 5.92490774e-07 1.19527885e-08 5.92590774e-07 1.19527883e-08 5.92690774e-07 1.19527885e-08 5.92790774e-07 1.19527883e-08
+ 5.92890774e-07 1.19527885e-08 5.92990774e-07 1.19527883e-08 5.93090774e-07 1.19527885e-08 5.93190774e-07 1.19527883e-08 5.93290774e-07 1.19527884e-08 5.93390774e-07 1.19527883e-08 5.93490774e-07 1.19527885e-08 5.93590774e-07 1.19527883e-08
+ 5.93690774e-07 1.19527885e-08 5.93790774e-07 1.19527883e-08 5.93890774e-07 1.19527885e-08 5.93990774e-07 1.19527883e-08 5.94090774e-07 1.19527885e-08 5.94190774e-07 1.19527883e-08 5.94290774e-07 1.19527885e-08 5.94390774e-07 1.19527883e-08
+ 5.94490774e-07 1.19527885e-08 5.94590774e-07 1.19527883e-08 5.94690774e-07 1.19527885e-08 5.94790774e-07 1.19527883e-08 5.94890774e-07 1.19527885e-08 5.94990774e-07 1.19527883e-08 5.95090774e-07 1.19527885e-08 5.95190774e-07 1.19527883e-08
+ 5.95290774e-07 1.19527885e-08 5.95390774e-07 1.19527883e-08 5.95490774e-07 1.19527885e-08 5.95590774e-07 1.19527883e-08 5.95690774e-07 1.19527885e-08 5.95790774e-07 1.19527883e-08 5.95890774e-07 1.19527885e-08 5.95990774e-07 1.19527883e-08
+ 5.96090774e-07 1.19527885e-08 5.96190774e-07 1.19527883e-08 5.96290774e-07 1.19527885e-08 5.96390774e-07 1.19527883e-08 5.96490774e-07 1.19527885e-08 5.96590774e-07 1.19527883e-08 5.96690774e-07 1.19527885e-08 5.96790774e-07 1.19527883e-08
+ 5.96890774e-07 1.19527885e-08 5.96990774e-07 1.19527883e-08 5.97090774e-07 1.19527885e-08 5.97190774e-07 1.19527883e-08 5.97290774e-07 1.19527885e-08 5.97390774e-07 1.19527883e-08 5.97490774e-07 1.19527885e-08 5.97590774e-07 1.19527883e-08
+ 5.97690774e-07 1.19527885e-08 5.97790774e-07 1.19527883e-08 5.97890774e-07 1.19527885e-08 5.97990774e-07 1.19527883e-08 5.98090774e-07 1.19527885e-08 5.98190774e-07 1.19527883e-08 5.98290774e-07 1.19527885e-08 5.98390774e-07 1.19527883e-08
+ 5.98490774e-07 1.19527885e-08 5.98590774e-07 1.19527883e-08 5.98690774e-07 1.19527885e-08 5.98790774e-07 1.19527883e-08 5.98890774e-07 1.19527885e-08 5.98990774e-07 1.19527883e-08 5.99090774e-07 1.19527885e-08 5.99190774e-07 1.19527883e-08
+ 5.99290774e-07 1.19527885e-08 5.99390774e-07 1.19527883e-08 5.99490774e-07 1.19527885e-08 5.99590774e-07 1.19527883e-08 5.99690774e-07 1.19527885e-08 5.99790774e-07 1.19527883e-08 5.99890774e-07 1.19527885e-08 5.99990774e-07 1.19527883e-08
+ 6e-07 1.19527881e-08 6.0001e-07 1.45272736e-08 6.0003e-07 1.23606658e-09 6.0007e-07 2.76445088e-08 6.0015e-07 -4.38735015e-09 6.0025e-07 2.82154677e-08 6.0035e-07 -3.18927074e-09 6.0045e-07 2.52177594e-08
+ 6.0055e-07 2.59408309e-09 6.0065e-07 -4.06359281e-08 6.0075e-07 3.06902814e-06 6.0085e-07 9.48375612e-05 6.00932239e-07 -0.0448088436 6.01e-07 1.97425329 6.01008502e-07 3.1007477 6.01025505e-07 4.14453646
+ 6.01059511e-07 4.88397722 6.01090728e-07 4.98064226 6.01143656e-07 5.00336705 6.01199398e-07 4.99900033 6.01276452e-07 5.00049859 6.01342062e-07 4.99975148 6.01411951e-07 5.00013732 6.01487979e-07 4.99991579
+ 6.01566956e-07 5.00005277 6.01643585e-07 4.99996651 6.01743585e-07 5.00002357 6.01843585e-07 4.9999831 6.01943585e-07 5.00001203 6.02043585e-07 4.99999123 6.02143585e-07 5.00000632 6.02243585e-07 4.99999529
+ 6.02343585e-07 5.00000343 6.02443585e-07 4.99999737 6.02543585e-07 5.00000193 6.02643585e-07 4.99999847 6.02743585e-07 5.00000113 6.02843585e-07 4.99999907 6.02943585e-07 5.00000068 6.03043585e-07 4.99999941
+ 6.03143585e-07 5.00000042 6.03243585e-07 4.99999961 6.03343585e-07 5.00000026 6.03443585e-07 4.99999974 6.03543585e-07 5.00000017 6.03643585e-07 4.99999981 6.03743585e-07 5.0000001 6.03843585e-07 4.99999986
+ 6.03943585e-07 5.00000006 6.04043585e-07 4.9999999 6.04143585e-07 5.00000003 6.04243585e-07 4.99999992 6.04343585e-07 5.00000001 6.04443585e-07 4.99999994 6.04543585e-07 5.0 6.04643585e-07 4.99999995
+ 6.04743585e-07 4.99999999 6.04843585e-07 4.99999996 6.04943585e-07 4.99999999 6.05043585e-07 4.99999996 6.05143585e-07 4.99999998 6.05243585e-07 4.99999996 6.05343585e-07 4.99999998 6.05443585e-07 4.99999997
+ 6.05543585e-07 4.99999998 6.05643585e-07 4.99999997 6.05743585e-07 4.99999998 6.05843585e-07 4.99999997 6.05943585e-07 4.99999997 6.06043585e-07 4.99999997 6.06143585e-07 4.99999997 6.06243585e-07 4.99999997
+ 6.06343585e-07 4.99999997 6.06443585e-07 4.99999997 6.06543585e-07 4.99999997 6.06643585e-07 4.99999997 6.06743585e-07 4.99999997 6.06843585e-07 4.99999997 6.06943585e-07 4.99999997 6.07043585e-07 4.99999997
+ 6.07143585e-07 4.99999997 6.07243585e-07 4.99999997 6.07343585e-07 4.99999997 6.07443585e-07 4.99999997 6.07543585e-07 4.99999997 6.07643585e-07 4.99999997 6.07743585e-07 4.99999997 6.07843585e-07 4.99999997
+ 6.07943585e-07 4.99999997 6.08043585e-07 4.99999997 6.08143585e-07 4.99999997 6.08243585e-07 4.99999997 6.08343585e-07 4.99999997 6.08443585e-07 4.99999997 6.08543585e-07 4.99999997 6.08643585e-07 4.99999997
+ 6.08743585e-07 4.99999997 6.08843585e-07 4.99999997 6.08943585e-07 4.99999997 6.09043585e-07 4.99999997 6.09143585e-07 4.99999997 6.09243585e-07 4.99999997 6.09343585e-07 4.99999997 6.09443585e-07 4.99999997
+ 6.09543585e-07 4.99999997 6.09643585e-07 4.99999997 6.09743585e-07 4.99999997 6.09843585e-07 4.99999997 6.09943585e-07 4.99999997 6.10043585e-07 4.99999997 6.10143585e-07 4.99999997 6.10243585e-07 4.99999997
+ 6.10343585e-07 4.99999997 6.10443585e-07 4.99999997 6.10543585e-07 4.99999997 6.10643585e-07 4.99999997 6.10743585e-07 4.99999997 6.10843585e-07 4.99999997 6.10943585e-07 4.99999997 6.11043585e-07 4.99999997
+ 6.11143585e-07 4.99999997 6.11243585e-07 4.99999997 6.11343585e-07 4.99999997 6.11443585e-07 4.99999997 6.11543585e-07 4.99999997 6.11643585e-07 4.99999997 6.11743585e-07 4.99999997 6.11843585e-07 4.99999997
+ 6.11943585e-07 4.99999997 6.12043585e-07 4.99999997 6.12143585e-07 4.99999997 6.12243585e-07 4.99999997 6.12343585e-07 4.99999997 6.12443585e-07 4.99999997 6.12543585e-07 4.99999997 6.12643585e-07 4.99999997
+ 6.12743585e-07 4.99999997 6.12843585e-07 4.99999997 6.12943585e-07 4.99999997 6.13043585e-07 4.99999997 6.13143585e-07 4.99999997 6.13243585e-07 4.99999997 6.13343585e-07 4.99999997 6.13443585e-07 4.99999997
+ 6.13543585e-07 4.99999997 6.13643585e-07 4.99999997 6.13743585e-07 4.99999997 6.13843585e-07 4.99999997 6.13943585e-07 4.99999997 6.14043585e-07 4.99999997 6.14143585e-07 4.99999997 6.14243585e-07 4.99999997
+ 6.14343585e-07 4.99999997 6.14443585e-07 4.99999997 6.14543585e-07 4.99999997 6.14643585e-07 4.99999997 6.14743585e-07 4.99999997 6.14843585e-07 4.99999997 6.14943585e-07 4.99999997 6.15043585e-07 4.99999997
+ 6.15143585e-07 4.99999997 6.15243585e-07 4.99999997 6.15343585e-07 4.99999997 6.15443585e-07 4.99999997 6.15543585e-07 4.99999997 6.15643585e-07 4.99999997 6.15743585e-07 4.99999997 6.15843585e-07 4.99999997
+ 6.15943585e-07 4.99999997 6.16043585e-07 4.99999997 6.16143585e-07 4.99999997 6.16243585e-07 4.99999997 6.16343585e-07 4.99999997 6.16443585e-07 4.99999997 6.16543585e-07 4.99999997 6.16643585e-07 4.99999997
+ 6.16743585e-07 4.99999997 6.16843585e-07 4.99999997 6.16943585e-07 4.99999997 6.17043585e-07 4.99999997 6.17143585e-07 4.99999997 6.17243585e-07 4.99999997 6.17343585e-07 4.99999997 6.17443585e-07 4.99999997
+ 6.17543585e-07 4.99999997 6.17643585e-07 4.99999997 6.17743585e-07 4.99999997 6.17843585e-07 4.99999997 6.17943585e-07 4.99999997 6.18043585e-07 4.99999997 6.18143585e-07 4.99999997 6.18243585e-07 4.99999997
+ 6.18343585e-07 4.99999997 6.18443585e-07 4.99999997 6.18543585e-07 4.99999997 6.18643585e-07 4.99999997 6.18743585e-07 4.99999997 6.18843585e-07 4.99999997 6.18943585e-07 4.99999997 6.19043585e-07 4.99999997
+ 6.19143585e-07 4.99999997 6.19243585e-07 4.99999997 6.19343585e-07 4.99999997 6.19443585e-07 4.99999997 6.19543585e-07 4.99999997 6.19643585e-07 4.99999997 6.19743585e-07 4.99999997 6.19843585e-07 4.99999997
+ 6.19943585e-07 4.99999997 6.20043585e-07 4.99999997 6.20143585e-07 4.99999997 6.20243585e-07 4.99999997 6.20343585e-07 4.99999997 6.20443585e-07 4.99999997 6.20543585e-07 4.99999997 6.20643585e-07 4.99999997
+ 6.20743585e-07 4.99999997 6.20843585e-07 4.99999997 6.20943585e-07 4.99999997 6.21043585e-07 4.99999997 6.21143585e-07 4.99999997 6.21243585e-07 4.99999997 6.21343585e-07 4.99999997 6.21443585e-07 4.99999997
+ 6.21543585e-07 4.99999997 6.21643585e-07 4.99999997 6.21743585e-07 4.99999997 6.21843585e-07 4.99999997 6.21943585e-07 4.99999997 6.22043585e-07 4.99999997 6.22143585e-07 4.99999997 6.22243585e-07 4.99999997
+ 6.22343585e-07 4.99999997 6.22443585e-07 4.99999997 6.22543585e-07 4.99999997 6.22643585e-07 4.99999997 6.22743585e-07 4.99999997 6.22843585e-07 4.99999997 6.22943585e-07 4.99999997 6.23043585e-07 4.99999997
+ 6.23143585e-07 4.99999997 6.23243585e-07 4.99999997 6.23343585e-07 4.99999997 6.23443585e-07 4.99999997 6.23543585e-07 4.99999997 6.23643585e-07 4.99999997 6.23743585e-07 4.99999997 6.23843585e-07 4.99999997
+ 6.23943585e-07 4.99999997 6.24043585e-07 4.99999997 6.24143585e-07 4.99999997 6.24243585e-07 4.99999997 6.24343585e-07 4.99999997 6.24443585e-07 4.99999997 6.24543585e-07 4.99999997 6.24643585e-07 4.99999997
+ 6.24743585e-07 4.99999997 6.24843585e-07 4.99999997 6.24943585e-07 4.99999997 6.25043585e-07 4.99999997 6.25143585e-07 4.99999997 6.25243585e-07 4.99999997 6.25343585e-07 4.99999997 6.25443585e-07 4.99999997
+ 6.25543585e-07 4.99999997 6.25643585e-07 4.99999997 6.25743585e-07 4.99999997 6.25843585e-07 4.99999997 6.25943585e-07 4.99999997 6.26043585e-07 4.99999997 6.26143585e-07 4.99999997 6.26243585e-07 4.99999997
+ 6.26343585e-07 4.99999997 6.26443585e-07 4.99999997 6.26543585e-07 4.99999997 6.26643585e-07 4.99999997 6.26743585e-07 4.99999997 6.26843585e-07 4.99999997 6.26943585e-07 4.99999997 6.27043585e-07 4.99999997
+ 6.27143585e-07 4.99999997 6.27243585e-07 4.99999997 6.27343585e-07 4.99999997 6.27443585e-07 4.99999997 6.27543585e-07 4.99999997 6.27643585e-07 4.99999997 6.27743585e-07 4.99999997 6.27843585e-07 4.99999997
+ 6.27943585e-07 4.99999997 6.28043585e-07 4.99999997 6.28143585e-07 4.99999997 6.28243585e-07 4.99999997 6.28343585e-07 4.99999997 6.28443585e-07 4.99999997 6.28543585e-07 4.99999997 6.28643585e-07 4.99999997
+ 6.28743585e-07 4.99999997 6.28843585e-07 4.99999997 6.28943585e-07 4.99999997 6.29043585e-07 4.99999997 6.29143585e-07 4.99999997 6.29243585e-07 4.99999997 6.29343585e-07 4.99999997 6.29443585e-07 4.99999997
+ 6.29543585e-07 4.99999997 6.29643585e-07 4.99999997 6.29743585e-07 4.99999997 6.29843585e-07 4.99999997 6.29943585e-07 4.99999997 6.30043585e-07 4.99999997 6.30143585e-07 4.99999997 6.30243585e-07 4.99999997
+ 6.30343585e-07 4.99999997 6.30443585e-07 4.99999997 6.30543585e-07 4.99999997 6.30643585e-07 4.99999997 6.30743585e-07 4.99999997 6.30843585e-07 4.99999997 6.30943585e-07 4.99999997 6.31043585e-07 4.99999997
+ 6.31143585e-07 4.99999997 6.31243585e-07 4.99999997 6.31343585e-07 4.99999997 6.31443585e-07 4.99999997 6.31543585e-07 4.99999997 6.31643585e-07 4.99999997 6.31743585e-07 4.99999997 6.31843585e-07 4.99999997
+ 6.31943585e-07 4.99999997 6.32043585e-07 4.99999997 6.32143585e-07 4.99999997 6.32243585e-07 4.99999997 6.32343585e-07 4.99999997 6.32443585e-07 4.99999997 6.32543585e-07 4.99999997 6.32643585e-07 4.99999997
+ 6.32743585e-07 4.99999997 6.32843585e-07 4.99999997 6.32943585e-07 4.99999997 6.33043585e-07 4.99999997 6.33143585e-07 4.99999997 6.33243585e-07 4.99999997 6.33343585e-07 4.99999997 6.33443585e-07 4.99999997
+ 6.33543585e-07 4.99999997 6.33643585e-07 4.99999997 6.33743585e-07 4.99999997 6.33843585e-07 4.99999997 6.33943585e-07 4.99999997 6.34043585e-07 4.99999997 6.34143585e-07 4.99999997 6.34243585e-07 4.99999997
+ 6.34343585e-07 4.99999997 6.34443585e-07 4.99999997 6.34543585e-07 4.99999997 6.34643585e-07 4.99999997 6.34743585e-07 4.99999997 6.34843585e-07 4.99999997 6.34943585e-07 4.99999997 6.35043585e-07 4.99999997
+ 6.35143585e-07 4.99999997 6.35243585e-07 4.99999997 6.35343585e-07 4.99999997 6.35443585e-07 4.99999997 6.35543585e-07 4.99999997 6.35643585e-07 4.99999997 6.35743585e-07 4.99999997 6.35843585e-07 4.99999997
+ 6.35943585e-07 4.99999997 6.36043585e-07 4.99999997 6.36143585e-07 4.99999997 6.36243585e-07 4.99999997 6.36343585e-07 4.99999997 6.36443585e-07 4.99999997 6.36543585e-07 4.99999997 6.36643585e-07 4.99999997
+ 6.36743585e-07 4.99999997 6.36843585e-07 4.99999997 6.36943585e-07 4.99999997 6.37043585e-07 4.99999997 6.37143585e-07 4.99999997 6.37243585e-07 4.99999997 6.37343585e-07 4.99999997 6.37443585e-07 4.99999997
+ 6.37543585e-07 4.99999997 6.37643585e-07 4.99999997 6.37743585e-07 4.99999997 6.37843585e-07 4.99999997 6.37943585e-07 4.99999997 6.38043585e-07 4.99999997 6.38143585e-07 4.99999997 6.38243585e-07 4.99999997
+ 6.38343585e-07 4.99999997 6.38443585e-07 4.99999997 6.38543585e-07 4.99999997 6.38643585e-07 4.99999997 6.38743585e-07 4.99999997 6.38843585e-07 4.99999997 6.38943585e-07 4.99999997 6.39043585e-07 4.99999997
+ 6.39143585e-07 4.99999997 6.39243585e-07 4.99999997 6.39343585e-07 4.99999997 6.39443585e-07 4.99999997 6.39543585e-07 4.99999997 6.39643585e-07 4.99999997 6.39743585e-07 4.99999997 6.39843585e-07 4.99999997
+ 6.39943585e-07 4.99999997 6.40043585e-07 4.99999997 6.40143585e-07 4.99999997 6.40243585e-07 4.99999997 6.40343585e-07 4.99999997 6.40443585e-07 4.99999997 6.40543585e-07 4.99999997 6.40643585e-07 4.99999997
+ 6.40743585e-07 4.99999997 6.40843585e-07 4.99999997 6.40943585e-07 4.99999997 6.41043585e-07 4.99999997 6.41143585e-07 4.99999997 6.41243585e-07 4.99999997 6.41343585e-07 4.99999997 6.41443585e-07 4.99999997
+ 6.41543585e-07 4.99999997 6.41643585e-07 4.99999997 6.41743585e-07 4.99999997 6.41843585e-07 4.99999997 6.41943585e-07 4.99999997 6.42043585e-07 4.99999997 6.42143585e-07 4.99999997 6.42243585e-07 4.99999997
+ 6.42343585e-07 4.99999997 6.42443585e-07 4.99999997 6.42543585e-07 4.99999997 6.42643585e-07 4.99999997 6.42743585e-07 4.99999997 6.42843585e-07 4.99999997 6.42943585e-07 4.99999997 6.43043585e-07 4.99999997
+ 6.43143585e-07 4.99999997 6.43243585e-07 4.99999997 6.43343585e-07 4.99999997 6.43443585e-07 4.99999997 6.43543585e-07 4.99999997 6.43643585e-07 4.99999997 6.43743585e-07 4.99999997 6.43843585e-07 4.99999997
+ 6.43943585e-07 4.99999997 6.44043585e-07 4.99999997 6.44143585e-07 4.99999997 6.44243585e-07 4.99999997 6.44343585e-07 4.99999997 6.44443585e-07 4.99999997 6.44543585e-07 4.99999997 6.44643585e-07 4.99999997
+ 6.44743585e-07 4.99999997 6.44843585e-07 4.99999997 6.44943585e-07 4.99999997 6.45043585e-07 4.99999997 6.45143585e-07 4.99999997 6.45243585e-07 4.99999997 6.45343585e-07 4.99999997 6.45443585e-07 4.99999997
+ 6.45543585e-07 4.99999997 6.45643585e-07 4.99999997 6.45743585e-07 4.99999997 6.45843585e-07 4.99999997 6.45943585e-07 4.99999997 6.46043585e-07 4.99999997 6.46143585e-07 4.99999997 6.46243585e-07 4.99999997
+ 6.46343585e-07 4.99999997 6.46443585e-07 4.99999997 6.46543585e-07 4.99999997 6.46643585e-07 4.99999997 6.46743585e-07 4.99999997 6.46843585e-07 4.99999997 6.46943585e-07 4.99999997 6.47043585e-07 4.99999997
+ 6.47143585e-07 4.99999997 6.47243585e-07 4.99999997 6.47343585e-07 4.99999997 6.47443585e-07 4.99999997 6.47543585e-07 4.99999997 6.47643585e-07 4.99999997 6.47743585e-07 4.99999997 6.47843585e-07 4.99999997
+ 6.47943585e-07 4.99999997 6.48043585e-07 4.99999997 6.48143585e-07 4.99999997 6.48243585e-07 4.99999997 6.48343585e-07 4.99999997 6.48443585e-07 4.99999997 6.48543585e-07 4.99999997 6.48643585e-07 4.99999997
+ 6.48743585e-07 4.99999997 6.48843585e-07 4.99999997 6.48943585e-07 4.99999997 6.49043585e-07 4.99999997 6.49143585e-07 4.99999997 6.49243585e-07 4.99999997 6.49343585e-07 4.99999997 6.49443585e-07 4.99999997
+ 6.49543585e-07 4.99999997 6.49643585e-07 4.99999997 6.49743585e-07 4.99999997 6.49843585e-07 4.99999997 6.49943585e-07 4.99999997 6.50043585e-07 4.99999997 6.50143585e-07 4.99999997 6.50243585e-07 4.99999997
+ 6.50343585e-07 4.99999997 6.50443585e-07 4.99999997 6.50543585e-07 4.99999997 6.50643585e-07 4.99999997 6.50743585e-07 4.99999997 6.50843585e-07 4.99999997 6.50943585e-07 4.99999997 6.51e-07 4.99999997
+ 6.5101e-07 4.99999997 6.5103e-07 4.99999998 6.5107e-07 4.99999996 6.5115e-07 4.99999998 6.5125e-07 4.99999997 6.5135e-07 4.99999997 6.5145e-07 4.99999998 6.5155e-07 4.99999996
+ 6.5165e-07 4.99999998 6.5175e-07 4.99999996 6.5185e-07 4.99999999 6.51930828e-07 5.00006476 6.52e-07 4.99916064 6.52008608e-07 4.99761638 6.52025825e-07 4.99311194 6.52060258e-07 5.01027326
+ 6.52106181e-07 5.09906166 6.52150081e-07 4.21228987 6.52198026e-07 0.290284563 6.5225538e-07 -0.0554589573 6.52312019e-07 0.0719466825 6.52404231e-07 -0.0579814231 6.52504231e-07 0.052890252 6.52604231e-07 -0.0475728397
+ 6.52704231e-07 0.0435755801 6.52804231e-07 -0.0393282951 6.52904231e-07 0.0359988053 6.53004231e-07 -0.0325571519 6.53104231e-07 0.029786221 6.53204231e-07 -0.0269830488 6.53304231e-07 0.0246778153 6.53404231e-07 -0.0223853345
+ 6.53504231e-07 0.0204675598 6.53604231e-07 -0.0185864689 6.53704231e-07 0.0169907803 6.53804231e-07 -0.0154430156 6.53904231e-07 0.0141150275 6.54004231e-07 -0.0128386436 6.54104231e-07 0.0117331852 6.54204231e-07 -0.0106786325
+ 6.54304231e-07 0.00975820759 6.54404231e-07 -0.00888558601 6.54504231e-07 0.00811906716 6.54604231e-07 -0.00739606596 6.54704231e-07 0.00675760434 6.54804231e-07 -0.00615793428 6.54904231e-07 0.00562605481 6.55004231e-07 -0.00512824045
+ 6.55104231e-07 0.00468509345 6.55204231e-07 -0.0042715328 6.55304231e-07 0.00390227528 6.55404231e-07 -0.00355850054 6.55504231e-07 0.00325078477 6.55604231e-07 -0.00296487618 6.55704231e-07 0.00270842653 6.55804231e-07 -0.00247054424
+ 6.55904231e-07 0.00225680687 6.56004231e-07 -0.00205881459 6.56104231e-07 0.00188066709 6.56204231e-07 -0.0017158279 6.56304231e-07 0.00156733843 6.56404231e-07 -0.00143006768 6.56504231e-07 0.00130629509 6.56604231e-07 -0.00119195888
+ 6.56704231e-07 0.0010887866 6.56804231e-07 -0.000993536867 6.56904231e-07 0.000907534878 6.57004231e-07 -0.000828173997 6.57104231e-07 0.000756484035 6.57204231e-07 -0.000690353405 6.57304231e-07 0.000630593448 6.57404231e-07 -0.000575481614
+ 6.57504231e-07 0.000525666393 6.57604231e-07 -0.000479733137 6.57704231e-07 0.000438207956 6.57804231e-07 -0.00039992149 6.57904231e-07 0.000365307115 6.58004231e-07 -0.000333392049 6.58104231e-07 0.000304538809 6.58204231e-07 -0.000277932999
+ 6.58304231e-07 0.000253882545 6.58404231e-07 -0.000231701277 6.58504231e-07 0.000211654724 6.58604231e-07 -0.000193160962 6.58704231e-07 0.000176452339 6.58804231e-07 -0.000161031999 6.58904231e-07 0.000147106127 6.59004231e-07 -0.000134247508
+ 6.59104231e-07 0.000122641562 6.59204231e-07 -0.000111918243 6.59304231e-07 0.000102246385 6.59404231e-07 -9.33029846e-05 6.59504231e-07 8.52435523e-05 6.59604231e-07 -7.77838768e-05 6.59704231e-07 7.10687098e-05 6.59804231e-07 -6.4845882e-05
+ 6.59904231e-07 5.925142e-05 6.60004231e-07 -5.40596605e-05 6.60104231e-07 4.93995251e-05 6.60204231e-07 -4.50673043e-05 6.60304231e-07 4.11861142e-05 6.60404231e-07 -3.75704478e-05 6.60504231e-07 3.4338663e-05 6.60604231e-07 -3.13203588e-05
+ 6.60704231e-07 2.86299828e-05 6.60804231e-07 -2.61096797e-05 6.60904231e-07 2.38706765e-05 6.61004231e-07 -2.17655435e-05 6.61104231e-07 1.99028504e-05 6.61204231e-07 -1.81438359e-05 6.61304231e-07 1.65948732e-05 6.61404231e-07 -1.5124412e-05
+ 6.61504231e-07 1.38370073e-05 6.61604231e-07 -1.26071091e-05 6.61704231e-07 1.15377661e-05 6.61804231e-07 -1.0508423e-05 6.61904231e-07 9.62087887e-06 6.62004231e-07 -8.75873714e-06 6.62104231e-07 8.02275961e-06 6.62204231e-07 -7.3000129e-06
+ 6.62304231e-07 6.69039716e-06 6.62404231e-07 -6.08386372e-06 6.62504231e-07 5.5795965e-06 6.62604231e-07 -5.06994998e-06 6.62704231e-07 4.65351243e-06 6.62804231e-07 -4.22464061e-06 6.62904231e-07 3.88142724e-06 6.63004231e-07 -3.51989747e-06
+ 6.63104231e-07 3.2377316e-06 6.63204231e-07 -2.93234513e-06 6.63304231e-07 2.70107501e-06 6.63404231e-07 -2.44249547e-06 6.63504231e-07 2.25365756e-06 6.63604231e-07 -2.03410123e-06 6.63704231e-07 1.88063941e-06 6.63804231e-07 -1.693617e-06
+ 6.63904231e-07 1.56964859e-06 6.64004231e-07 -1.40079315e-06 6.64104231e-07 1.32022001e-06 6.64204231e-07 -1.16494992e-06 6.64304231e-07 1.10220937e-06 6.64404231e-07 -9.68844208e-07 6.64504231e-07 9.20524047e-07 6.64604231e-07 -8.05377433e-07
+ 6.64704231e-07 7.69072859e-07 6.64804231e-07 -6.69112641e-07 6.64904231e-07 6.42823883e-07 6.65004231e-07 -5.55522921e-07 6.65104231e-07 5.37583103e-07 6.65204231e-07 -4.60834721e-07 6.65304231e-07 4.49854148e-07 6.65404231e-07 -3.81902181e-07
+ 6.65504231e-07 3.76722907e-07 6.65604231e-07 -3.16103905e-07 6.65704231e-07 3.15760619e-07 6.65804231e-07 -2.61254327e-07 6.65904231e-07 2.64942218e-07 6.66004231e-07 -2.15531651e-07 6.66104231e-07 2.22580083e-07 6.66204231e-07 -1.77427235e-07
+ 6.66304231e-07 1.87287055e-07 6.66404231e-07 -1.45682225e-07 6.66504231e-07 1.57884166e-07 6.66604231e-07 -1.192351e-07 6.66704231e-07 1.33388171e-07 6.66804231e-07 -9.72015e-08 6.66904231e-07 1.12980002e-07 6.67004231e-07 -7.88447312e-08
+ 6.67104231e-07 9.59773838e-08 6.67204231e-07 -6.35512259e-08 6.67304231e-07 8.18121369e-08 6.67404231e-07 -5.07714673e-08 6.67504231e-07 6.99716868e-08 6.67604231e-07 -4.01611717e-08 6.67704231e-07 6.01481946e-08 6.67804231e-07 -3.13254486e-08
+ 6.67904231e-07 5.19644651e-08 6.68004231e-07 -2.39643281e-08 6.68104231e-07 4.51465265e-08 6.68204231e-07 -1.78317312e-08 6.68304231e-07 3.94662537e-08 6.68404231e-07 -1.27220455e-08 6.68504231e-07 3.47335097e-08 6.68604231e-07 -8.4651863e-09
+ 6.68704231e-07 3.07909066e-08 6.68804231e-07 -4.91900451e-09 6.68904231e-07 2.75064927e-08 6.69004231e-07 -1.96481137e-09 6.69104231e-07 2.47703488e-08 6.69204231e-07 4.96254204e-10 6.69304231e-07 2.24974266e-08 6.69404231e-07 2.54098009e-09
+ 6.69504231e-07 2.06303728e-08 6.69604231e-07 4.22158863e-09 6.69704231e-07 1.90956559e-08 6.69804231e-07 5.60309754e-09 6.69904231e-07 1.78340381e-08 6.70004231e-07 6.73880063e-09 6.70104231e-07 1.67968683e-08 6.70204231e-07 7.67247987e-09
+ 6.70304231e-07 1.59441738e-08 6.70404231e-07 8.44010867e-09 6.70504231e-07 1.51438051e-08 6.70604231e-07 9.05738062e-09 6.70704231e-07 1.45796681e-08 6.70804231e-07 9.56953086e-09 6.70904231e-07 1.41150475e-08 6.71004231e-07 9.99100255e-09
+ 6.71104231e-07 1.37327182e-08 6.71204231e-07 1.03378268e-08 6.71304231e-07 1.34180995e-08 6.71404231e-07 1.06232328e-08 6.71504231e-07 1.31591913e-08 6.71604231e-07 1.08581058e-08 6.71704231e-07 1.29461201e-08 6.71804231e-07 1.10514011e-08
+ 6.71904231e-07 1.27707631e-08 6.72004231e-07 1.12104866e-08 6.72104231e-07 1.26264374e-08 6.72204231e-07 1.13414235e-08 6.72304231e-07 1.25076454e-08 6.72404231e-07 1.1449199e-08 6.72504231e-07 1.24098633e-08 6.72604231e-07 1.15379161e-08
+ 6.72704231e-07 1.23293694e-08 6.72804231e-07 1.16109497e-08 6.72904231e-07 1.22631032e-08 6.73004231e-07 1.16710778e-08 6.73104231e-07 1.22085437e-08 6.73204231e-07 1.17205851e-08 6.73304231e-07 1.21636197e-08 6.73404231e-07 1.17613514e-08
+ 6.73504231e-07 1.21266251e-08 6.73604231e-07 1.17949241e-08 6.73704231e-07 1.20961567e-08 6.73804231e-07 1.18225762e-08 6.73904231e-07 1.207106e-08 6.74004231e-07 1.18453544e-08 6.74104231e-07 1.20503851e-08 6.74204231e-07 1.18641205e-08
+ 6.74304231e-07 1.20333505e-08 6.74404231e-07 1.18795842e-08 6.74504231e-07 1.20193127e-08 6.74604231e-07 1.18923286e-08 6.74704231e-07 1.2007742e-08 6.74804231e-07 1.19028339e-08 6.74904231e-07 1.19982031e-08 6.75004231e-07 1.19114958e-08
+ 6.75104231e-07 1.19903374e-08 6.75204231e-07 1.19186389e-08 6.75304231e-07 1.19838498e-08 6.75404231e-07 1.19245313e-08 6.75504231e-07 1.19784976e-08 6.75604231e-07 1.19293935e-08 6.75704231e-07 1.19740805e-08 6.75804231e-07 1.19334068e-08
+ 6.75904231e-07 1.1970434e-08 6.76004231e-07 1.19367204e-08 6.76104231e-07 1.19674223e-08 6.76204231e-07 1.19394575e-08 6.76304231e-07 1.19649342e-08 6.76404231e-07 1.19417194e-08 6.76504231e-07 1.19628779e-08 6.76604231e-07 1.19435894e-08
+ 6.76704231e-07 1.19611773e-08 6.76804231e-07 1.19451362e-08 6.76904231e-07 1.19597701e-08 6.77004231e-07 1.19464165e-08 6.77104231e-07 1.19586052e-08 6.77204231e-07 1.19474764e-08 6.77304231e-07 1.19576405e-08 6.77404231e-07 1.19483549e-08
+ 6.77504231e-07 1.19568404e-08 6.77604231e-07 1.19490833e-08 6.77704231e-07 1.1956177e-08 6.77804231e-07 1.1949688e-08 6.77904231e-07 1.1955626e-08 6.78004231e-07 1.19501898e-08 6.78104231e-07 1.19551684e-08 6.78204231e-07 1.19506072e-08
+ 6.78304231e-07 1.19547877e-08 6.78404231e-07 1.19509546e-08 6.78504231e-07 1.19544707e-08 6.78604231e-07 1.19512439e-08 6.78704231e-07 1.19542066e-08 6.78804231e-07 1.19514852e-08 6.78904231e-07 1.19539859e-08 6.79004231e-07 1.19516868e-08
+ 6.79104231e-07 1.19538021e-08 6.79204231e-07 1.19518552e-08 6.79304231e-07 1.19536477e-08 6.79404231e-07 1.19519963e-08 6.79504231e-07 1.19535188e-08 6.79604231e-07 1.19521143e-08 6.79704231e-07 1.19534103e-08 6.79804231e-07 1.19522136e-08
+ 6.79904231e-07 1.19533192e-08 6.80004231e-07 1.19522975e-08 6.80104231e-07 1.19532427e-08 6.80204231e-07 1.19523677e-08 6.80304231e-07 1.19531781e-08 6.80404231e-07 1.1952427e-08 6.80504231e-07 1.19531235e-08 6.80604231e-07 1.19524772e-08
+ 6.80704231e-07 1.19530771e-08 6.80804231e-07 1.19525199e-08 6.80904231e-07 1.19530381e-08 6.81004231e-07 1.19525559e-08 6.81104231e-07 1.19530049e-08 6.81204231e-07 1.19525865e-08 6.81304231e-07 1.19529765e-08 6.81404231e-07 1.1952613e-08
+ 6.81504231e-07 1.19529518e-08 6.81604231e-07 1.19526357e-08 6.81704231e-07 1.19529311e-08 6.81804231e-07 1.19526548e-08 6.81904231e-07 1.19529132e-08 6.82004231e-07 1.19526713e-08 6.82104231e-07 1.19528979e-08 6.82204231e-07 1.19526857e-08
+ 6.82304231e-07 1.19528845e-08 6.82404231e-07 1.19526981e-08 6.82504231e-07 1.1952873e-08 6.82604231e-07 1.19527087e-08 6.82704231e-07 1.19528631e-08 6.82804231e-07 1.19527177e-08 6.82904231e-07 1.19528546e-08 6.83004231e-07 1.19527261e-08
+ 6.83104231e-07 1.19528468e-08 6.83204231e-07 1.1952733e-08 6.83304231e-07 1.19528402e-08 6.83404231e-07 1.19527394e-08 6.83504231e-07 1.19528344e-08 6.83604231e-07 1.1952745e-08 6.83704231e-07 1.19528293e-08 6.83804231e-07 1.19527495e-08
+ 6.83904231e-07 1.19528252e-08 6.84004231e-07 1.19527538e-08 6.84104231e-07 1.19528209e-08 6.84204231e-07 1.19527573e-08 6.84304231e-07 1.19528176e-08 6.84404231e-07 1.19527606e-08 6.84504231e-07 1.19528146e-08 6.84604231e-07 1.19527635e-08
+ 6.84704231e-07 1.19528116e-08 6.84804231e-07 1.19527659e-08 6.84904231e-07 1.19528095e-08 6.85004231e-07 1.19527684e-08 6.85104231e-07 1.19528072e-08 6.85204231e-07 1.19527702e-08 6.85304231e-07 1.19528054e-08 6.85404231e-07 1.1952772e-08
+ 6.85504231e-07 1.19528036e-08 6.85604231e-07 1.19527738e-08 6.85704231e-07 1.19528021e-08 6.85804231e-07 1.19527753e-08 6.85904231e-07 1.19528006e-08 6.86004231e-07 1.19527763e-08 6.86104231e-07 1.19527997e-08 6.86204231e-07 1.19527777e-08
+ 6.86304231e-07 1.19527986e-08 6.86404231e-07 1.19527785e-08 6.86504231e-07 1.19527976e-08 6.86604231e-07 1.19527795e-08 6.86704231e-07 1.19527966e-08 6.86804231e-07 1.19527805e-08 6.86904231e-07 1.19527955e-08 6.87004231e-07 1.19527813e-08
+ 6.87104231e-07 1.19527948e-08 6.87204231e-07 1.19527821e-08 6.87304231e-07 1.19527942e-08 6.87404231e-07 1.19527828e-08 6.87504231e-07 1.19527936e-08 6.87604231e-07 1.19527831e-08 6.87704231e-07 1.19527933e-08 6.87804231e-07 1.19527835e-08
+ 6.87904231e-07 1.19527929e-08 6.88004231e-07 1.19527842e-08 6.88104231e-07 1.19527924e-08 6.88204231e-07 1.19527844e-08 6.88304231e-07 1.19527919e-08 6.88404231e-07 1.19527848e-08 6.88504231e-07 1.19527918e-08 6.88604231e-07 1.19527851e-08
+ 6.88704231e-07 1.19527915e-08 6.88804231e-07 1.19527854e-08 6.88904231e-07 1.1952791e-08 6.89004231e-07 1.19527858e-08 6.89104231e-07 1.19527906e-08 6.89204231e-07 1.1952786e-08 6.89304231e-07 1.19527906e-08 6.89404231e-07 1.19527863e-08
+ 6.89504231e-07 1.19527901e-08 6.89604231e-07 1.19527865e-08 6.89704231e-07 1.19527899e-08 6.89804231e-07 1.19527868e-08 6.89904231e-07 1.19527898e-08 6.90004231e-07 1.19527869e-08 6.90104231e-07 1.19527897e-08 6.90204231e-07 1.19527868e-08
+ 6.90304231e-07 1.19527897e-08 6.90404231e-07 1.19527869e-08 6.90504231e-07 1.19527898e-08 6.90604231e-07 1.1952787e-08 6.90704231e-07 1.19527898e-08 6.90804231e-07 1.19527871e-08 6.90904231e-07 1.19527897e-08 6.91004231e-07 1.1952787e-08
+ 6.91104231e-07 1.19527894e-08 6.91204231e-07 1.19527872e-08 6.91304231e-07 1.19527894e-08 6.91404231e-07 1.19527872e-08 6.91504231e-07 1.19527896e-08 6.91604231e-07 1.19527872e-08 6.91704231e-07 1.19527893e-08 6.91804231e-07 1.19527872e-08
+ 6.91904231e-07 1.19527894e-08 6.92004231e-07 1.19527874e-08 6.92104231e-07 1.1952789e-08 6.92204231e-07 1.19527874e-08 6.92304231e-07 1.19527892e-08 6.92404231e-07 1.19527876e-08 6.92504231e-07 1.19527892e-08 6.92604231e-07 1.19527876e-08
+ 6.92704231e-07 1.1952789e-08 6.92804231e-07 1.19527876e-08 6.92904231e-07 1.1952789e-08 6.93004231e-07 1.19527876e-08 6.93104231e-07 1.1952789e-08 6.93204231e-07 1.19527878e-08 6.93304231e-07 1.19527889e-08 6.93404231e-07 1.19527879e-08
+ 6.93504231e-07 1.1952789e-08 6.93604231e-07 1.19527879e-08 6.93704231e-07 1.19527889e-08 6.93804231e-07 1.1952788e-08 6.93904231e-07 1.19527888e-08 6.94004231e-07 1.1952788e-08 6.94104231e-07 1.19527888e-08 6.94204231e-07 1.1952788e-08
+ 6.94304231e-07 1.19527888e-08 6.94404231e-07 1.1952788e-08 6.94504231e-07 1.19527889e-08 6.94604231e-07 1.1952788e-08 6.94704231e-07 1.19527886e-08 6.94804231e-07 1.1952788e-08 6.94904231e-07 1.19527888e-08 6.95004231e-07 1.1952788e-08
+ 6.95104231e-07 1.19527887e-08 6.95204231e-07 1.19527881e-08 6.95304231e-07 1.19527887e-08 6.95404231e-07 1.19527881e-08 6.95504231e-07 1.19527886e-08 6.95604231e-07 1.19527881e-08 6.95704231e-07 1.19527887e-08 6.95804231e-07 1.19527881e-08
+ 6.95904231e-07 1.19527886e-08 6.96004231e-07 1.19527882e-08 6.96104231e-07 1.19527885e-08 6.96204231e-07 1.19527882e-08 6.96304231e-07 1.19527885e-08 6.96404231e-07 1.19527882e-08 6.96504231e-07 1.19527885e-08 6.96604231e-07 1.19527882e-08
+ 6.96704231e-07 1.19527885e-08 6.96804231e-07 1.19527882e-08 6.96904231e-07 1.19527885e-08 6.97004231e-07 1.19527882e-08 6.97104231e-07 1.19527885e-08 6.97204231e-07 1.19527882e-08 6.97304231e-07 1.19527885e-08 6.97404231e-07 1.19527883e-08
+ 6.97504231e-07 1.19527884e-08 6.97604231e-07 1.19527883e-08 6.97704231e-07 1.19527885e-08 6.97804231e-07 1.19527883e-08 6.97904231e-07 1.19527885e-08 6.98004231e-07 1.19527883e-08 6.98104231e-07 1.19527885e-08 6.98204231e-07 1.19527883e-08
+ 6.98304231e-07 1.19527885e-08 6.98404231e-07 1.19527883e-08 6.98504231e-07 1.19527885e-08 6.98604231e-07 1.19527883e-08 6.98704231e-07 1.19527885e-08 6.98804231e-07 1.19527883e-08 6.98904231e-07 1.19527885e-08 6.99004231e-07 1.19527883e-08
+ 6.99104231e-07 1.19527885e-08 6.99204231e-07 1.19527883e-08 6.99304231e-07 1.19527885e-08 6.99404231e-07 1.19527883e-08 6.99504231e-07 1.19527885e-08 6.99604231e-07 1.19527883e-08 6.99704231e-07 1.19527885e-08 6.99804231e-07 1.19527883e-08
+ 6.99904231e-07 1.19527885e-08 7e-07 1.19527882e-08 7.0001e-07 1.45267506e-08 7.0003e-07 1.23970145e-09 7.0007e-07 2.76375265e-08 7.0015e-07 -4.37848938e-09 7.0025e-07 2.82049112e-08 7.0035e-07 -3.17728036e-09
+ 7.0045e-07 2.52046196e-08 7.0055e-07 2.60783975e-09 7.0065e-07 -4.0648491e-08 7.0075e-07 3.06912282e-06 7.0085e-07 9.51416557e-05 7.00931988e-07 -0.0447690188 7.01e-07 1.97565125 7.01008484e-07 3.09900368
+ 7.01025451e-07 4.14251596 7.01059385e-07 4.88272691 7.01090588e-07 4.97988863 7.01143428e-07 5.00280497 7.011991e-07 4.99920014 7.012991e-07 5.00046356 7.013991e-07 4.99971393 7.014991e-07 5.00018225
+ 7.01578678e-07 4.99989094 7.01663998e-07 5.00006899 7.01763998e-07 4.99995201 7.01858547e-07 5.00003258 7.01958547e-07 4.99997704 7.02058547e-07 5.00001602 7.02158547e-07 4.99998864 7.02258547e-07 5.00000791
+ 7.02358547e-07 4.99999437 7.02458547e-07 5.00000389 7.02558547e-07 4.99999721 7.02658547e-07 5.0000019 7.02758547e-07 4.99999862 7.02858547e-07 5.00000091 7.02958547e-07 4.99999932 7.03058547e-07 5.00000042
+ 7.03158547e-07 4.99999966 7.03258547e-07 5.00000018 7.03358547e-07 4.99999983 7.03458547e-07 5.00000007 7.03558547e-07 4.99999991 7.03658547e-07 5.00000001 7.03758547e-07 4.99999995 7.03858547e-07 4.99999999
+ 7.03958547e-07 4.99999996 7.04058547e-07 4.99999998 7.04158547e-07 4.99999997 7.04258547e-07 4.99999997 7.04358547e-07 4.99999997 7.04458547e-07 4.99999997 7.04558547e-07 4.99999997 7.04658547e-07 4.99999997
+ 7.04758547e-07 4.99999997 7.04858547e-07 4.99999997 7.04958547e-07 4.99999997 7.05058547e-07 4.99999997 7.05158547e-07 4.99999997 7.05258547e-07 4.99999997 7.05358547e-07 4.99999997 7.05458547e-07 4.99999997
+ 7.05558547e-07 4.99999997 7.05658547e-07 4.99999997 7.05758547e-07 4.99999997 7.05858547e-07 4.99999997 7.05958547e-07 4.99999997 7.06058547e-07 4.99999997 7.06158547e-07 4.99999997 7.06258547e-07 4.99999997
+ 7.06358547e-07 4.99999997 7.06458547e-07 4.99999997 7.06558547e-07 4.99999997 7.06658547e-07 4.99999997 7.06758547e-07 4.99999997 7.06858547e-07 4.99999997 7.06958547e-07 4.99999997 7.07058547e-07 4.99999997
+ 7.07158547e-07 4.99999997 7.07258547e-07 4.99999997 7.07358547e-07 4.99999997 7.07458547e-07 4.99999997 7.07558547e-07 4.99999997 7.07658547e-07 4.99999997 7.07758547e-07 4.99999997 7.07858547e-07 4.99999997
+ 7.07958547e-07 4.99999997 7.08058547e-07 4.99999997 7.08158547e-07 4.99999997 7.08258547e-07 4.99999997 7.08358547e-07 4.99999997 7.08458547e-07 4.99999997 7.08558547e-07 4.99999997 7.08658547e-07 4.99999997
+ 7.08758547e-07 4.99999997 7.08858547e-07 4.99999997 7.08958547e-07 4.99999997 7.09058547e-07 4.99999997 7.09158547e-07 4.99999997 7.09258547e-07 4.99999997 7.09358547e-07 4.99999997 7.09458547e-07 4.99999997
+ 7.09558547e-07 4.99999997 7.09658547e-07 4.99999997 7.09758547e-07 4.99999997 7.09858547e-07 4.99999997 7.09958547e-07 4.99999997 7.10058547e-07 4.99999997 7.10158547e-07 4.99999997 7.10258547e-07 4.99999997
+ 7.10358547e-07 4.99999997 7.10458547e-07 4.99999997 7.10558547e-07 4.99999997 7.10658547e-07 4.99999997 7.10758547e-07 4.99999997 7.10858547e-07 4.99999997 7.10958547e-07 4.99999997 7.11058547e-07 4.99999997
+ 7.11158547e-07 4.99999997 7.11258547e-07 4.99999997 7.11358547e-07 4.99999997 7.11458547e-07 4.99999997 7.11558547e-07 4.99999997 7.11658547e-07 4.99999997 7.11758547e-07 4.99999997 7.11858547e-07 4.99999997
+ 7.11958547e-07 4.99999997 7.12058547e-07 4.99999997 7.12158547e-07 4.99999997 7.12258547e-07 4.99999997 7.12358547e-07 4.99999997 7.12458547e-07 4.99999997 7.12558547e-07 4.99999997 7.12658547e-07 4.99999997
+ 7.12758547e-07 4.99999997 7.12858547e-07 4.99999997 7.12958547e-07 4.99999997 7.13058547e-07 4.99999997 7.13158547e-07 4.99999997 7.13258547e-07 4.99999997 7.13358547e-07 4.99999997 7.13458547e-07 4.99999997
+ 7.13558547e-07 4.99999997 7.13658547e-07 4.99999997 7.13758547e-07 4.99999997 7.13858547e-07 4.99999997 7.13958547e-07 4.99999997 7.14058547e-07 4.99999997 7.14158547e-07 4.99999997 7.14258547e-07 4.99999997
+ 7.14358547e-07 4.99999997 7.14458547e-07 4.99999997 7.14558547e-07 4.99999997 7.14658547e-07 4.99999997 7.14758547e-07 4.99999997 7.14858547e-07 4.99999997 7.14958547e-07 4.99999997 7.15058547e-07 4.99999997
+ 7.15158547e-07 4.99999997 7.15258547e-07 4.99999997 7.15358547e-07 4.99999997 7.15458547e-07 4.99999997 7.15558547e-07 4.99999997 7.15658547e-07 4.99999997 7.15758547e-07 4.99999997 7.15858547e-07 4.99999997
+ 7.15958547e-07 4.99999997 7.16058547e-07 4.99999997 7.16158547e-07 4.99999997 7.16258547e-07 4.99999997 7.16358547e-07 4.99999997 7.16458547e-07 4.99999997 7.16558547e-07 4.99999997 7.16658547e-07 4.99999997
+ 7.16758547e-07 4.99999997 7.16858547e-07 4.99999997 7.16958547e-07 4.99999997 7.17058547e-07 4.99999997 7.17158547e-07 4.99999997 7.17258547e-07 4.99999997 7.17358547e-07 4.99999997 7.17458547e-07 4.99999997
+ 7.17558547e-07 4.99999997 7.17658547e-07 4.99999997 7.17758547e-07 4.99999997 7.17858547e-07 4.99999997 7.17958547e-07 4.99999997 7.18058547e-07 4.99999997 7.18158547e-07 4.99999997 7.18258547e-07 4.99999997
+ 7.18358547e-07 4.99999997 7.18458547e-07 4.99999997 7.18558547e-07 4.99999997 7.18658547e-07 4.99999997 7.18758547e-07 4.99999997 7.18858547e-07 4.99999997 7.18958547e-07 4.99999997 7.19058547e-07 4.99999997
+ 7.19158547e-07 4.99999997 7.19258547e-07 4.99999997 7.19358547e-07 4.99999997 7.19458547e-07 4.99999997 7.19558547e-07 4.99999997 7.19658547e-07 4.99999997 7.19758547e-07 4.99999997 7.19858547e-07 4.99999997
+ 7.19958547e-07 4.99999997 7.20058547e-07 4.99999997 7.20158547e-07 4.99999997 7.20258547e-07 4.99999997 7.20358547e-07 4.99999997 7.20458547e-07 4.99999997 7.20558547e-07 4.99999997 7.20658547e-07 4.99999997
+ 7.20758547e-07 4.99999997 7.20858547e-07 4.99999997 7.20958547e-07 4.99999997 7.21058547e-07 4.99999997 7.21158547e-07 4.99999997 7.21258547e-07 4.99999997 7.21358547e-07 4.99999997 7.21458547e-07 4.99999997
+ 7.21558547e-07 4.99999997 7.21658547e-07 4.99999997 7.21758547e-07 4.99999997 7.21858547e-07 4.99999997 7.21958547e-07 4.99999997 7.22058547e-07 4.99999997 7.22158547e-07 4.99999997 7.22258547e-07 4.99999997
+ 7.22358547e-07 4.99999997 7.22458547e-07 4.99999997 7.22558547e-07 4.99999997 7.22658547e-07 4.99999997 7.22758547e-07 4.99999997 7.22858547e-07 4.99999997 7.22958547e-07 4.99999997 7.23058547e-07 4.99999997
+ 7.23158547e-07 4.99999997 7.23258547e-07 4.99999997 7.23358547e-07 4.99999997 7.23458547e-07 4.99999997 7.23558547e-07 4.99999997 7.23658547e-07 4.99999997 7.23758547e-07 4.99999997 7.23858547e-07 4.99999997
+ 7.23958547e-07 4.99999997 7.24058547e-07 4.99999997 7.24158547e-07 4.99999997 7.24258547e-07 4.99999997 7.24358547e-07 4.99999997 7.24458547e-07 4.99999997 7.24558547e-07 4.99999997 7.24658547e-07 4.99999997
+ 7.24758547e-07 4.99999997 7.24858547e-07 4.99999997 7.24958547e-07 4.99999997 7.25058547e-07 4.99999997 7.25158547e-07 4.99999997 7.25258547e-07 4.99999997 7.25358547e-07 4.99999997 7.25458547e-07 4.99999997
+ 7.25558547e-07 4.99999997 7.25658547e-07 4.99999997 7.25758547e-07 4.99999997 7.25858547e-07 4.99999997 7.25958547e-07 4.99999997 7.26058547e-07 4.99999997 7.26158547e-07 4.99999997 7.26258547e-07 4.99999997
+ 7.26358547e-07 4.99999997 7.26458547e-07 4.99999997 7.26558547e-07 4.99999997 7.26658547e-07 4.99999997 7.26758547e-07 4.99999997 7.26858547e-07 4.99999997 7.26958547e-07 4.99999997 7.27058547e-07 4.99999997
+ 7.27158547e-07 4.99999997 7.27258547e-07 4.99999997 7.27358547e-07 4.99999997 7.27458547e-07 4.99999997 7.27558547e-07 4.99999997 7.27658547e-07 4.99999997 7.27758547e-07 4.99999997 7.27858547e-07 4.99999997
+ 7.27958547e-07 4.99999997 7.28058547e-07 4.99999997 7.28158547e-07 4.99999997 7.28258547e-07 4.99999997 7.28358547e-07 4.99999997 7.28458547e-07 4.99999997 7.28558547e-07 4.99999997 7.28658547e-07 4.99999997
+ 7.28758547e-07 4.99999997 7.28858547e-07 4.99999997 7.28958547e-07 4.99999997 7.29058547e-07 4.99999997 7.29158547e-07 4.99999997 7.29258547e-07 4.99999997 7.29358547e-07 4.99999997 7.29458547e-07 4.99999997
+ 7.29558547e-07 4.99999997 7.29658547e-07 4.99999997 7.29758547e-07 4.99999997 7.29858547e-07 4.99999997 7.29958547e-07 4.99999997 7.30058547e-07 4.99999997 7.30158547e-07 4.99999997 7.30258547e-07 4.99999997
+ 7.30358547e-07 4.99999997 7.30458547e-07 4.99999997 7.30558547e-07 4.99999997 7.30658547e-07 4.99999997 7.30758547e-07 4.99999997 7.30858547e-07 4.99999997 7.30958547e-07 4.99999997 7.31058547e-07 4.99999997
+ 7.31158547e-07 4.99999997 7.31258547e-07 4.99999997 7.31358547e-07 4.99999997 7.31458547e-07 4.99999997 7.31558547e-07 4.99999997 7.31658547e-07 4.99999997 7.31758547e-07 4.99999997 7.31858547e-07 4.99999997
+ 7.31958547e-07 4.99999997 7.32058547e-07 4.99999997 7.32158547e-07 4.99999997 7.32258547e-07 4.99999997 7.32358547e-07 4.99999997 7.32458547e-07 4.99999997 7.32558547e-07 4.99999997 7.32658547e-07 4.99999997
+ 7.32758547e-07 4.99999997 7.32858547e-07 4.99999997 7.32958547e-07 4.99999997 7.33058547e-07 4.99999997 7.33158547e-07 4.99999997 7.33258547e-07 4.99999997 7.33358547e-07 4.99999997 7.33458547e-07 4.99999997
+ 7.33558547e-07 4.99999997 7.33658547e-07 4.99999997 7.33758547e-07 4.99999997 7.33858547e-07 4.99999997 7.33958547e-07 4.99999997 7.34058547e-07 4.99999997 7.34158547e-07 4.99999997 7.34258547e-07 4.99999997
+ 7.34358547e-07 4.99999997 7.34458547e-07 4.99999997 7.34558547e-07 4.99999997 7.34658547e-07 4.99999997 7.34758547e-07 4.99999997 7.34858547e-07 4.99999997 7.34958547e-07 4.99999997 7.35058547e-07 4.99999997
+ 7.35158547e-07 4.99999997 7.35258547e-07 4.99999997 7.35358547e-07 4.99999997 7.35458547e-07 4.99999997 7.35558547e-07 4.99999997 7.35658547e-07 4.99999997 7.35758547e-07 4.99999997 7.35858547e-07 4.99999997
+ 7.35958547e-07 4.99999997 7.36058547e-07 4.99999997 7.36158547e-07 4.99999997 7.36258547e-07 4.99999997 7.36358547e-07 4.99999997 7.36458547e-07 4.99999997 7.36558547e-07 4.99999997 7.36658547e-07 4.99999997
+ 7.36758547e-07 4.99999997 7.36858547e-07 4.99999997 7.36958547e-07 4.99999997 7.37058547e-07 4.99999997 7.37158547e-07 4.99999997 7.37258547e-07 4.99999997 7.37358547e-07 4.99999997 7.37458547e-07 4.99999997
+ 7.37558547e-07 4.99999997 7.37658547e-07 4.99999997 7.37758547e-07 4.99999997 7.37858547e-07 4.99999997 7.37958547e-07 4.99999997 7.38058547e-07 4.99999997 7.38158547e-07 4.99999997 7.38258547e-07 4.99999997
+ 7.38358547e-07 4.99999997 7.38458547e-07 4.99999997 7.38558547e-07 4.99999997 7.38658547e-07 4.99999997 7.38758547e-07 4.99999997 7.38858547e-07 4.99999997 7.38958547e-07 4.99999997 7.39058547e-07 4.99999997
+ 7.39158547e-07 4.99999997 7.39258547e-07 4.99999997 7.39358547e-07 4.99999997 7.39458547e-07 4.99999997 7.39558547e-07 4.99999997 7.39658547e-07 4.99999997 7.39758547e-07 4.99999997 7.39858547e-07 4.99999997
+ 7.39958547e-07 4.99999997 7.40058547e-07 4.99999997 7.40158547e-07 4.99999997 7.40258547e-07 4.99999997 7.40358547e-07 4.99999997 7.40458547e-07 4.99999997 7.40558547e-07 4.99999997 7.40658547e-07 4.99999997
+ 7.40758547e-07 4.99999997 7.40858547e-07 4.99999997 7.40958547e-07 4.99999997 7.41058547e-07 4.99999997 7.41158547e-07 4.99999997 7.41258547e-07 4.99999997 7.41358547e-07 4.99999997 7.41458547e-07 4.99999997
+ 7.41558547e-07 4.99999997 7.41658547e-07 4.99999997 7.41758547e-07 4.99999997 7.41858547e-07 4.99999997 7.41958547e-07 4.99999997 7.42058547e-07 4.99999997 7.42158547e-07 4.99999997 7.42258547e-07 4.99999997
+ 7.42358547e-07 4.99999997 7.42458547e-07 4.99999997 7.42558547e-07 4.99999997 7.42658547e-07 4.99999997 7.42758547e-07 4.99999997 7.42858547e-07 4.99999997 7.42958547e-07 4.99999997 7.43058547e-07 4.99999997
+ 7.43158547e-07 4.99999997 7.43258547e-07 4.99999997 7.43358547e-07 4.99999997 7.43458547e-07 4.99999997 7.43558547e-07 4.99999997 7.43658547e-07 4.99999997 7.43758547e-07 4.99999997 7.43858547e-07 4.99999997
+ 7.43958547e-07 4.99999997 7.44058547e-07 4.99999997 7.44158547e-07 4.99999997 7.44258547e-07 4.99999997 7.44358547e-07 4.99999997 7.44458547e-07 4.99999997 7.44558547e-07 4.99999997 7.44658547e-07 4.99999997
+ 7.44758547e-07 4.99999997 7.44858547e-07 4.99999997 7.44958547e-07 4.99999997 7.45058547e-07 4.99999997 7.45158547e-07 4.99999997 7.45258547e-07 4.99999997 7.45358547e-07 4.99999997 7.45458547e-07 4.99999997
+ 7.45558547e-07 4.99999997 7.45658547e-07 4.99999997 7.45758547e-07 4.99999997 7.45858547e-07 4.99999997 7.45958547e-07 4.99999997 7.46058547e-07 4.99999997 7.46158547e-07 4.99999997 7.46258547e-07 4.99999997
+ 7.46358547e-07 4.99999997 7.46458547e-07 4.99999997 7.46558547e-07 4.99999997 7.46658547e-07 4.99999997 7.46758547e-07 4.99999997 7.46858547e-07 4.99999997 7.46958547e-07 4.99999997 7.47058547e-07 4.99999997
+ 7.47158547e-07 4.99999997 7.47258547e-07 4.99999997 7.47358547e-07 4.99999997 7.47458547e-07 4.99999997 7.47558547e-07 4.99999997 7.47658547e-07 4.99999997 7.47758547e-07 4.99999997 7.47858547e-07 4.99999997
+ 7.47958547e-07 4.99999997 7.48058547e-07 4.99999997 7.48158547e-07 4.99999997 7.48258547e-07 4.99999997 7.48358547e-07 4.99999997 7.48458547e-07 4.99999997 7.48558547e-07 4.99999997 7.48658547e-07 4.99999997
+ 7.48758547e-07 4.99999997 7.48858547e-07 4.99999997 7.48958547e-07 4.99999997 7.49058547e-07 4.99999997 7.49158547e-07 4.99999997 7.49258547e-07 4.99999997 7.49358547e-07 4.99999997 7.49458547e-07 4.99999997
+ 7.49558547e-07 4.99999997 7.49658547e-07 4.99999997 7.49758547e-07 4.99999997 7.49858547e-07 4.99999997 7.49958547e-07 4.99999997 7.50058547e-07 4.99999997 7.50158547e-07 4.99999997 7.50258547e-07 4.99999997
+ 7.50358547e-07 4.99999997 7.50458547e-07 4.99999997 7.50558547e-07 4.99999997 7.50658547e-07 4.99999997 7.50758547e-07 4.99999997 7.50858547e-07 4.99999997 7.50958547e-07 4.99999997 7.51e-07 4.99999997
+ 7.5101e-07 4.99999997 7.5103e-07 4.99999998 7.5107e-07 4.99999996 7.5115e-07 4.99999998 7.5125e-07 4.99999997 7.5135e-07 4.99999997 7.5145e-07 4.99999998 7.5155e-07 4.99999996
+ 7.5165e-07 4.99999998 7.5175e-07 4.99999996 7.5185e-07 4.99999999 7.51930828e-07 5.00006471 7.52e-07 4.99916173 7.52008608e-07 4.99761842 7.52025825e-07 4.99312391 7.52060258e-07 5.01021642
+ 7.52106188e-07 5.09915302 7.52150118e-07 4.2138351 7.5219811e-07 0.290132927 7.522555e-07 -0.055559802 7.52312176e-07 0.0719919946 7.52404431e-07 -0.0580528341 7.52490759e-07 0.0521271683 7.52590759e-07 -0.0468986726
+ 7.52690759e-07 0.0429726694 7.52790759e-07 -0.0387916891 7.52890759e-07 0.0355067968 7.52990759e-07 -0.0321238152 7.53090759e-07 0.0293826519 7.53190759e-07 -0.0266208089 7.53290759e-07 0.0243463628 7.53390759e-07 -0.0220869282
+ 7.53490759e-07 0.0201946558 7.53590759e-07 -0.018340188 7.53690759e-07 0.0167656294 7.53790759e-07 -0.0152394344 7.53890759e-07 0.0139289603 7.53990759e-07 -0.0126701333 7.54090759e-07 0.0115791999 7.54190759e-07 -0.0105389933
+ 7.54290759e-07 0.00963062169 7.54390759e-07 -0.00876976083 7.54490759e-07 0.00801325014 7.54590759e-07 -0.00729991652 7.54690759e-07 0.00666976939 7.54790759e-07 -0.00607806441 7.54890759e-07 0.00555309574 7.54990759e-07 -0.00506185631
+ 7.55090759e-07 0.00462445582 7.55190759e-07 -0.00421633125 7.55290759e-07 0.00385185386 7.55390759e-07 -0.00351257961 7.55490759e-07 0.00320884134 7.55590759e-07 -0.00292666284 7.55690759e-07 0.00267352374 7.55790759e-07 -0.00243873589
+ 7.55890759e-07 0.00222775459 7.55990759e-07 -0.00203233144 7.56090759e-07 0.00185647883 7.56190759e-07 -0.00169377401 7.56290759e-07 0.00154719576 7.56390759e-07 -0.00141169917 7.56490759e-07 0.00128951848 7.56590759e-07 -0.00117744179
+ 7.56690759e-07 0.00107519826 7.56790759e-07 -0.000980224982 7.56890759e-07 0.000896201859 7.56990759e-07 -0.000816256475 7.57090759e-07 0.000747091622 7.57190759e-07 -0.000679905625 7.57290759e-07 0.000622853518 7.57390759e-07 -0.000568158092
+ 7.57490759e-07 0.000518950145 7.57590759e-07 -0.000473602727 7.57690759e-07 0.000432609181 7.57790759e-07 -0.000394813042 7.57890759e-07 0.000360641794 7.57990759e-07 -0.00032913503 7.58090759e-07 0.000300650957 7.58190759e-07 -0.000274385188
+ 7.58290759e-07 0.000250642317 7.58390759e-07 -0.000227597045 7.58490759e-07 0.000209143757 7.58590759e-07 -0.000189777838 7.58690759e-07 0.000174428486 7.58790759e-07 -0.000158243287 7.58890759e-07 0.000146480534 7.58990759e-07 -0.000131798715
+ 7.59090759e-07 0.000122072762 7.59190759e-07 -0.000109833166 7.59290759e-07 0.000101741072 7.59390759e-07 -9.15328229e-05 7.59490759e-07 8.4798664e-05 7.59590759e-07 -7.62841394e-05 7.59690759e-07 7.06796878e-05 7.59790759e-07 -6.3577359e-05
+ 7.59890759e-07 5.89130619e-05 7.59990759e-07 -5.29881514e-05 7.60090759e-07 4.91064763e-05 7.60190759e-07 -4.41632069e-05 7.60290759e-07 4.09331671e-05 7.60390759e-07 -3.68082931e-05 7.60490759e-07 3.41209287e-05 7.60590759e-07 -3.06783363e-05
+ 7.60690759e-07 2.84429787e-05 7.60790759e-07 -2.55691818e-05 7.60890759e-07 2.37103609e-05 7.60990759e-07 -2.13107424e-05 7.61090759e-07 1.97656238e-05 7.61190759e-07 -1.77613005e-05 7.61290759e-07 1.64775595e-05 7.61390759e-07 -1.48027673e-05
+ 7.61490759e-07 1.37368234e-05 7.61590759e-07 -1.23367368e-05 7.61690759e-07 1.14522874e-05 7.61790759e-07 -1.02812005e-05 7.61890759e-07 9.54800221e-06 7.61990759e-07 -8.56781254e-06 7.62090759e-07 7.96066694e-06 7.62190759e-07 -7.13961088e-06
+ 7.62290759e-07 6.63752161e-06 7.62390759e-07 -5.94912011e-06 7.62490759e-07 5.5345908e-06 7.62590759e-07 -4.95677035e-06 7.62690759e-07 4.61522039e-06 7.62790759e-07 -4.1295802e-06 7.62890759e-07 3.84885826e-06 7.62990759e-07 -3.44005922e-06
+ 7.63090759e-07 3.21003811e-06 7.63190759e-07 -2.86529346e-06 7.63290759e-07 2.67753269e-06 7.63390759e-07 -2.38618332e-06 7.63490759e-07 2.23364797e-06 7.63590759e-07 -1.98680848e-06 7.63690759e-07 1.86363501e-06 7.63790759e-07 -1.65389859e-06
+ 7.63890759e-07 1.55519979e-06 7.63990759e-07 -1.37639223e-06 7.64090759e-07 1.29809458e-06 7.64190759e-07 -1.14506907e-06 7.64290759e-07 1.08377708e-06 7.64390759e-07 -9.52243233e-07 7.64490759e-07 9.05126584e-07 7.64590759e-07 -7.91507923e-07
+ 7.64690759e-07 7.56207395e-07 7.64790759e-07 -6.57522578e-07 7.64890759e-07 6.32071612e-07 7.64990759e-07 -5.4583533e-07 7.65090759e-07 5.28594424e-07 7.65190759e-07 -4.52734886e-07 7.65290759e-07 4.42337866e-07 7.65390759e-07 -3.7512853e-07
+ 7.65490759e-07 3.70436518e-07 7.65590759e-07 -3.10437819e-07 7.65690759e-07 3.10501328e-07 7.65790759e-07 -2.56513247e-07 7.65890759e-07 2.60540816e-07 7.65990759e-07 -2.11564427e-07 7.66090759e-07 2.18897721e-07 7.66190759e-07 -1.74107636e-07
+ 7.66290759e-07 1.84205259e-07 7.66390759e-07 -1.42903498e-07 7.66490759e-07 1.55303991e-07 7.66590759e-07 -1.16908189e-07 7.66690759e-07 1.31227074e-07 7.66790759e-07 -9.52521048e-08 7.66890759e-07 1.11169114e-07 7.66990759e-07 -7.72108561e-08
+ 7.67090759e-07 9.44592506e-08 7.67190759e-07 -6.21811991e-08 7.67290759e-07 8.05388985e-08 7.67390759e-07 -4.96223675e-08 7.67490759e-07 6.89035346e-08 7.67590759e-07 -3.91967475e-08 7.67690759e-07 5.925146e-08 7.67790759e-07 -3.05155715e-08
+ 7.67890759e-07 5.12112145e-08 7.67990759e-07 -2.32838321e-08 7.68090759e-07 4.45134133e-08 7.68190759e-07 -1.72595827e-08 7.68290759e-07 3.89337721e-08 7.68390759e-07 -1.22406801e-08 7.68490759e-07 3.42853598e-08 7.68590759e-07 -8.05990238e-09
+ 7.68690759e-07 3.04134398e-08 7.68790759e-07 -4.57750143e-09 7.68890759e-07 2.71882931e-08 7.68990759e-07 -1.6768002e-09 7.69090759e-07 2.45018676e-08 7.69190759e-07 7.39380002e-10 7.69290759e-07 2.22738645e-08 7.69390759e-07 2.74369907e-09
+ 7.69490759e-07 2.04438307e-08 7.69590759e-07 4.39085443e-09 7.69690759e-07 1.89397882e-08 7.69790759e-07 5.74463149e-09 7.69890759e-07 1.77036111e-08 7.69990759e-07 6.85732449e-09 7.70090759e-07 1.66875591e-08 7.70190759e-07 7.77189338e-09
+ 7.70290759e-07 1.58524128e-08 7.70390759e-07 8.52363424e-09 7.70490759e-07 1.50671434e-08 7.70590759e-07 9.1277538e-09 7.70690759e-07 1.45150394e-08 7.70790759e-07 9.62891197e-09 7.70890759e-07 1.40604611e-08 7.70990759e-07 1.00412061e-08
+ 7.71090759e-07 1.36865218e-08 7.71190759e-07 1.0380358e-08 7.71290759e-07 1.33789217e-08 7.71390759e-07 1.06593411e-08 7.71490759e-07 1.31258937e-08 7.71590759e-07 1.08888288e-08 7.71690759e-07 1.29177566e-08 7.71790759e-07 1.10776014e-08
+ 7.71890759e-07 1.27465466e-08 7.71990759e-07 1.12328827e-08 7.72090759e-07 1.26057123e-08 7.72190759e-07 1.13606136e-08 7.72290759e-07 1.24898659e-08 7.72390759e-07 1.14656821e-08 7.72490759e-07 1.23945729e-08 7.72590759e-07 1.15521088e-08
+ 7.72690759e-07 1.23161874e-08 7.72790759e-07 1.1623201e-08 7.72890759e-07 1.22517097e-08 7.72990759e-07 1.168168e-08 7.73090759e-07 1.21986718e-08 7.73190759e-07 1.17297829e-08 7.73290759e-07 1.21550446e-08 7.73390759e-07 1.1769351e-08
+ 7.73490759e-07 1.2119158e-08 7.73590759e-07 1.18018983e-08 7.73690759e-07 1.20896388e-08 7.73790759e-07 1.18286712e-08 7.73890759e-07 1.2065357e-08 7.73990759e-07 1.18506934e-08 7.74090759e-07 1.20453836e-08 7.74190759e-07 1.18688085e-08
+ 7.74290759e-07 1.20289542e-08 7.74390759e-07 1.18837093e-08 7.74490759e-07 1.20154397e-08 7.74590759e-07 1.18959663e-08 7.74690759e-07 1.20043232e-08 7.74790759e-07 1.19060486e-08 7.74890759e-07 1.19951791e-08 7.74990759e-07 1.19143419e-08
+ 7.75090759e-07 1.19876572e-08 7.75190759e-07 1.19211634e-08 7.75290759e-07 1.19814704e-08 7.75390759e-07 1.19267747e-08 7.75490759e-07 1.19763814e-08 7.75590759e-07 1.19313903e-08 7.75690759e-07 1.19721951e-08 7.75790759e-07 1.19351871e-08
+ 7.75890759e-07 1.19687517e-08 7.75990759e-07 1.19383102e-08 7.76090759e-07 1.19659193e-08 7.76190759e-07 1.19408791e-08 7.76290759e-07 1.19635895e-08 7.76390759e-07 1.19429921e-08 7.76490759e-07 1.1961673e-08 7.76590759e-07 1.19447306e-08
+ 7.76690759e-07 1.19600964e-08 7.76790759e-07 1.19461605e-08 7.76890759e-07 1.19587996e-08 7.76990759e-07 1.19473365e-08 7.77090759e-07 1.19577328e-08 7.77190759e-07 1.19483038e-08 7.77290759e-07 1.19568556e-08 7.77390759e-07 1.19490997e-08
+ 7.77490759e-07 1.19561337e-08 7.77590759e-07 1.19497542e-08 7.77690759e-07 1.19555399e-08 7.77790759e-07 1.19502925e-08 7.77890759e-07 1.19550519e-08 7.77990759e-07 1.19507354e-08 7.78090759e-07 1.19546501e-08 7.78190759e-07 1.19510996e-08
+ 7.78290759e-07 1.195432e-08 7.78390759e-07 1.19513991e-08 7.78490759e-07 1.19540482e-08 7.78590759e-07 1.19516455e-08 7.78690759e-07 1.19538247e-08 7.78790759e-07 1.19518482e-08 7.78890759e-07 1.19536407e-08 7.78990759e-07 1.19520152e-08
+ 7.79090759e-07 1.19534895e-08 7.79190759e-07 1.19521527e-08 7.79290759e-07 1.19533653e-08 7.79390759e-07 1.19522651e-08 7.79490759e-07 1.19532625e-08 7.79590759e-07 1.1952358e-08 7.79690759e-07 1.19531783e-08 7.79790759e-07 1.19524344e-08
+ 7.79890759e-07 1.19531093e-08 7.79990759e-07 1.19524974e-08 7.80090759e-07 1.19530524e-08 7.80190759e-07 1.19525491e-08 7.80290759e-07 1.19530054e-08 7.80390759e-07 1.19525914e-08 7.80490759e-07 1.1952967e-08 7.80590759e-07 1.19526266e-08
+ 7.80690759e-07 1.19529351e-08 7.80790759e-07 1.19526554e-08 7.80890759e-07 1.1952909e-08 7.80990759e-07 1.19526787e-08 7.81090759e-07 1.19528876e-08 7.81190759e-07 1.19526981e-08 7.81290759e-07 1.195287e-08 7.81390759e-07 1.19527143e-08
+ 7.81490759e-07 1.19528555e-08 7.81590759e-07 1.19527272e-08 7.81690759e-07 1.19528438e-08 7.81790759e-07 1.19527383e-08 7.81890759e-07 1.19528339e-08 7.81990759e-07 1.19527472e-08 7.82090759e-07 1.19528258e-08 7.82190759e-07 1.19527544e-08
+ 7.82290759e-07 1.19528192e-08 7.82390759e-07 1.19527604e-08 7.82490759e-07 1.19528135e-08 7.82590759e-07 1.19527654e-08 7.82690759e-07 1.19528093e-08 7.82790759e-07 1.19527694e-08 7.82890759e-07 1.19528054e-08 7.82990759e-07 1.19527727e-08
+ 7.83090759e-07 1.19528023e-08 7.83190759e-07 1.19527756e-08 7.83290759e-07 1.19527999e-08 7.83390759e-07 1.1952778e-08 7.83490759e-07 1.19527975e-08 7.83590759e-07 1.19527798e-08 7.83690759e-07 1.19527961e-08 7.83790759e-07 1.19527814e-08
+ 7.83890759e-07 1.19527945e-08 7.83990759e-07 1.19527827e-08 7.84090759e-07 1.19527936e-08 7.84190759e-07 1.19527836e-08 7.84290759e-07 1.19527927e-08 7.84390759e-07 1.19527843e-08 7.84490759e-07 1.19527919e-08 7.84590759e-07 1.1952785e-08
+ 7.84690759e-07 1.19527911e-08 7.84790759e-07 1.19527855e-08 7.84890759e-07 1.19527909e-08 7.84990759e-07 1.19527858e-08 7.85090759e-07 1.19527904e-08 7.85190759e-07 1.19527864e-08 7.85290759e-07 1.195279e-08 7.85390759e-07 1.19527868e-08
+ 7.85490759e-07 1.19527897e-08 7.85590759e-07 1.19527869e-08 7.85690759e-07 1.19527898e-08 7.85790759e-07 1.1952787e-08 7.85890759e-07 1.19527893e-08 7.85990759e-07 1.19527872e-08 7.86090759e-07 1.19527894e-08 7.86190759e-07 1.19527874e-08
+ 7.86290759e-07 1.19527892e-08 7.86390759e-07 1.19527876e-08 7.86490759e-07 1.1952789e-08 7.86590759e-07 1.19527878e-08 7.86690759e-07 1.19527891e-08 7.86790759e-07 1.19527876e-08 7.86890759e-07 1.19527887e-08 7.86990759e-07 1.19527878e-08
+ 7.87090759e-07 1.19527888e-08 7.87190759e-07 1.1952788e-08 7.87290759e-07 1.19527888e-08 7.87390759e-07 1.19527881e-08 7.87490759e-07 1.19527887e-08 7.87590759e-07 1.19527881e-08 7.87690759e-07 1.19527886e-08 7.87790759e-07 1.19527883e-08
+ 7.87890759e-07 1.19527886e-08 7.87990759e-07 1.19527881e-08 7.88090759e-07 1.19527886e-08 7.88190759e-07 1.19527882e-08 7.88290759e-07 1.19527885e-08 7.88390759e-07 1.19527882e-08 7.88490759e-07 1.19527885e-08 7.88590759e-07 1.19527882e-08
+ 7.88690759e-07 1.19527885e-08 7.88790759e-07 1.19527882e-08 7.88890759e-07 1.19527885e-08 7.88990759e-07 1.19527882e-08 7.89090759e-07 1.19527885e-08 7.89190759e-07 1.19527882e-08 7.89290759e-07 1.19527885e-08 7.89390759e-07 1.19527882e-08
+ 7.89490759e-07 1.19527885e-08 7.89590759e-07 1.19527882e-08 7.89690759e-07 1.19527885e-08 7.89790759e-07 1.19527882e-08 7.89890759e-07 1.19527885e-08 7.89990759e-07 1.19527882e-08 7.90090759e-07 1.19527885e-08 7.90190759e-07 1.19527882e-08
+ 7.90290759e-07 1.19527885e-08 7.90390759e-07 1.19527882e-08 7.90490759e-07 1.19527885e-08 7.90590759e-07 1.19527882e-08 7.90690759e-07 1.19527885e-08 7.90790759e-07 1.19527882e-08 7.90890759e-07 1.19527885e-08 7.90990759e-07 1.19527882e-08
+ 7.91090759e-07 1.19527885e-08 7.91190759e-07 1.19527882e-08 7.91290759e-07 1.19527885e-08 7.91390759e-07 1.19527882e-08 7.91490759e-07 1.19527885e-08 7.91590759e-07 1.19527882e-08 7.91690759e-07 1.19527885e-08 7.91790759e-07 1.19527882e-08
+ 7.91890759e-07 1.19527885e-08 7.91990759e-07 1.19527882e-08 7.92090759e-07 1.19527885e-08 7.92190759e-07 1.19527882e-08 7.92290759e-07 1.19527885e-08 7.92390759e-07 1.19527882e-08 7.92490759e-07 1.19527885e-08 7.92590759e-07 1.19527882e-08
+ 7.92690759e-07 1.19527885e-08 7.92790759e-07 1.19527882e-08 7.92890759e-07 1.19527885e-08 7.92990759e-07 1.19527882e-08 7.93090759e-07 1.19527885e-08 7.93190759e-07 1.19527882e-08 7.93290759e-07 1.19527885e-08 7.93390759e-07 1.19527882e-08
+ 7.93490759e-07 1.19527885e-08 7.93590759e-07 1.19527882e-08 7.93690759e-07 1.19527885e-08 7.93790759e-07 1.19527882e-08 7.93890759e-07 1.19527885e-08 7.93990759e-07 1.19527882e-08 7.94090759e-07 1.19527885e-08 7.94190759e-07 1.19527882e-08
+ 7.94290759e-07 1.19527885e-08 7.94390759e-07 1.19527882e-08 7.94490759e-07 1.19527885e-08 7.94590759e-07 1.19527882e-08 7.94690759e-07 1.19527885e-08 7.94790759e-07 1.19527882e-08 7.94890759e-07 1.19527885e-08 7.94990759e-07 1.19527882e-08
+ 7.95090759e-07 1.19527885e-08 7.95190759e-07 1.19527882e-08 7.95290759e-07 1.19527885e-08 7.95390759e-07 1.19527882e-08 7.95490759e-07 1.19527885e-08 7.95590759e-07 1.19527882e-08 7.95690759e-07 1.19527885e-08 7.95790759e-07 1.19527882e-08
+ 7.95890759e-07 1.19527885e-08 7.95990759e-07 1.19527882e-08 7.96090759e-07 1.19527885e-08 7.96190759e-07 1.19527882e-08 7.96290759e-07 1.19527885e-08 7.96390759e-07 1.19527882e-08 7.96490759e-07 1.19527885e-08 7.96590759e-07 1.19527882e-08
+ 7.96690759e-07 1.19527885e-08 7.96790759e-07 1.19527882e-08 7.96890759e-07 1.19527885e-08 7.96990759e-07 1.19527882e-08 7.97090759e-07 1.19527885e-08 7.97190759e-07 1.19527882e-08 7.97290759e-07 1.19527885e-08 7.97390759e-07 1.19527882e-08
+ 7.97490759e-07 1.19527885e-08 7.97590759e-07 1.19527882e-08 7.97690759e-07 1.19527885e-08 7.97790759e-07 1.19527882e-08 7.97890759e-07 1.19527885e-08 7.97990759e-07 1.19527882e-08 7.98090759e-07 1.19527885e-08 7.98190759e-07 1.19527882e-08
+ 7.98290759e-07 1.19527885e-08 7.98390759e-07 1.19527882e-08 7.98490759e-07 1.19527885e-08 7.98590759e-07 1.19527882e-08 7.98690759e-07 1.19527885e-08 7.98790759e-07 1.19527882e-08 7.98890759e-07 1.19527885e-08 7.98990759e-07 1.19527882e-08
+ 7.99090759e-07 1.19527885e-08 7.99190759e-07 1.19527882e-08 7.99290759e-07 1.19527885e-08 7.99390759e-07 1.19527882e-08 7.99490759e-07 1.19527885e-08 7.99590759e-07 1.19527882e-08 7.99690759e-07 1.19527885e-08 7.99790759e-07 1.19527882e-08
+ 7.99890759e-07 1.19527885e-08 7.99990759e-07 1.19527882e-08 8e-07 1.19527883e-08 8.0001e-07 1.45272738e-08 8.0003e-07 1.23606558e-09 8.0007e-07 2.76445113e-08 8.0015e-07 -4.38735373e-09 8.0025e-07 2.82154724e-08
+ 8.0035e-07 -3.1892772e-09 8.0045e-07 2.52177674e-08 8.0055e-07 2.59407318e-09 8.0065e-07 -4.06359157e-08 8.0075e-07 3.06902779e-06 8.0085e-07 9.4837652e-05 8.00931913e-07 -0.0447404595 8.01e-07 1.97335451
+ 8.01008477e-07 3.09581876 8.01025432e-07 4.14108237 8.01059342e-07 4.88215046 8.01090545e-07 4.98042869 8.01143412e-07 5.00336525 8.01199108e-07 4.99901157 8.01266691e-07 5.00044073 8.01329415e-07 4.99978464
+ 8.01394829e-07 5.00011532 8.01464618e-07 4.99993177 8.01533535e-07 5.00004011 8.01610366e-07 4.99997429 8.01709241e-07 5.00001814 8.01809241e-07 4.99998689 8.01909241e-07 5.00000939 8.02009241e-07 4.99999309
+ 8.02109241e-07 5.000005 8.02209241e-07 4.99999625 8.02309241e-07 5.00000274 8.02409241e-07 4.99999789 8.02509241e-07 5.00000154 8.02609241e-07 4.99999877 8.02709241e-07 5.00000089 8.02809241e-07 4.99999926
+ 8.02909241e-07 5.00000052 8.03009241e-07 4.99999954 8.03109241e-07 5.00000031 8.03209241e-07 4.9999997 8.03309241e-07 5.00000019 8.03409241e-07 4.9999998 8.03509241e-07 5.00000011 8.03609241e-07 4.99999986
+ 8.03709241e-07 5.00000006 8.03809241e-07 4.9999999 8.03909241e-07 5.00000003 8.04009241e-07 4.99999992 8.04109241e-07 5.00000001 8.04209241e-07 4.99999994 8.04309241e-07 5.0 8.04409241e-07 4.99999995
+ 8.04509241e-07 4.99999999 8.04609241e-07 4.99999996 8.04709241e-07 4.99999999 8.04809241e-07 4.99999996 8.04909241e-07 4.99999998 8.05009241e-07 4.99999996 8.05109241e-07 4.99999998 8.05209241e-07 4.99999997
+ 8.05309241e-07 4.99999998 8.05409241e-07 4.99999997 8.05509241e-07 4.99999998 8.05609241e-07 4.99999997 8.05709241e-07 4.99999997 8.05809241e-07 4.99999997 8.05909241e-07 4.99999997 8.06009241e-07 4.99999997
+ 8.06109241e-07 4.99999997 8.06209241e-07 4.99999997 8.06309241e-07 4.99999997 8.06409241e-07 4.99999997 8.06509241e-07 4.99999997 8.06609241e-07 4.99999997 8.06709241e-07 4.99999997 8.06809241e-07 4.99999997
+ 8.06909241e-07 4.99999997 8.07009241e-07 4.99999997 8.07109241e-07 4.99999997 8.07209241e-07 4.99999997 8.07309241e-07 4.99999997 8.07409241e-07 4.99999997 8.07509241e-07 4.99999997 8.07609241e-07 4.99999997
+ 8.07709241e-07 4.99999997 8.07809241e-07 4.99999997 8.07909241e-07 4.99999997 8.08009241e-07 4.99999997 8.08109241e-07 4.99999997 8.08209241e-07 4.99999997 8.08309241e-07 4.99999997 8.08409241e-07 4.99999997
+ 8.08509241e-07 4.99999997 8.08609241e-07 4.99999997 8.08709241e-07 4.99999997 8.08809241e-07 4.99999997 8.08909241e-07 4.99999997 8.09009241e-07 4.99999997 8.09109241e-07 4.99999997 8.09209241e-07 4.99999997
+ 8.09309241e-07 4.99999997 8.09409241e-07 4.99999997 8.09509241e-07 4.99999997 8.09609241e-07 4.99999997 8.09709241e-07 4.99999997 8.09809241e-07 4.99999997 8.09909241e-07 4.99999997 8.10009241e-07 4.99999997
+ 8.10109241e-07 4.99999997 8.10209241e-07 4.99999997 8.10309241e-07 4.99999997 8.10409241e-07 4.99999997 8.10509241e-07 4.99999997 8.10609241e-07 4.99999997 8.10709241e-07 4.99999997 8.10809241e-07 4.99999997
+ 8.10909241e-07 4.99999997 8.11009241e-07 4.99999997 8.11109241e-07 4.99999997 8.11209241e-07 4.99999997 8.11309241e-07 4.99999997 8.11409241e-07 4.99999997 8.11509241e-07 4.99999997 8.11609241e-07 4.99999997
+ 8.11709241e-07 4.99999997 8.11809241e-07 4.99999997 8.11909241e-07 4.99999997 8.12009241e-07 4.99999997 8.12109241e-07 4.99999997 8.12209241e-07 4.99999997 8.12309241e-07 4.99999997 8.12409241e-07 4.99999997
+ 8.12509241e-07 4.99999997 8.12609241e-07 4.99999997 8.12709241e-07 4.99999997 8.12809241e-07 4.99999997 8.12909241e-07 4.99999997 8.13009241e-07 4.99999997 8.13109241e-07 4.99999997 8.13209241e-07 4.99999997
+ 8.13309241e-07 4.99999997 8.13409241e-07 4.99999997 8.13509241e-07 4.99999997 8.13609241e-07 4.99999997 8.13709241e-07 4.99999997 8.13809241e-07 4.99999997 8.13909241e-07 4.99999997 8.14009241e-07 4.99999997
+ 8.14109241e-07 4.99999997 8.14209241e-07 4.99999997 8.14309241e-07 4.99999997 8.14409241e-07 4.99999997 8.14509241e-07 4.99999997 8.14609241e-07 4.99999997 8.14709241e-07 4.99999997 8.14809241e-07 4.99999997
+ 8.14909241e-07 4.99999997 8.15009241e-07 4.99999997 8.15109241e-07 4.99999997 8.15209241e-07 4.99999997 8.15309241e-07 4.99999997 8.15409241e-07 4.99999997 8.15509241e-07 4.99999997 8.15609241e-07 4.99999997
+ 8.15709241e-07 4.99999997 8.15809241e-07 4.99999997 8.15909241e-07 4.99999997 8.16009241e-07 4.99999997 8.16109241e-07 4.99999997 8.16209241e-07 4.99999997 8.16309241e-07 4.99999997 8.16409241e-07 4.99999997
+ 8.16509241e-07 4.99999997 8.16609241e-07 4.99999997 8.16709241e-07 4.99999997 8.16809241e-07 4.99999997 8.16909241e-07 4.99999997 8.17009241e-07 4.99999997 8.17109241e-07 4.99999997 8.17209241e-07 4.99999997
+ 8.17309241e-07 4.99999997 8.17409241e-07 4.99999997 8.17509241e-07 4.99999997 8.17609241e-07 4.99999997 8.17709241e-07 4.99999997 8.17809241e-07 4.99999997 8.17909241e-07 4.99999997 8.18009241e-07 4.99999997
+ 8.18109241e-07 4.99999997 8.18209241e-07 4.99999997 8.18309241e-07 4.99999997 8.18409241e-07 4.99999997 8.18509241e-07 4.99999997 8.18609241e-07 4.99999997 8.18709241e-07 4.99999997 8.18809241e-07 4.99999997
+ 8.18909241e-07 4.99999997 8.19009241e-07 4.99999997 8.19109241e-07 4.99999997 8.19209241e-07 4.99999997 8.19309241e-07 4.99999997 8.19409241e-07 4.99999997 8.19509241e-07 4.99999997 8.19609241e-07 4.99999997
+ 8.19709241e-07 4.99999997 8.19809241e-07 4.99999997 8.19909241e-07 4.99999997 8.20009241e-07 4.99999997 8.20109241e-07 4.99999997 8.20209241e-07 4.99999997 8.20309241e-07 4.99999997 8.20409241e-07 4.99999997
+ 8.20509241e-07 4.99999997 8.20609241e-07 4.99999997 8.20709241e-07 4.99999997 8.20809241e-07 4.99999997 8.20909241e-07 4.99999997 8.21009241e-07 4.99999997 8.21109241e-07 4.99999997 8.21209241e-07 4.99999997
+ 8.21309241e-07 4.99999997 8.21409241e-07 4.99999997 8.21509241e-07 4.99999997 8.21609241e-07 4.99999997 8.21709241e-07 4.99999997 8.21809241e-07 4.99999997 8.21909241e-07 4.99999997 8.22009241e-07 4.99999997
+ 8.22109241e-07 4.99999997 8.22209241e-07 4.99999997 8.22309241e-07 4.99999997 8.22409241e-07 4.99999997 8.22509241e-07 4.99999997 8.22609241e-07 4.99999997 8.22709241e-07 4.99999997 8.22809241e-07 4.99999997
+ 8.22909241e-07 4.99999997 8.23009241e-07 4.99999997 8.23109241e-07 4.99999997 8.23209241e-07 4.99999997 8.23309241e-07 4.99999997 8.23409241e-07 4.99999997 8.23509241e-07 4.99999997 8.23609241e-07 4.99999997
+ 8.23709241e-07 4.99999997 8.23809241e-07 4.99999997 8.23909241e-07 4.99999997 8.24009241e-07 4.99999997 8.24109241e-07 4.99999997 8.24209241e-07 4.99999997 8.24309241e-07 4.99999997 8.24409241e-07 4.99999997
+ 8.24509241e-07 4.99999997 8.24609241e-07 4.99999997 8.24709241e-07 4.99999997 8.24809241e-07 4.99999997 8.24909241e-07 4.99999997 8.25009241e-07 4.99999997 8.25109241e-07 4.99999997 8.25209241e-07 4.99999997
+ 8.25309241e-07 4.99999997 8.25409241e-07 4.99999997 8.25509241e-07 4.99999997 8.25609241e-07 4.99999997 8.25709241e-07 4.99999997 8.25809241e-07 4.99999997 8.25909241e-07 4.99999997 8.26009241e-07 4.99999997
+ 8.26109241e-07 4.99999997 8.26209241e-07 4.99999997 8.26309241e-07 4.99999997 8.26409241e-07 4.99999997 8.26509241e-07 4.99999997 8.26609241e-07 4.99999997 8.26709241e-07 4.99999997 8.26809241e-07 4.99999997
+ 8.26909241e-07 4.99999997 8.27009241e-07 4.99999997 8.27109241e-07 4.99999997 8.27209241e-07 4.99999997 8.27309241e-07 4.99999997 8.27409241e-07 4.99999997 8.27509241e-07 4.99999997 8.27609241e-07 4.99999997
+ 8.27709241e-07 4.99999997 8.27809241e-07 4.99999997 8.27909241e-07 4.99999997 8.28009241e-07 4.99999997 8.28109241e-07 4.99999997 8.28209241e-07 4.99999997 8.28309241e-07 4.99999997 8.28409241e-07 4.99999997
+ 8.28509241e-07 4.99999997 8.28609241e-07 4.99999997 8.28709241e-07 4.99999997 8.28809241e-07 4.99999997 8.28909241e-07 4.99999997 8.29009241e-07 4.99999997 8.29109241e-07 4.99999997 8.29209241e-07 4.99999997
+ 8.29309241e-07 4.99999997 8.29409241e-07 4.99999997 8.29509241e-07 4.99999997 8.29609241e-07 4.99999997 8.29709241e-07 4.99999997 8.29809241e-07 4.99999997 8.29909241e-07 4.99999997 8.30009241e-07 4.99999997
+ 8.30109241e-07 4.99999997 8.30209241e-07 4.99999997 8.30309241e-07 4.99999997 8.30409241e-07 4.99999997 8.30509241e-07 4.99999997 8.30609241e-07 4.99999997 8.30709241e-07 4.99999997 8.30809241e-07 4.99999997
+ 8.30909241e-07 4.99999997 8.31009241e-07 4.99999997 8.31109241e-07 4.99999997 8.31209241e-07 4.99999997 8.31309241e-07 4.99999997 8.31409241e-07 4.99999997 8.31509241e-07 4.99999997 8.31609241e-07 4.99999997
+ 8.31709241e-07 4.99999997 8.31809241e-07 4.99999997 8.31909241e-07 4.99999997 8.32009241e-07 4.99999997 8.32109241e-07 4.99999997 8.32209241e-07 4.99999997 8.32309241e-07 4.99999997 8.32409241e-07 4.99999997
+ 8.32509241e-07 4.99999997 8.32609241e-07 4.99999997 8.32709241e-07 4.99999997 8.32809241e-07 4.99999997 8.32909241e-07 4.99999997 8.33009241e-07 4.99999997 8.33109241e-07 4.99999997 8.33209241e-07 4.99999997
+ 8.33309241e-07 4.99999997 8.33409241e-07 4.99999997 8.33509241e-07 4.99999997 8.33609241e-07 4.99999997 8.33709241e-07 4.99999997 8.33809241e-07 4.99999997 8.33909241e-07 4.99999997 8.34009241e-07 4.99999997
+ 8.34109241e-07 4.99999997 8.34209241e-07 4.99999997 8.34309241e-07 4.99999997 8.34409241e-07 4.99999997 8.34509241e-07 4.99999997 8.34609241e-07 4.99999997 8.34709241e-07 4.99999997 8.34809241e-07 4.99999997
+ 8.34909241e-07 4.99999997 8.35009241e-07 4.99999997 8.35109241e-07 4.99999997 8.35209241e-07 4.99999997 8.35309241e-07 4.99999997 8.35409241e-07 4.99999997 8.35509241e-07 4.99999997 8.35609241e-07 4.99999997
+ 8.35709241e-07 4.99999997 8.35809241e-07 4.99999997 8.35909241e-07 4.99999997 8.36009241e-07 4.99999997 8.36109241e-07 4.99999997 8.36209241e-07 4.99999997 8.36309241e-07 4.99999997 8.36409241e-07 4.99999997
+ 8.36509241e-07 4.99999997 8.36609241e-07 4.99999997 8.36709241e-07 4.99999997 8.36809241e-07 4.99999997 8.36909241e-07 4.99999997 8.37009241e-07 4.99999997 8.37109241e-07 4.99999997 8.37209241e-07 4.99999997
+ 8.37309241e-07 4.99999997 8.37409241e-07 4.99999997 8.37509241e-07 4.99999997 8.37609241e-07 4.99999997 8.37709241e-07 4.99999997 8.37809241e-07 4.99999997 8.37909241e-07 4.99999997 8.38009241e-07 4.99999997
+ 8.38109241e-07 4.99999997 8.38209241e-07 4.99999997 8.38309241e-07 4.99999997 8.38409241e-07 4.99999997 8.38509241e-07 4.99999997 8.38609241e-07 4.99999997 8.38709241e-07 4.99999997 8.38809241e-07 4.99999997
+ 8.38909241e-07 4.99999997 8.39009241e-07 4.99999997 8.39109241e-07 4.99999997 8.39209241e-07 4.99999997 8.39309241e-07 4.99999997 8.39409241e-07 4.99999997 8.39509241e-07 4.99999997 8.39609241e-07 4.99999997
+ 8.39709241e-07 4.99999997 8.39809241e-07 4.99999997 8.39909241e-07 4.99999997 8.40009241e-07 4.99999997 8.40109241e-07 4.99999997 8.40209241e-07 4.99999997 8.40309241e-07 4.99999997 8.40409241e-07 4.99999997
+ 8.40509241e-07 4.99999997 8.40609241e-07 4.99999997 8.40709241e-07 4.99999997 8.40809241e-07 4.99999997 8.40909241e-07 4.99999997 8.41009241e-07 4.99999997 8.41109241e-07 4.99999997 8.41209241e-07 4.99999997
+ 8.41309241e-07 4.99999997 8.41409241e-07 4.99999997 8.41509241e-07 4.99999997 8.41609241e-07 4.99999997 8.41709241e-07 4.99999997 8.41809241e-07 4.99999997 8.41909241e-07 4.99999997 8.42009241e-07 4.99999997
+ 8.42109241e-07 4.99999997 8.42209241e-07 4.99999997 8.42309241e-07 4.99999997 8.42409241e-07 4.99999997 8.42509241e-07 4.99999997 8.42609241e-07 4.99999997 8.42709241e-07 4.99999997 8.42809241e-07 4.99999997
+ 8.42909241e-07 4.99999997 8.43009241e-07 4.99999997 8.43109241e-07 4.99999997 8.43209241e-07 4.99999997 8.43309241e-07 4.99999997 8.43409241e-07 4.99999997 8.43509241e-07 4.99999997 8.43609241e-07 4.99999997
+ 8.43709241e-07 4.99999997 8.43809241e-07 4.99999997 8.43909241e-07 4.99999997 8.44009241e-07 4.99999997 8.44109241e-07 4.99999997 8.44209241e-07 4.99999997 8.44309241e-07 4.99999997 8.44409241e-07 4.99999997
+ 8.44509241e-07 4.99999997 8.44609241e-07 4.99999997 8.44709241e-07 4.99999997 8.44809241e-07 4.99999997 8.44909241e-07 4.99999997 8.45009241e-07 4.99999997 8.45109241e-07 4.99999997 8.45209241e-07 4.99999997
+ 8.45309241e-07 4.99999997 8.45409241e-07 4.99999997 8.45509241e-07 4.99999997 8.45609241e-07 4.99999997 8.45709241e-07 4.99999997 8.45809241e-07 4.99999997 8.45909241e-07 4.99999997 8.46009241e-07 4.99999997
+ 8.46109241e-07 4.99999997 8.46209241e-07 4.99999997 8.46309241e-07 4.99999997 8.46409241e-07 4.99999997 8.46509241e-07 4.99999997 8.46609241e-07 4.99999997 8.46709241e-07 4.99999997 8.46809241e-07 4.99999997
+ 8.46909241e-07 4.99999997 8.47009241e-07 4.99999997 8.47109241e-07 4.99999997 8.47209241e-07 4.99999997 8.47309241e-07 4.99999997 8.47409241e-07 4.99999997 8.47509241e-07 4.99999997 8.47609241e-07 4.99999997
+ 8.47709241e-07 4.99999997 8.47809241e-07 4.99999997 8.47909241e-07 4.99999997 8.48009241e-07 4.99999997 8.48109241e-07 4.99999997 8.48209241e-07 4.99999997 8.48309241e-07 4.99999997 8.48409241e-07 4.99999997
+ 8.48509241e-07 4.99999997 8.48609241e-07 4.99999997 8.48709241e-07 4.99999997 8.48809241e-07 4.99999997 8.48909241e-07 4.99999997 8.49009241e-07 4.99999997 8.49109241e-07 4.99999997 8.49209241e-07 4.99999997
+ 8.49309241e-07 4.99999997 8.49409241e-07 4.99999997 8.49509241e-07 4.99999997 8.49609241e-07 4.99999997 8.49709241e-07 4.99999997 8.49809241e-07 4.99999997 8.49909241e-07 4.99999997 8.50009241e-07 4.99999997
+ 8.50109241e-07 4.99999997 8.50209241e-07 4.99999997 8.50309241e-07 4.99999997 8.50409241e-07 4.99999997 8.50509241e-07 4.99999997 8.50609241e-07 4.99999997 8.50709241e-07 4.99999997 8.50809241e-07 4.99999997
+ 8.50909241e-07 4.99999997 8.51e-07 4.99999997 8.5101e-07 4.99999997 8.5103e-07 4.99999998 8.5107e-07 4.99999996 8.5115e-07 4.99999998 8.5125e-07 4.99999997 8.5135e-07 4.99999997
+ 8.5145e-07 4.99999998 8.5155e-07 4.99999996 8.5165e-07 4.99999998 8.5175e-07 4.99999996 8.5185e-07 4.99999999 8.51930828e-07 5.00006476 8.52e-07 4.99916064 8.52008608e-07 4.99761639
+ 8.52025825e-07 4.99311196 8.52060258e-07 5.01027311 8.52106181e-07 5.09906218 8.52150081e-07 4.21229454 8.52198026e-07 0.290284903 8.5225538e-07 -0.0554592023 8.52312019e-07 0.0719468597 8.52404232e-07 -0.0579815953
+ 8.52504232e-07 0.0528904133 8.52604232e-07 -0.0475729854 8.52704232e-07 0.0435757158 8.52804232e-07 -0.0393284178 8.52904232e-07 0.0359989191 8.53004232e-07 -0.0325572549 8.53104232e-07 0.0297863163 8.53204232e-07 -0.0269831353
+ 8.53304232e-07 0.024677895 8.53404232e-07 -0.0223854069 8.53504232e-07 0.0204676265 8.53604232e-07 -0.0185865295 8.53704232e-07 0.0169908361 8.53804232e-07 -0.0154430663 8.53904232e-07 0.0141150741 8.54004232e-07 -0.0128386861
+ 8.54104232e-07 0.0117332242 8.54204232e-07 -0.0106786681 8.54304232e-07 0.00975824024 8.54404232e-07 -0.00888561579 8.54504232e-07 0.00811909449 8.54604232e-07 -0.00739609091 8.54704232e-07 0.00675762723 8.54804232e-07 -0.00615795518
+ 8.54904232e-07 0.00562607399 8.55004232e-07 -0.00512825797 8.55104232e-07 0.00468510952 8.55204232e-07 -0.00427154749 8.55304232e-07 0.00390228875 8.55404232e-07 -0.00355851286 8.55504232e-07 0.00325079606 8.55604232e-07 -0.00296488651
+ 8.55704232e-07 0.002708436 8.55804232e-07 -0.0024705529 8.55904232e-07 0.00225681481 8.56004232e-07 -0.00205882186 8.56104232e-07 0.00188067375 8.56204232e-07 -0.00171583399 8.56304232e-07 0.00156734401 8.56404232e-07 -0.00143007279
+ 8.56504232e-07 0.00130629977 8.56604232e-07 -0.00119196316 8.56704232e-07 0.00108879052 8.56804232e-07 -0.000993540456 8.56904232e-07 0.000907538165 8.57004232e-07 -0.000828177003 8.57104232e-07 0.000756486787 8.57204232e-07 -0.000690355922
+ 8.57304232e-07 0.000630595752 8.57404232e-07 -0.00057548372 8.57504232e-07 0.00052566832 8.57604232e-07 -0.000479734899 8.57704232e-07 0.000438209567 8.57804232e-07 -0.000399922963 8.57904232e-07 0.000365308462 8.58004232e-07 -0.000333393279
+ 8.58104232e-07 0.000304539933 8.58204232e-07 -0.000277934025 8.58304232e-07 0.000253883483 8.58404232e-07 -0.000231702133 8.58504232e-07 0.000211655506 8.58604232e-07 -0.000193161676 8.58704232e-07 0.00017645299 8.58804232e-07 -0.000161032592
+ 8.58904232e-07 0.000147106668 8.59004232e-07 -0.000134248002 8.59104232e-07 0.000122642012 8.59204232e-07 -0.000111918653 8.59304232e-07 0.000102246759 8.59404232e-07 -9.33033251e-05 8.59504232e-07 8.52438625e-05 8.59604232e-07 -7.7784159e-05
+ 8.59704232e-07 7.10689667e-05 8.59804232e-07 -6.48461156e-05 8.59904232e-07 5.92516325e-05 8.60004232e-07 -5.40598536e-05 8.60104232e-07 4.93997006e-05 8.60204232e-07 -4.50674637e-05 8.60304232e-07 4.11862589e-05 8.60404232e-07 -3.75705791e-05
+ 8.60504232e-07 3.43387821e-05 8.60604232e-07 -3.13204668e-05 8.60704232e-07 2.86300807e-05 8.60804232e-07 -2.61097683e-05 8.60904232e-07 2.38707567e-05 8.61004232e-07 -2.17656161e-05 8.61104232e-07 1.9902916e-05 8.61204232e-07 -1.81438953e-05
+ 8.61304232e-07 1.65949268e-05 8.61404232e-07 -1.51244604e-05 8.61504232e-07 1.38370509e-05 8.61604232e-07 -1.26071484e-05 8.61704232e-07 1.15378015e-05 8.61804232e-07 -1.05084548e-05 8.61904232e-07 9.62090748e-06 8.62004232e-07 -8.75876282e-06
+ 8.62104232e-07 8.02278265e-06 8.62204232e-07 -7.30003353e-06 8.62304232e-07 6.69041563e-06 8.62404232e-07 -6.08388022e-06 8.62504232e-07 5.57961123e-06 8.62604232e-07 -5.0699631e-06 8.62704232e-07 4.65352411e-06 8.62804232e-07 -4.22465098e-06
+ 8.62904232e-07 3.88143644e-06 8.63004232e-07 -3.5199056e-06 8.63104232e-07 3.23773878e-06 8.63204232e-07 -2.93235145e-06 8.63304232e-07 2.70108056e-06 8.63404232e-07 -2.44250033e-06 8.63504232e-07 2.2536618e-06 8.63604232e-07 -2.03410491e-06
+ 8.63704232e-07 1.88064259e-06 8.63804232e-07 -1.69361974e-06 8.63904232e-07 1.56965094e-06 8.64004232e-07 -1.40079513e-06 8.64104232e-07 1.32022171e-06 8.64204232e-07 -1.16495131e-06 8.64304232e-07 1.10221054e-06 8.64404232e-07 -9.68845144e-07
+ 8.64504232e-07 9.20524804e-07 8.64604232e-07 -8.05378012e-07 8.64704232e-07 7.69073298e-07 8.64804232e-07 -6.69112945e-07 8.64904232e-07 6.42824079e-07 8.65004232e-07 -5.55523018e-07 8.65104232e-07 5.37583117e-07 8.65204232e-07 -4.60834663e-07
+ 8.65304232e-07 4.49854028e-07 8.65404232e-07 -3.81902011e-07 8.65504232e-07 3.76722692e-07 8.65604232e-07 -3.16103657e-07 8.65704232e-07 3.15760337e-07 8.65804232e-07 -2.61254025e-07 8.65904232e-07 2.64941894e-07 8.66004232e-07 -2.15531318e-07
+ 8.66104232e-07 2.22579736e-07 8.66204232e-07 -1.77426888e-07 8.66304232e-07 1.87286699e-07 8.66404232e-07 -1.45681874e-07 8.66504232e-07 1.57883812e-07 8.66604232e-07 -1.19234754e-07 8.66704232e-07 1.33387825e-07 8.66804232e-07 -9.72011649e-08
+ 8.66904232e-07 1.1297967e-07 8.67004232e-07 -7.88444124e-08 8.67104232e-07 9.59770695e-08 8.67204232e-07 -6.35509263e-08 8.67304232e-07 8.18118435e-08 8.67404232e-07 -5.07711887e-08 8.67504232e-07 6.9971415e-08 8.67604232e-07 -4.0160915e-08
+ 8.67704232e-07 6.01479455e-08 8.67804232e-07 -3.13252139e-08 8.67904232e-07 5.19642377e-08 8.68004232e-07 -2.39641146e-08 8.68104232e-07 4.51463207e-08 8.68204232e-07 -1.78315385e-08 8.68304232e-07 3.94660683e-08 8.68404232e-07 -1.27218723e-08
+ 8.68504232e-07 3.47333431e-08 8.68604232e-07 -8.46503109e-09 8.68704232e-07 3.07907579e-08 8.68804232e-07 -4.91886643e-09 8.68904232e-07 2.75063606e-08 8.69004232e-07 -1.96468886e-09 8.69104232e-07 2.47702319e-08 8.69204232e-07 4.96362257e-10
+ 8.69304232e-07 2.24973247e-08 8.69404232e-07 2.54107424e-09 8.69504232e-07 2.06302844e-08 8.69604232e-07 4.22167007e-09 8.69704232e-07 1.90955799e-08 8.69804232e-07 5.60316776e-09 8.69904232e-07 1.78339727e-08 8.70004232e-07 6.73886072e-09
+ 8.70104232e-07 1.67968122e-08 8.70204232e-07 7.67253122e-09 8.70304232e-07 1.59441262e-08 8.70404232e-07 8.44015208e-09 8.70504232e-07 1.51437649e-08 8.70604232e-07 9.05741751e-09 8.70704232e-07 1.45796341e-08 8.70804232e-07 9.56956192e-09
+ 8.70904232e-07 1.41150189e-08 8.71004232e-07 9.99102842e-09 8.71104232e-07 1.37326948e-08 8.71204232e-07 1.03378478e-08 8.71304232e-07 1.34180805e-08 8.71404232e-07 1.062325e-08 8.71504232e-07 1.31591759e-08 8.71604232e-07 1.08581193e-08
+ 8.71704232e-07 1.29461078e-08 8.71804232e-07 1.1051412e-08 8.71904232e-07 1.27707535e-08 8.72004232e-07 1.12104951e-08 8.72104232e-07 1.26264302e-08 8.72204232e-07 1.13414299e-08 8.72304232e-07 1.25076398e-08 8.72404232e-07 1.14492037e-08
+ 8.72504232e-07 1.24098594e-08 8.72604232e-07 1.15379188e-08 8.72704232e-07 1.23293674e-08 8.72804232e-07 1.16109513e-08 8.72904232e-07 1.22631016e-08 8.73004232e-07 1.16710786e-08 8.73104232e-07 1.22085435e-08 8.73204232e-07 1.17205849e-08
+ 8.73304232e-07 1.216362e-08 8.73404232e-07 1.17613505e-08 8.73504232e-07 1.21266263e-08 8.73604232e-07 1.17949223e-08 8.73704232e-07 1.20961589e-08 8.73804232e-07 1.18225738e-08 8.73904232e-07 1.20710628e-08 8.74004232e-07 1.1845351e-08
+ 8.74104232e-07 1.20503885e-08 8.74204232e-07 1.18641174e-08 8.74304232e-07 1.2033354e-08 8.74404232e-07 1.18795806e-08 8.74504232e-07 1.20193161e-08 8.74604232e-07 1.18923248e-08 8.74704232e-07 1.20077457e-08 8.74804232e-07 1.19028304e-08
+ 8.74904232e-07 1.19982068e-08 8.75004232e-07 1.19114921e-08 8.75104232e-07 1.19903411e-08 8.75204232e-07 1.19186353e-08 8.75304232e-07 1.19838534e-08 8.75404232e-07 1.19245281e-08 8.75504232e-07 1.19785009e-08 8.75604232e-07 1.19293903e-08
+ 8.75704232e-07 1.19740838e-08 8.75804232e-07 1.19334034e-08 8.75904232e-07 1.19704372e-08 8.76004232e-07 1.19367173e-08 8.76104232e-07 1.19674256e-08 8.76204232e-07 1.19394546e-08 8.76304232e-07 1.19649375e-08 8.76404232e-07 1.19417165e-08
+ 8.76504232e-07 1.19628807e-08 8.76604232e-07 1.19435865e-08 8.76704232e-07 1.19611799e-08 8.76804232e-07 1.19451337e-08 8.76904232e-07 1.19597724e-08 8.77004232e-07 1.19464139e-08 8.77104232e-07 1.19586076e-08 8.77204232e-07 1.19474744e-08
+ 8.77304232e-07 1.19576424e-08 8.77404232e-07 1.19483528e-08 8.77504232e-07 1.19568426e-08 8.77604232e-07 1.19490811e-08 8.77704232e-07 1.19561789e-08 8.77804232e-07 1.19496861e-08 8.77904232e-07 1.19556278e-08 8.78004232e-07 1.19501883e-08
+ 8.78104232e-07 1.19551703e-08 8.78204232e-07 1.19506056e-08 8.78304232e-07 1.19547895e-08 8.78404232e-07 1.19509529e-08 8.78504232e-07 1.19544726e-08 8.78604232e-07 1.19512422e-08 8.78704232e-07 1.19542082e-08 8.78804232e-07 1.19514836e-08
+ 8.78904232e-07 1.19539877e-08 8.79004232e-07 1.1951685e-08 8.79104232e-07 1.19538037e-08 8.79204232e-07 1.19518534e-08 8.79304232e-07 1.19536496e-08 8.79404232e-07 1.19519948e-08 8.79504232e-07 1.19535203e-08 8.79604232e-07 1.1952113e-08
+ 8.79704232e-07 1.19534118e-08 8.79804232e-07 1.19522123e-08 8.79904232e-07 1.19533209e-08 8.80004232e-07 1.19522957e-08 8.80104232e-07 1.19532443e-08 8.80204232e-07 1.19523663e-08 8.80304232e-07 1.1953179e-08 8.80404232e-07 1.19524258e-08
+ 8.80504232e-07 1.19531248e-08 8.80604232e-07 1.19524759e-08 8.80704232e-07 1.19530782e-08 8.80804232e-07 1.19525187e-08 8.80904232e-07 1.19530389e-08 8.81004232e-07 1.19525548e-08 8.81104232e-07 1.19530057e-08 8.81204232e-07 1.19525861e-08
+ 8.81304232e-07 1.19529769e-08 8.81404232e-07 1.19526123e-08 8.81504232e-07 1.19529525e-08 8.81604232e-07 1.19526349e-08 8.81704232e-07 1.19529316e-08 8.81804232e-07 1.19526543e-08 8.81904232e-07 1.19529136e-08 8.82004232e-07 1.19526709e-08
+ 8.82104232e-07 1.19528984e-08 8.82204232e-07 1.19526852e-08 8.82304232e-07 1.19528849e-08 8.82404232e-07 1.19526977e-08 8.82504232e-07 1.19528734e-08 8.82604232e-07 1.19527084e-08 8.82704232e-07 1.19528634e-08 8.82804232e-07 1.19527176e-08
+ 8.82904232e-07 1.19528547e-08 8.83004232e-07 1.19527259e-08 8.83104232e-07 1.19528473e-08 8.83204232e-07 1.19527328e-08 8.83304232e-07 1.19528405e-08 8.83404232e-07 1.19527392e-08 8.83504232e-07 1.19528347e-08 8.83604232e-07 1.19527446e-08
+ 8.83704232e-07 1.19528297e-08 8.83804232e-07 1.19527493e-08 8.83904232e-07 1.19528252e-08 8.84004232e-07 1.19527537e-08 8.84104232e-07 1.19528209e-08 8.84204232e-07 1.19527572e-08 8.84304232e-07 1.19528177e-08 8.84404232e-07 1.19527603e-08
+ 8.84504232e-07 1.19528145e-08 8.84604232e-07 1.19527634e-08 8.84704232e-07 1.19528118e-08 8.84804232e-07 1.19527659e-08 8.84904232e-07 1.19528095e-08 8.85004232e-07 1.19527683e-08 8.85104232e-07 1.19528072e-08 8.85204232e-07 1.19527702e-08
+ 8.85304232e-07 1.19528053e-08 8.85404232e-07 1.1952772e-08 8.85504232e-07 1.19528037e-08 8.85604232e-07 1.19527738e-08 8.85704232e-07 1.1952802e-08 8.85804232e-07 1.19527753e-08 8.85904232e-07 1.19528006e-08 8.86004232e-07 1.19527765e-08
+ 8.86104232e-07 1.19527997e-08 8.86204232e-07 1.19527775e-08 8.86304232e-07 1.19527985e-08 8.86404232e-07 1.19527786e-08 8.86504232e-07 1.19527974e-08 8.86604232e-07 1.19527795e-08 8.86704232e-07 1.19527965e-08 8.86804232e-07 1.19527808e-08
+ 8.86904232e-07 1.19527956e-08 8.87004232e-07 1.19527814e-08 8.87104232e-07 1.19527948e-08 8.87204232e-07 1.1952782e-08 8.87304232e-07 1.19527943e-08 8.87404232e-07 1.19527827e-08 8.87504232e-07 1.19527937e-08 8.87604232e-07 1.1952783e-08
+ 8.87704232e-07 1.19527933e-08 8.87804232e-07 1.19527837e-08 8.87904232e-07 1.1952793e-08 8.88004232e-07 1.19527841e-08 8.88104232e-07 1.19527925e-08 8.88204232e-07 1.19527846e-08 8.88304232e-07 1.19527922e-08 8.88404232e-07 1.19527849e-08
+ 8.88504232e-07 1.19527915e-08 8.88604232e-07 1.19527853e-08 8.88704232e-07 1.19527913e-08 8.88804232e-07 1.19527855e-08 8.88904232e-07 1.1952791e-08 8.89004232e-07 1.19527859e-08 8.89104232e-07 1.19527907e-08 8.89204232e-07 1.19527863e-08
+ 8.89304232e-07 1.19527905e-08 8.89404232e-07 1.19527863e-08 8.89504232e-07 1.19527903e-08 8.89604232e-07 1.19527866e-08 8.89704232e-07 1.19527898e-08 8.89804232e-07 1.19527869e-08 8.89904232e-07 1.19527899e-08 8.90004232e-07 1.19527869e-08
+ 8.90104232e-07 1.19527897e-08 8.90204232e-07 1.19527869e-08 8.90304232e-07 1.19527899e-08 8.90404232e-07 1.19527869e-08 8.90504232e-07 1.19527898e-08 8.90604232e-07 1.1952787e-08 8.90704232e-07 1.19527898e-08 8.90804232e-07 1.1952787e-08
+ 8.90904232e-07 1.19527898e-08 8.91004232e-07 1.1952787e-08 8.91104232e-07 1.19527894e-08 8.91204232e-07 1.19527871e-08 8.91304232e-07 1.19527895e-08 8.91404232e-07 1.19527872e-08 8.91504232e-07 1.19527896e-08 8.91604232e-07 1.19527873e-08
+ 8.91704232e-07 1.19527891e-08 8.91804232e-07 1.19527873e-08 8.91904232e-07 1.19527894e-08 8.92004232e-07 1.19527875e-08 8.92104232e-07 1.19527893e-08 8.92204232e-07 1.19527874e-08 8.92304232e-07 1.19527892e-08 8.92404232e-07 1.19527876e-08
+ 8.92504232e-07 1.1952789e-08 8.92604232e-07 1.19527877e-08 8.92704232e-07 1.19527891e-08 8.92804232e-07 1.19527876e-08 8.92904232e-07 1.19527891e-08 8.93004232e-07 1.19527877e-08 8.93104232e-07 1.1952789e-08 8.93204232e-07 1.19527878e-08
+ 8.93304232e-07 1.19527891e-08 8.93404232e-07 1.19527877e-08 8.93504232e-07 1.1952789e-08 8.93604232e-07 1.19527879e-08 8.93704232e-07 1.19527889e-08 8.93804232e-07 1.19527879e-08 8.93904232e-07 1.19527889e-08 8.94004232e-07 1.19527879e-08
+ 8.94104232e-07 1.19527888e-08 8.94204232e-07 1.1952788e-08 8.94304232e-07 1.19527889e-08 8.94404232e-07 1.19527879e-08 8.94504232e-07 1.19527889e-08 8.94604232e-07 1.1952788e-08 8.94704232e-07 1.19527888e-08 8.94804232e-07 1.1952788e-08
+ 8.94904232e-07 1.19527887e-08 8.95004232e-07 1.1952788e-08 8.95104232e-07 1.19527888e-08 8.95204232e-07 1.19527881e-08 8.95304232e-07 1.19527887e-08 8.95404232e-07 1.1952788e-08 8.95504232e-07 1.19527887e-08 8.95604232e-07 1.1952788e-08
+ 8.95704232e-07 1.19527887e-08 8.95804232e-07 1.19527881e-08 8.95904232e-07 1.19527887e-08 8.96004232e-07 1.19527881e-08 8.96104232e-07 1.19527886e-08 8.96204232e-07 1.1952788e-08 8.96304232e-07 1.19527887e-08 8.96404232e-07 1.19527881e-08
+ 8.96504232e-07 1.19527886e-08 8.96604232e-07 1.19527882e-08 8.96704232e-07 1.19527887e-08 8.96804232e-07 1.1952788e-08 8.96904232e-07 1.19527886e-08 8.97004232e-07 1.19527882e-08 8.97104232e-07 1.19527886e-08 8.97204232e-07 1.19527882e-08
+ 8.97304232e-07 1.19527886e-08 8.97404232e-07 1.19527881e-08 8.97504232e-07 1.19527886e-08 8.97604232e-07 1.19527881e-08 8.97704232e-07 1.19527886e-08 8.97804232e-07 1.19527883e-08 8.97904232e-07 1.19527884e-08 8.98004232e-07 1.19527882e-08
+ 8.98104232e-07 1.19527885e-08 8.98204232e-07 1.19527883e-08 8.98304232e-07 1.19527885e-08 8.98404232e-07 1.19527883e-08 8.98504232e-07 1.19527885e-08 8.98604232e-07 1.19527883e-08 8.98704232e-07 1.19527885e-08 8.98804232e-07 1.19527883e-08
+ 8.98904232e-07 1.19527885e-08 8.99004232e-07 1.19527883e-08 8.99104232e-07 1.19527885e-08 8.99204232e-07 1.19527883e-08 8.99304232e-07 1.19527885e-08 8.99404232e-07 1.19527883e-08 8.99504232e-07 1.19527885e-08 8.99604232e-07 1.19527883e-08
+ 8.99704232e-07 1.19527885e-08 8.99804232e-07 1.19527883e-08 8.99904232e-07 1.19527885e-08 9e-07 1.19527883e-08 9.0001e-07 1.45267509e-08 9.0003e-07 1.23970223e-09 9.0007e-07 2.7637525e-08 9.0015e-07 -4.37848716e-09
+ 9.0025e-07 2.82049084e-08 9.0035e-07 -3.17727716e-09 9.0045e-07 2.52046159e-08 9.0055e-07 2.60784397e-09 9.0065e-07 -4.06484961e-08 9.0075e-07 3.06912285e-06 9.0085e-07 9.51416721e-05 9.00932051e-07 -0.0447831027
+ 9.01e-07 1.97583273 9.01008488e-07 3.09989962 9.01025463e-07 4.14313244 9.01059414e-07 4.88304728 9.0109062e-07 4.97992695 9.0114347e-07 5.00280645 9.01199151e-07 4.99919782 9.01299151e-07 5.00046536
+ 9.01399151e-07 4.99971259 9.01499151e-07 5.00018323 9.01599151e-07 4.99987811 9.01699151e-07 5.00008217 9.01799151e-07 4.99994319 9.01893327e-07 5.00003835 9.01993327e-07 4.99997304 9.02093327e-07 5.00001879
+ 9.02193327e-07 4.99998671 9.02293327e-07 5.00000926 9.02393327e-07 4.99999342 9.02493327e-07 5.00000455 9.02593327e-07 4.99999675 9.02693327e-07 5.00000222 9.02793327e-07 4.9999984 9.02893327e-07 5.00000107
+ 9.02993327e-07 4.99999921 9.03093327e-07 5.0000005 9.03193327e-07 4.99999961 9.03293327e-07 5.00000022 9.03393327e-07 4.9999998 9.03493327e-07 5.00000008 9.03593327e-07 4.9999999 9.03693327e-07 5.00000002
+ 9.03793327e-07 4.99999994 9.03893327e-07 4.99999999 9.03993327e-07 4.99999996 9.04093327e-07 4.99999998 9.04193327e-07 4.99999997 9.04293327e-07 4.99999997 9.04393327e-07 4.99999997 9.04493327e-07 4.99999997
+ 9.04593327e-07 4.99999997 9.04693327e-07 4.99999997 9.04793327e-07 4.99999997 9.04893327e-07 4.99999997 9.04993327e-07 4.99999997 9.05093327e-07 4.99999997 9.05193327e-07 4.99999997 9.05293327e-07 4.99999997
+ 9.05393327e-07 4.99999997 9.05493327e-07 4.99999997 9.05593327e-07 4.99999997 9.05693327e-07 4.99999997 9.05793327e-07 4.99999997 9.05893327e-07 4.99999997 9.05993327e-07 4.99999997 9.06093327e-07 4.99999997
+ 9.06193327e-07 4.99999997 9.06293327e-07 4.99999997 9.06393327e-07 4.99999997 9.06493327e-07 4.99999997 9.06593327e-07 4.99999997 9.06693327e-07 4.99999997 9.06793327e-07 4.99999997 9.06893327e-07 4.99999997
+ 9.06993327e-07 4.99999997 9.07093327e-07 4.99999997 9.07193327e-07 4.99999997 9.07293327e-07 4.99999997 9.07393327e-07 4.99999997 9.07493327e-07 4.99999997 9.07593327e-07 4.99999997 9.07693327e-07 4.99999997
+ 9.07793327e-07 4.99999997 9.07893327e-07 4.99999997 9.07993327e-07 4.99999997 9.08093327e-07 4.99999997 9.08193327e-07 4.99999997 9.08293327e-07 4.99999997 9.08393327e-07 4.99999997 9.08493327e-07 4.99999997
+ 9.08593327e-07 4.99999997 9.08693327e-07 4.99999997 9.08793327e-07 4.99999997 9.08893327e-07 4.99999997 9.08993327e-07 4.99999997 9.09093327e-07 4.99999997 9.09193327e-07 4.99999997 9.09293327e-07 4.99999997
+ 9.09393327e-07 4.99999997 9.09493327e-07 4.99999997 9.09593327e-07 4.99999997 9.09693327e-07 4.99999997 9.09793327e-07 4.99999997 9.09893327e-07 4.99999997 9.09993327e-07 4.99999997 9.10093327e-07 4.99999997
+ 9.10193327e-07 4.99999997 9.10293327e-07 4.99999997 9.10393327e-07 4.99999997 9.10493327e-07 4.99999997 9.10593327e-07 4.99999997 9.10693327e-07 4.99999997 9.10793327e-07 4.99999997 9.10893327e-07 4.99999997
+ 9.10993327e-07 4.99999997 9.11093327e-07 4.99999997 9.11193327e-07 4.99999997 9.11293327e-07 4.99999997 9.11393327e-07 4.99999997 9.11493327e-07 4.99999997 9.11593327e-07 4.99999997 9.11693327e-07 4.99999997
+ 9.11793327e-07 4.99999997 9.11893327e-07 4.99999997 9.11993327e-07 4.99999997 9.12093327e-07 4.99999997 9.12193327e-07 4.99999997 9.12293327e-07 4.99999997 9.12393327e-07 4.99999997 9.12493327e-07 4.99999997
+ 9.12593327e-07 4.99999997 9.12693327e-07 4.99999997 9.12793327e-07 4.99999997 9.12893327e-07 4.99999997 9.12993327e-07 4.99999997 9.13093327e-07 4.99999997 9.13193327e-07 4.99999997 9.13293327e-07 4.99999997
+ 9.13393327e-07 4.99999997 9.13493327e-07 4.99999997 9.13593327e-07 4.99999997 9.13693327e-07 4.99999997 9.13793327e-07 4.99999997 9.13893327e-07 4.99999997 9.13993327e-07 4.99999997 9.14093327e-07 4.99999997
+ 9.14193327e-07 4.99999997 9.14293327e-07 4.99999997 9.14393327e-07 4.99999997 9.14493327e-07 4.99999997 9.14593327e-07 4.99999997 9.14693327e-07 4.99999997 9.14793327e-07 4.99999997 9.14893327e-07 4.99999997
+ 9.14993327e-07 4.99999997 9.15093327e-07 4.99999997 9.15193327e-07 4.99999997 9.15293327e-07 4.99999997 9.15393327e-07 4.99999997 9.15493327e-07 4.99999997 9.15593327e-07 4.99999997 9.15693327e-07 4.99999997
+ 9.15793327e-07 4.99999997 9.15893327e-07 4.99999997 9.15993327e-07 4.99999997 9.16093327e-07 4.99999997 9.16193327e-07 4.99999997 9.16293327e-07 4.99999997 9.16393327e-07 4.99999997 9.16493327e-07 4.99999997
+ 9.16593327e-07 4.99999997 9.16693327e-07 4.99999997 9.16793327e-07 4.99999997 9.16893327e-07 4.99999997 9.16993327e-07 4.99999997 9.17093327e-07 4.99999997 9.17193327e-07 4.99999997 9.17293327e-07 4.99999997
+ 9.17393327e-07 4.99999997 9.17493327e-07 4.99999997 9.17593327e-07 4.99999997 9.17693327e-07 4.99999997 9.17793327e-07 4.99999997 9.17893327e-07 4.99999997 9.17993327e-07 4.99999997 9.18093327e-07 4.99999997
+ 9.18193327e-07 4.99999997 9.18293327e-07 4.99999997 9.18393327e-07 4.99999997 9.18493327e-07 4.99999997 9.18593327e-07 4.99999997 9.18693327e-07 4.99999997 9.18793327e-07 4.99999997 9.18893327e-07 4.99999997
+ 9.18993327e-07 4.99999997 9.19093327e-07 4.99999997 9.19193327e-07 4.99999997 9.19293327e-07 4.99999997 9.19393327e-07 4.99999997 9.19493327e-07 4.99999997 9.19593327e-07 4.99999997 9.19693327e-07 4.99999997
+ 9.19793327e-07 4.99999997 9.19893327e-07 4.99999997 9.19993327e-07 4.99999997 9.20093327e-07 4.99999997 9.20193327e-07 4.99999997 9.20293327e-07 4.99999997 9.20393327e-07 4.99999997 9.20493327e-07 4.99999997
+ 9.20593327e-07 4.99999997 9.20693327e-07 4.99999997 9.20793327e-07 4.99999997 9.20893327e-07 4.99999997 9.20993327e-07 4.99999997 9.21093327e-07 4.99999997 9.21193327e-07 4.99999997 9.21293327e-07 4.99999997
+ 9.21393327e-07 4.99999997 9.21493327e-07 4.99999997 9.21593327e-07 4.99999997 9.21693327e-07 4.99999997 9.21793327e-07 4.99999997 9.21893327e-07 4.99999997 9.21993327e-07 4.99999997 9.22093327e-07 4.99999997
+ 9.22193327e-07 4.99999997 9.22293327e-07 4.99999997 9.22393327e-07 4.99999997 9.22493327e-07 4.99999997 9.22593327e-07 4.99999997 9.22693327e-07 4.99999997 9.22793327e-07 4.99999997 9.22893327e-07 4.99999997
+ 9.22993327e-07 4.99999997 9.23093327e-07 4.99999997 9.23193327e-07 4.99999997 9.23293327e-07 4.99999997 9.23393327e-07 4.99999997 9.23493327e-07 4.99999997 9.23593327e-07 4.99999997 9.23693327e-07 4.99999997
+ 9.23793327e-07 4.99999997 9.23893327e-07 4.99999997 9.23993327e-07 4.99999997 9.24093327e-07 4.99999997 9.24193327e-07 4.99999997 9.24293327e-07 4.99999997 9.24393327e-07 4.99999997 9.24493327e-07 4.99999997
+ 9.24593327e-07 4.99999997 9.24693327e-07 4.99999997 9.24793327e-07 4.99999997 9.24893327e-07 4.99999997 9.24993327e-07 4.99999997 9.25093327e-07 4.99999997 9.25193327e-07 4.99999997 9.25293327e-07 4.99999997
+ 9.25393327e-07 4.99999997 9.25493327e-07 4.99999997 9.25593327e-07 4.99999997 9.25693327e-07 4.99999997 9.25793327e-07 4.99999997 9.25893327e-07 4.99999997 9.25993327e-07 4.99999997 9.26093327e-07 4.99999997
+ 9.26193327e-07 4.99999997 9.26293327e-07 4.99999997 9.26393327e-07 4.99999997 9.26493327e-07 4.99999997 9.26593327e-07 4.99999997 9.26693327e-07 4.99999997 9.26793327e-07 4.99999997 9.26893327e-07 4.99999997
+ 9.26993327e-07 4.99999997 9.27093327e-07 4.99999997 9.27193327e-07 4.99999997 9.27293327e-07 4.99999997 9.27393327e-07 4.99999997 9.27493327e-07 4.99999997 9.27593327e-07 4.99999997 9.27693327e-07 4.99999997
+ 9.27793327e-07 4.99999997 9.27893327e-07 4.99999997 9.27993327e-07 4.99999997 9.28093327e-07 4.99999997 9.28193327e-07 4.99999997 9.28293327e-07 4.99999997 9.28393327e-07 4.99999997 9.28493327e-07 4.99999997
+ 9.28593327e-07 4.99999997 9.28693327e-07 4.99999997 9.28793327e-07 4.99999997 9.28893327e-07 4.99999997 9.28993327e-07 4.99999997 9.29093327e-07 4.99999997 9.29193327e-07 4.99999997 9.29293327e-07 4.99999997
+ 9.29393327e-07 4.99999997 9.29493327e-07 4.99999997 9.29593327e-07 4.99999997 9.29693327e-07 4.99999997 9.29793327e-07 4.99999997 9.29893327e-07 4.99999997 9.29993327e-07 4.99999997 9.30093327e-07 4.99999997
+ 9.30193327e-07 4.99999997 9.30293327e-07 4.99999997 9.30393327e-07 4.99999997 9.30493327e-07 4.99999997 9.30593327e-07 4.99999997 9.30693327e-07 4.99999997 9.30793327e-07 4.99999997 9.30893327e-07 4.99999997
+ 9.30993327e-07 4.99999997 9.31093327e-07 4.99999997 9.31193327e-07 4.99999997 9.31293327e-07 4.99999997 9.31393327e-07 4.99999997 9.31493327e-07 4.99999997 9.31593327e-07 4.99999997 9.31693327e-07 4.99999997
+ 9.31793327e-07 4.99999997 9.31893327e-07 4.99999997 9.31993327e-07 4.99999997 9.32093327e-07 4.99999997 9.32193327e-07 4.99999997 9.32293327e-07 4.99999997 9.32393327e-07 4.99999997 9.32493327e-07 4.99999997
+ 9.32593327e-07 4.99999997 9.32693327e-07 4.99999997 9.32793327e-07 4.99999997 9.32893327e-07 4.99999997 9.32993327e-07 4.99999997 9.33093327e-07 4.99999997 9.33193327e-07 4.99999997 9.33293327e-07 4.99999997
+ 9.33393327e-07 4.99999997 9.33493327e-07 4.99999997 9.33593327e-07 4.99999997 9.33693327e-07 4.99999997 9.33793327e-07 4.99999997 9.33893327e-07 4.99999997 9.33993327e-07 4.99999997 9.34093327e-07 4.99999997
+ 9.34193327e-07 4.99999997 9.34293327e-07 4.99999997 9.34393327e-07 4.99999997 9.34493327e-07 4.99999997 9.34593327e-07 4.99999997 9.34693327e-07 4.99999997 9.34793327e-07 4.99999997 9.34893327e-07 4.99999997
+ 9.34993327e-07 4.99999997 9.35093327e-07 4.99999997 9.35193327e-07 4.99999997 9.35293327e-07 4.99999997 9.35393327e-07 4.99999997 9.35493327e-07 4.99999997 9.35593327e-07 4.99999997 9.35693327e-07 4.99999997
+ 9.35793327e-07 4.99999997 9.35893327e-07 4.99999997 9.35993327e-07 4.99999997 9.36093327e-07 4.99999997 9.36193327e-07 4.99999997 9.36293327e-07 4.99999997 9.36393327e-07 4.99999997 9.36493327e-07 4.99999997
+ 9.36593327e-07 4.99999997 9.36693327e-07 4.99999997 9.36793327e-07 4.99999997 9.36893327e-07 4.99999997 9.36993327e-07 4.99999997 9.37093327e-07 4.99999997 9.37193327e-07 4.99999997 9.37293327e-07 4.99999997
+ 9.37393327e-07 4.99999997 9.37493327e-07 4.99999997 9.37593327e-07 4.99999997 9.37693327e-07 4.99999997 9.37793327e-07 4.99999997 9.37893327e-07 4.99999997 9.37993327e-07 4.99999997 9.38093327e-07 4.99999997
+ 9.38193327e-07 4.99999997 9.38293327e-07 4.99999997 9.38393327e-07 4.99999997 9.38493327e-07 4.99999997 9.38593327e-07 4.99999997 9.38693327e-07 4.99999997 9.38793327e-07 4.99999997 9.38893327e-07 4.99999997
+ 9.38993327e-07 4.99999997 9.39093327e-07 4.99999997 9.39193327e-07 4.99999997 9.39293327e-07 4.99999997 9.39393327e-07 4.99999997 9.39493327e-07 4.99999997 9.39593327e-07 4.99999997 9.39693327e-07 4.99999997
+ 9.39793327e-07 4.99999997 9.39893327e-07 4.99999997 9.39993327e-07 4.99999997 9.40093327e-07 4.99999997 9.40193327e-07 4.99999997 9.40293327e-07 4.99999997 9.40393327e-07 4.99999997 9.40493327e-07 4.99999997
+ 9.40593327e-07 4.99999997 9.40693327e-07 4.99999997 9.40793327e-07 4.99999997 9.40893327e-07 4.99999997 9.40993327e-07 4.99999997 9.41093327e-07 4.99999997 9.41193327e-07 4.99999997 9.41293327e-07 4.99999997
+ 9.41393327e-07 4.99999997 9.41493327e-07 4.99999997 9.41593327e-07 4.99999997 9.41693327e-07 4.99999997 9.41793327e-07 4.99999997 9.41893327e-07 4.99999997 9.41993327e-07 4.99999997 9.42093327e-07 4.99999997
+ 9.42193327e-07 4.99999997 9.42293327e-07 4.99999997 9.42393327e-07 4.99999997 9.42493327e-07 4.99999997 9.42593327e-07 4.99999997 9.42693327e-07 4.99999997 9.42793327e-07 4.99999997 9.42893327e-07 4.99999997
+ 9.42993327e-07 4.99999997 9.43093327e-07 4.99999997 9.43193327e-07 4.99999997 9.43293327e-07 4.99999997 9.43393327e-07 4.99999997 9.43493327e-07 4.99999997 9.43593327e-07 4.99999997 9.43693327e-07 4.99999997
+ 9.43793327e-07 4.99999997 9.43893327e-07 4.99999997 9.43993327e-07 4.99999997 9.44093327e-07 4.99999997 9.44193327e-07 4.99999997 9.44293327e-07 4.99999997 9.44393327e-07 4.99999997 9.44493327e-07 4.99999997
+ 9.44593327e-07 4.99999997 9.44693327e-07 4.99999997 9.44793327e-07 4.99999997 9.44893327e-07 4.99999997 9.44993327e-07 4.99999997 9.45093327e-07 4.99999997 9.45193327e-07 4.99999997 9.45293327e-07 4.99999997
+ 9.45393327e-07 4.99999997 9.45493327e-07 4.99999997 9.45593327e-07 4.99999997 9.45693327e-07 4.99999997 9.45793327e-07 4.99999997 9.45893327e-07 4.99999997 9.45993327e-07 4.99999997 9.46093327e-07 4.99999997
+ 9.46193327e-07 4.99999997 9.46293327e-07 4.99999997 9.46393327e-07 4.99999997 9.46493327e-07 4.99999997 9.46593327e-07 4.99999997 9.46693327e-07 4.99999997 9.46793327e-07 4.99999997 9.46893327e-07 4.99999997
+ 9.46993327e-07 4.99999997 9.47093327e-07 4.99999997 9.47193327e-07 4.99999997 9.47293327e-07 4.99999997 9.47393327e-07 4.99999997 9.47493327e-07 4.99999997 9.47593327e-07 4.99999997 9.47693327e-07 4.99999997
+ 9.47793327e-07 4.99999997 9.47893327e-07 4.99999997 9.47993327e-07 4.99999997 9.48093327e-07 4.99999997 9.48193327e-07 4.99999997 9.48293327e-07 4.99999997 9.48393327e-07 4.99999997 9.48493327e-07 4.99999997
+ 9.48593327e-07 4.99999997 9.48693327e-07 4.99999997 9.48793327e-07 4.99999997 9.48893327e-07 4.99999997 9.48993327e-07 4.99999997 9.49093327e-07 4.99999997 9.49193327e-07 4.99999997 9.49293327e-07 4.99999997
+ 9.49393327e-07 4.99999997 9.49493327e-07 4.99999997 9.49593327e-07 4.99999997 9.49693327e-07 4.99999997 9.49793327e-07 4.99999997 9.49893327e-07 4.99999997 9.49993327e-07 4.99999997 9.50093327e-07 4.99999997
+ 9.50193327e-07 4.99999997 9.50293327e-07 4.99999997 9.50393327e-07 4.99999997 9.50493327e-07 4.99999997 9.50593327e-07 4.99999997 9.50693327e-07 4.99999997 9.50793327e-07 4.99999997 9.50893327e-07 4.99999997
+ 9.50993327e-07 4.99999997 9.51e-07 4.99999997 9.5101e-07 4.99999997 9.5103e-07 4.99999998 9.5107e-07 4.99999996 9.5115e-07 4.99999998 9.5125e-07 4.99999997 9.5135e-07 4.99999997
+ 9.5145e-07 4.99999998 9.5155e-07 4.99999996 9.5165e-07 4.99999998 9.5175e-07 4.99999996 9.5185e-07 4.99999999 9.51930828e-07 5.00006471 9.52e-07 4.99916174 9.52008608e-07 4.99761843
+ 9.52025825e-07 4.99312395 9.52060258e-07 5.01021614 9.52106188e-07 5.09915398 9.52150118e-07 4.21384241 9.5219811e-07 0.290133164 9.52255501e-07 -0.0555601235 9.52312176e-07 0.071992207 9.52404431e-07 -0.0580455459
+ 9.52490774e-07 0.0521266462 9.52590774e-07 -0.046900588 9.52690774e-07 0.042974581 9.52790774e-07 -0.0387934186 9.52890774e-07 0.0355083829 9.52990774e-07 -0.0321185209 9.53090774e-07 0.0293845439 9.53190774e-07 -0.0266224795
+ 9.53290774e-07 0.0243478875 9.53390774e-07 -0.0220883003 9.53490774e-07 0.0201959102 9.53590774e-07 -0.0183413196 9.53690774e-07 0.0167666634 9.53790774e-07 -0.0152403688 9.53890774e-07 0.0139298139 9.53990774e-07 -0.0126709058
+ 9.54090774e-07 0.0115799054 9.54190774e-07 -0.0105396326 9.54290774e-07 0.00963120539 9.54390774e-07 -0.00877029031 9.54490774e-07 0.00801373348 9.54590774e-07 -0.00730035533 9.54690774e-07 0.00667016991 9.54790774e-07 -0.0060784283
+ 9.54890774e-07 0.00555342785 9.54990774e-07 -0.00506215822 9.55090774e-07 0.00462473134 9.55190774e-07 -0.00421658185 9.55290774e-07 0.00385208255 9.55390774e-07 -0.0035127877 9.55490774e-07 0.00320903124 9.55590774e-07 -0.0029268357
+ 9.55690774e-07 0.00267368149 9.55790774e-07 -0.00243887954 9.55890774e-07 0.00222788568 9.55990774e-07 -0.00203245084 9.56090774e-07 0.0018565878 9.56190774e-07 -0.0016938733 9.56290774e-07 0.00154728638 9.56390774e-07 -0.00141178176
+ 9.56490774e-07 0.00128959387 9.56590774e-07 -0.00117672642 9.56690774e-07 0.00107487425 9.56790774e-07 -0.000980846434 9.56890774e-07 0.000895944254 9.56990774e-07 -0.000817600267 9.57090774e-07 0.000746826659 9.57190774e-07 -0.000681542527
+ 9.57290774e-07 0.000622546127 9.57390774e-07 -0.000568139108 9.57490774e-07 0.000518960166 9.57590774e-07 -0.00047361387 9.57690774e-07 0.000432618935 9.57790774e-07 -0.00039482136 9.57890774e-07 0.000360648892 9.57990774e-07 -0.000329141088
+ 9.58090774e-07 0.000300656148 9.58190774e-07 -0.000274389641 9.58290774e-07 0.000250646154 9.58390774e-07 -0.000228747599 9.58490774e-07 0.0002089569 9.58590774e-07 -0.000190698721 9.58690774e-07 0.000174203358 9.58790774e-07 -0.00015897934
+ 9.58890774e-07 0.000145231232 9.58990774e-07 -0.000132536229 9.59090774e-07 0.000121078462 9.59190774e-07 -0.000110491511 9.59290774e-07 0.000100943174 9.59390774e-07 -9.21134357e-05 9.59490774e-07 8.4156973e-05 9.59590774e-07 -7.67920397e-05
+ 9.59690774e-07 7.01627124e-05 9.59790774e-07 -6.40188597e-05 9.59890774e-07 5.84959595e-05 9.59990774e-07 -5.33700348e-05 9.60090774e-07 4.87695597e-05 9.60190774e-07 -4.44922222e-05 9.60290774e-07 4.06607716e-05 9.60390774e-07 -3.70908606e-05
+ 9.60490774e-07 3.39005457e-05 9.60590774e-07 -3.09203885e-05 9.60690774e-07 2.82645887e-05 9.60790774e-07 -2.57760907e-05 9.60890774e-07 2.3565917e-05 9.60990774e-07 -2.14873027e-05 9.61090774e-07 1.96486482e-05 9.61190774e-07 -1.79117455e-05
+ 9.61290774e-07 1.63828276e-05 9.61390774e-07 -1.49308044e-05 9.61490774e-07 1.36601148e-05 9.61590774e-07 -1.24455918e-05 9.61690774e-07 1.1390188e-05 9.61790774e-07 -1.03736667e-05 9.61890774e-07 9.49774736e-06 9.61990774e-07 -8.6462987e-06
+ 9.62090774e-07 7.9200162e-06 9.62190774e-07 -7.20618766e-06 9.62290774e-07 6.60465801e-06 9.62390774e-07 -6.00556286e-06 9.62490774e-07 5.50804017e-06 9.62590774e-07 -5.004598e-06 9.62690774e-07 4.59378634e-06 9.62790774e-07 -4.17008995e-06
+ 9.62890774e-07 3.83156966e-06 9.62990774e-07 -3.47435733e-06 9.63090774e-07 3.19610667e-06 9.63190774e-07 -2.89432215e-06 9.63290774e-07 2.66631855e-06 9.63390774e-07 -2.41074428e-06 9.63490774e-07 2.22463188e-06 9.63590774e-07 -2.00758319e-06
+ 9.63690774e-07 1.85639569e-06 9.63790774e-07 -1.6714659e-06 9.63890774e-07 1.55939899e-06 9.63990774e-07 -1.38082138e-06 9.64090774e-07 1.30227747e-06 9.64190774e-07 -1.14884092e-06 9.64290774e-07 1.08727392e-06 9.64390774e-07 -9.55390912e-07
+ 9.64490774e-07 9.08044284e-07 9.64590774e-07 -7.94134405e-07 9.64690774e-07 7.58642143e-07 9.64790774e-07 -6.59714463e-07 9.64890774e-07 6.34103635e-07 9.64990774e-07 -5.47664793e-07 9.65090774e-07 5.30290583e-07 9.65190774e-07 -4.54262083e-07
+ 9.65290774e-07 4.43753895e-07 9.65390774e-07 -3.76403601e-07 9.65490774e-07 3.71618865e-07 9.65590774e-07 -3.11502551e-07 9.65690774e-07 3.11488709e-07 9.65790774e-07 -2.57402481e-07 9.65890774e-07 2.61365519e-07 9.65990774e-07 -2.12307012e-07
+ 9.66090774e-07 2.19586255e-07 9.66190774e-07 -1.74727651e-07 9.66290774e-07 1.84780202e-07 9.66390774e-07 -1.43421282e-07 9.66490774e-07 1.55784187e-07 9.66590774e-07 -1.17340694e-07 9.66690774e-07 1.3162823e-07 9.66790774e-07 -9.56134645e-08
+ 9.66890774e-07 1.11504323e-07 9.66990774e-07 -7.75128521e-08 9.67090774e-07 9.47394285e-08 9.67190774e-07 -6.24336459e-08 9.67290774e-07 8.0773134e-08 9.67390774e-07 -4.98334141e-08 9.67490774e-07 6.90993794e-08 9.67590774e-07 -3.93732593e-08
+ 9.67690774e-07 5.94152846e-08 9.67790774e-07 -3.06632475e-08 9.67890774e-07 5.13482989e-08 9.67990774e-07 -2.34074253e-08 9.68090774e-07 4.4628163e-08 9.68190774e-07 -1.73630595e-08 9.68290774e-07 3.90298632e-08 9.68390774e-07 -1.23273488e-08
+ 9.68490774e-07 3.43658604e-08 9.68590774e-07 -8.13252618e-09 9.68690774e-07 3.04809105e-08 9.68790774e-07 -4.6383857e-09 9.68890774e-07 2.72448725e-08 9.68990774e-07 -1.72787004e-09 9.69090774e-07 2.45493399e-08 9.69190774e-07 6.96517594e-10
+ 9.69290774e-07 2.23131571e-08 9.69390774e-07 2.70818332e-09 9.69490774e-07 2.0476404e-08 9.69590774e-07 4.36139957e-09 9.69690774e-07 1.89668154e-08 9.69790774e-07 5.72018077e-09 9.69890774e-07 1.77260565e-08 9.69990774e-07 6.83700865e-09
+ 9.70090774e-07 1.67062181e-08 9.70190774e-07 7.75499584e-09 9.70290774e-07 1.58679406e-08 9.70390774e-07 8.50956478e-09 9.70490774e-07 1.50799962e-08 9.70590774e-07 9.11601317e-09 9.70690774e-07 1.45257675e-08 9.70790774e-07 9.61910643e-09
+ 9.70890774e-07 1.40694267e-08 9.70990774e-07 1.00330061e-08 9.71090774e-07 1.36940246e-08 9.71190774e-07 1.03734906e-08 9.71290774e-07 1.33852096e-08 9.71390774e-07 1.06535815e-08 9.71490774e-07 1.31311713e-08 9.71590774e-07 1.08839909e-08
+ 9.71690774e-07 1.2922193e-08 9.71790774e-07 1.10735315e-08 9.71890774e-07 1.27502823e-08 9.71990774e-07 1.12294522e-08 9.72090774e-07 1.26088638e-08 9.72190774e-07 1.13577175e-08 9.72290774e-07 1.24925288e-08 9.72390774e-07 1.14632322e-08
+ 9.72490774e-07 1.23968276e-08 9.72590774e-07 1.15500324e-08 9.72690774e-07 1.23181003e-08 9.72790774e-07 1.16214378e-08 9.72890774e-07 1.22533358e-08 9.72990774e-07 1.16801792e-08 9.73090774e-07 1.2200057e-08 9.73190774e-07 1.17285029e-08
+ 9.73290774e-07 1.21562274e-08 9.73390774e-07 1.17682568e-08 9.73490774e-07 1.212017e-08 9.73590774e-07 1.18009615e-08 9.73690774e-07 1.20905067e-08 9.73790774e-07 1.18278667e-08 9.73890774e-07 1.20661032e-08 9.73990774e-07 1.18500012e-08
+ 9.74090774e-07 1.20460264e-08 9.74190774e-07 1.18682112e-08 9.74290774e-07 1.20295095e-08 9.74390774e-07 1.18831928e-08 9.74490774e-07 1.20159205e-08 9.74590774e-07 1.18955188e-08 9.74690774e-07 1.20047403e-08 9.74790774e-07 1.19056595e-08
+ 9.74890774e-07 1.1995542e-08 9.74990774e-07 1.19140032e-08 9.75090774e-07 1.19879736e-08 9.75190774e-07 1.19208679e-08 9.75290774e-07 1.19817468e-08 9.75390774e-07 1.19265163e-08 9.75490774e-07 1.19766235e-08 9.75590774e-07 1.19311635e-08
+ 9.75690774e-07 1.19724074e-08 9.75790774e-07 1.19349879e-08 9.75890774e-07 1.19689388e-08 9.75990774e-07 1.19381347e-08 9.76090774e-07 1.19660842e-08 9.76190774e-07 1.19407246e-08 9.76290774e-07 1.19637349e-08 9.76390774e-07 1.19428557e-08
+ 9.76490774e-07 1.19618013e-08 9.76590774e-07 1.19446092e-08 9.76690774e-07 1.19602104e-08 9.76790774e-07 1.19460527e-08 9.76890774e-07 1.1958901e-08 9.76990774e-07 1.19472407e-08 9.77090774e-07 1.19578234e-08 9.77190774e-07 1.19482187e-08
+ 9.77290774e-07 1.19569359e-08 9.77390774e-07 1.19490237e-08 9.77490774e-07 1.19562054e-08 9.77590774e-07 1.19496865e-08 9.77690774e-07 1.19556042e-08 9.77790774e-07 1.19502319e-08 9.77890774e-07 1.19551089e-08 9.77990774e-07 1.19506812e-08
+ 9.78090774e-07 1.19547013e-08 9.78190774e-07 1.19510511e-08 9.78290774e-07 1.19543659e-08 9.78390774e-07 1.19513556e-08 9.78490774e-07 1.19540894e-08 9.78590774e-07 1.19516065e-08 9.78690774e-07 1.19538617e-08 9.78790774e-07 1.1951813e-08
+ 9.78890774e-07 1.19536742e-08 9.78990774e-07 1.19519835e-08 9.79090774e-07 1.19535195e-08 9.79190774e-07 1.19521238e-08 9.79290774e-07 1.19533922e-08 9.79390774e-07 1.19522396e-08 9.79490774e-07 1.1953287e-08 9.79590774e-07 1.1952335e-08
+ 9.79690774e-07 1.19532002e-08 9.79790774e-07 1.19524136e-08 9.79890774e-07 1.19531291e-08 9.79990774e-07 1.19524781e-08 9.80090774e-07 1.19530704e-08 9.80190774e-07 1.19525316e-08 9.80290774e-07 1.19530218e-08 9.80390774e-07 1.19525759e-08
+ 9.80490774e-07 1.19529817e-08 9.80590774e-07 1.19526123e-08 9.80690774e-07 1.19529488e-08 9.80790774e-07 1.19526425e-08 9.80890774e-07 1.19529213e-08 9.80990774e-07 1.19526671e-08 9.81090774e-07 1.19528986e-08 9.81190774e-07 1.19526877e-08
+ 9.81290774e-07 1.19528799e-08 9.81390774e-07 1.19527047e-08 9.81490774e-07 1.19528645e-08 9.81590774e-07 1.1952719e-08 9.81690774e-07 1.19528518e-08 9.81790774e-07 1.19527305e-08 9.81890774e-07 1.19528411e-08 9.81990774e-07 1.19527405e-08
+ 9.82090774e-07 1.19528322e-08 9.82190774e-07 1.19527481e-08 9.82290774e-07 1.19528249e-08 9.82390774e-07 1.19527548e-08 9.82490774e-07 1.1952819e-08 9.82590774e-07 1.19527604e-08 9.82690774e-07 1.19528143e-08 9.82790774e-07 1.19527648e-08
+ 9.82890774e-07 1.19528102e-08 9.82990774e-07 1.19527685e-08 9.83090774e-07 1.19528064e-08 9.83190774e-07 1.19527717e-08 9.83290774e-07 1.19528034e-08 9.83390774e-07 1.19527742e-08 9.83490774e-07 1.19528011e-08 9.83590774e-07 1.19527765e-08
+ 9.83690774e-07 1.19527991e-08 9.83790774e-07 1.1952778e-08 9.83890774e-07 1.19527978e-08 9.83990774e-07 1.19527795e-08 9.84090774e-07 1.19527963e-08 9.84190774e-07 1.19527812e-08 9.84290774e-07 1.19527949e-08 9.84390774e-07 1.19527823e-08
+ 9.84490774e-07 1.1952794e-08 9.84590774e-07 1.19527833e-08 9.84690774e-07 1.19527931e-08 9.84790774e-07 1.19527838e-08 9.84890774e-07 1.19527926e-08 9.84990774e-07 1.19527845e-08 9.85090774e-07 1.19527918e-08 9.85190774e-07 1.1952785e-08
+ 9.85290774e-07 1.19527913e-08 9.85390774e-07 1.19527855e-08 9.85490774e-07 1.19527909e-08 9.85590774e-07 1.1952786e-08 9.85690774e-07 1.19527904e-08 9.85790774e-07 1.19527865e-08 9.85890774e-07 1.19527899e-08 9.85990774e-07 1.19527868e-08
+ 9.86090774e-07 1.19527899e-08 9.86190774e-07 1.19527868e-08 9.86290774e-07 1.195279e-08 9.86390774e-07 1.19527868e-08 9.86490774e-07 1.195279e-08 9.86590774e-07 1.19527868e-08 9.86690774e-07 1.19527897e-08 9.86790774e-07 1.19527869e-08
+ 9.86890774e-07 1.19527896e-08 9.86990774e-07 1.1952787e-08 9.87090774e-07 1.19527894e-08 9.87190774e-07 1.1952787e-08 9.87290774e-07 1.19527897e-08 9.87390774e-07 1.19527871e-08 9.87490774e-07 1.19527893e-08 9.87590774e-07 1.19527872e-08
+ 9.87690774e-07 1.19527895e-08 9.87790774e-07 1.19527874e-08 9.87890774e-07 1.19527891e-08 9.87990774e-07 1.19527874e-08 9.88090774e-07 1.19527891e-08 9.88190774e-07 1.19527876e-08 9.88290774e-07 1.1952789e-08 9.88390774e-07 1.19527878e-08
+ 9.88490774e-07 1.1952789e-08 9.88590774e-07 1.19527878e-08 9.88690774e-07 1.19527889e-08 9.88790774e-07 1.19527879e-08 9.88890774e-07 1.1952789e-08 9.88990774e-07 1.19527878e-08 9.89090774e-07 1.19527888e-08 9.89190774e-07 1.19527878e-08
+ 9.89290774e-07 1.19527889e-08 9.89390774e-07 1.19527879e-08 9.89490774e-07 1.19527889e-08 9.89590774e-07 1.1952788e-08 9.89690774e-07 1.19527889e-08 9.89790774e-07 1.1952788e-08 9.89890774e-07 1.19527888e-08 9.89990774e-07 1.1952788e-08
+ 9.90090774e-07 1.19527889e-08 9.90190774e-07 1.1952788e-08 9.90290774e-07 1.19527888e-08 9.90390774e-07 1.1952788e-08 9.90490774e-07 1.19527888e-08 9.90590774e-07 1.19527881e-08 9.90690774e-07 1.19527887e-08 9.90790774e-07 1.1952788e-08
+ 9.90890774e-07 1.19527888e-08 9.90990774e-07 1.1952788e-08 9.91090774e-07 1.19527888e-08 9.91190774e-07 1.19527879e-08 9.91290774e-07 1.19527888e-08 9.91390774e-07 1.19527881e-08 9.91490774e-07 1.19527887e-08 9.91590774e-07 1.19527881e-08
+ 9.91690774e-07 1.19527887e-08 9.91790774e-07 1.19527881e-08 9.91890774e-07 1.19527887e-08 9.91990774e-07 1.19527882e-08 9.92090774e-07 1.19527885e-08 9.92190774e-07 1.19527882e-08 9.92290774e-07 1.19527886e-08 9.92390774e-07 1.19527883e-08
+ 9.92490774e-07 1.19527886e-08 9.92590774e-07 1.19527881e-08 9.92690774e-07 1.19527886e-08 9.92790774e-07 1.19527883e-08 9.92890774e-07 1.19527885e-08 9.92990774e-07 1.19527881e-08 9.93090774e-07 1.19527886e-08 9.93190774e-07 1.19527882e-08
+ 9.93290774e-07 1.19527885e-08 9.93390774e-07 1.19527882e-08 9.93490774e-07 1.19527885e-08 9.93590774e-07 1.19527882e-08 9.93690774e-07 1.19527885e-08 9.93790774e-07 1.19527882e-08 9.93890774e-07 1.19527885e-08 9.93990774e-07 1.19527882e-08
+ 9.94090774e-07 1.19527885e-08 9.94190774e-07 1.19527882e-08 9.94290774e-07 1.19527885e-08 9.94390774e-07 1.19527882e-08 9.94490774e-07 1.19527885e-08 9.94590774e-07 1.19527882e-08 9.94690774e-07 1.19527885e-08 9.94790774e-07 1.19527882e-08
+ 9.94890774e-07 1.19527885e-08 9.94990774e-07 1.19527882e-08 9.95090774e-07 1.19527885e-08 9.95190774e-07 1.19527882e-08 9.95290774e-07 1.19527885e-08 9.95390774e-07 1.19527882e-08 9.95490774e-07 1.19527885e-08 9.95590774e-07 1.19527882e-08
+ 9.95690774e-07 1.19527886e-08 9.95790774e-07 1.19527883e-08 9.95890774e-07 1.19527884e-08 9.95990774e-07 1.19527883e-08 9.96090774e-07 1.19527885e-08 9.96190774e-07 1.19527883e-08 9.96290774e-07 1.19527885e-08 9.96390774e-07 1.19527883e-08
+ 9.96490774e-07 1.19527885e-08 9.96590774e-07 1.19527883e-08 9.96690774e-07 1.19527885e-08 9.96790774e-07 1.19527883e-08 9.96890774e-07 1.19527885e-08 9.96990774e-07 1.19527883e-08 9.97090774e-07 1.19527885e-08 9.97190774e-07 1.19527883e-08
+ 9.97290774e-07 1.19527885e-08 9.97390774e-07 1.19527883e-08 9.97490774e-07 1.19527885e-08 9.97590774e-07 1.19527883e-08 9.97690774e-07 1.19527885e-08 9.97790774e-07 1.19527883e-08 9.97890774e-07 1.19527885e-08 9.97990774e-07 1.19527883e-08
+ 9.98090774e-07 1.19527885e-08 9.98190774e-07 1.19527883e-08 9.98290774e-07 1.19527885e-08 9.98390774e-07 1.19527883e-08 9.98490774e-07 1.19527885e-08 9.98590774e-07 1.19527883e-08 9.98690774e-07 1.19527885e-08 9.98790774e-07 1.19527883e-08
+ 9.98890774e-07 1.19527885e-08 9.98990774e-07 1.19527883e-08 9.99090774e-07 1.19527885e-08 9.99190774e-07 1.19527883e-08 9.99290774e-07 1.19527885e-08 9.99390774e-07 1.19527883e-08 9.99490774e-07 1.19527885e-08 9.99590774e-07 1.19527883e-08
+ 9.99690774e-07 1.19527885e-08 9.99790774e-07 1.19527883e-08 9.99890774e-07 1.19527885e-08 9.99990774e-07 1.19527883e-08 1e-06 1.19527881e-08 )

Vclkin2 in2 0 PWL( 0.0 1.19527881e-08 1e-12 1.24792718e-08 2e-12 1.25186848e-08 4e-12 1.21631176e-08 8e-12 1.12795195e-08 1.6e-11 1.18109305e-08 3.2e-11 1.23719842e-08 6.4e-11 1.16333275e-08
+ 1.28e-10 1.21770584e-08 2.28e-10 1.17852892e-08 3.28e-10 1.20753204e-08 4.28e-10 1.18612976e-08 5.28e-10 1.20299297e-08 6.28e-10 1.18245968e-08 7.28e-10 1.38600423e-08 8.17641203e-10 -4.02920994e-07
+ 8.87939724e-10 3.97836068e-06 9.63955785e-10 -2.00790766e-06 1e-09 -3.65992502e-05 1.00713579e-09 -3.91179359e-06 1.02140738e-09 7.54784841e-06 1.04995055e-09 7.88235786e-06 1.09557449e-09 1.08375649e-05 1.1454732e-09 -7.23832858e-07
+ 1.21884515e-09 -8.61866769e-06 1.31884515e-09 5.17990034e-06 1.41884515e-09 -1.52120962e-06 1.51884515e-09 2.33511653e-07 1.61884515e-09 4.01624692e-07 1.71884515e-09 -6.92434146e-07 1.81884515e-09 8.89819171e-07 1.91884515e-09 -9.63936286e-07
+ 2.01884515e-09 1.03919308e-06 2.11884515e-09 -1.03623834e-06 2.21884515e-09 1.05968371e-06 2.31884515e-09 -1.01993892e-06 2.41884515e-09 1.01713978e-06 2.51884515e-09 -9.58452698e-07 2.61884515e-09 9.42421307e-07 2.71884515e-09 -8.74722477e-07
+ 2.81884515e-09 8.53062973e-07 2.91884515e-09 -7.82296098e-07 3.01884515e-09 7.59588916e-07 3.11884515e-09 -6.89314803e-07 3.21884515e-09 6.68262018e-07 3.31884515e-09 -6.00529173e-07 3.41884515e-09 5.82629049e-07 3.51884515e-09 -5.1851424e-07
+ 3.61884515e-09 5.0449337e-07 3.71884515e-09 -4.41670007e-07 3.81884515e-09 4.37771547e-07 3.91884515e-09 -3.76004654e-07 4.01884515e-09 3.75519474e-07 4.11884515e-09 -3.18601286e-07 4.21884515e-09 3.21152194e-07 4.31884515e-09 -2.68691983e-07
+ 4.41884515e-09 2.74063803e-07 4.51884515e-09 -2.2561747e-07 4.61884515e-09 2.33549616e-07 4.71884515e-09 -1.88658673e-07 4.81884515e-09 1.98872911e-07 4.91884515e-09 -1.57094897e-07 5.01884515e-09 1.69316027e-07 5.11884515e-09 -1.30239202e-07
+ 5.21884515e-09 1.44208636e-07 5.31884515e-09 -1.07460078e-07 5.41884515e-09 1.22940825e-07 5.51884515e-09 -8.81882992e-08 5.61884515e-09 1.04967793e-07 5.71884515e-09 -7.19185811e-08 5.81884515e-09 8.98081736e-08 5.91884515e-09 -5.82103102e-08
+ 6.01884515e-09 7.7047931e-08 6.11884515e-09 -4.66795699e-08 6.21884515e-09 6.63219972e-08 6.31884515e-09 -3.69933403e-08 6.41884515e-09 5.73169687e-08 6.51884515e-09 -2.88653901e-08 6.61884515e-09 4.97638871e-08 6.71884515e-09 -2.20504009e-08
+ 6.81884515e-09 4.34329868e-08 6.91884515e-09 -1.63400911e-08 7.01884515e-09 3.81300682e-08 7.11884515e-09 -1.15448655e-08 7.21884515e-09 3.36782729e-08 7.31884515e-09 -7.54564888e-09 7.41884515e-09 2.99660583e-08 7.51884515e-09 -4.19998974e-09
+ 7.61884515e-09 2.68613089e-08 7.71884515e-09 -1.40219222e-09 7.81884515e-09 2.42653431e-08 7.91884515e-09 9.36803607e-10 8.01884515e-09 2.21075072e-08 8.11884515e-09 2.88145136e-09 8.21884515e-09 2.03288801e-08 8.31884515e-09 4.48488657e-09
+ 8.41884515e-09 1.88624873e-08 8.51884515e-09 5.80674178e-09 8.61884515e-09 1.76536916e-08 8.71884515e-09 6.89631979e-09 8.81884515e-09 1.66573664e-08 8.91884515e-09 7.79433357e-09 9.01884515e-09 1.58362513e-08 9.11884515e-09 8.53438836e-09
+ 9.21884515e-09 1.50615762e-08 9.31884515e-09 9.13027823e-09 9.41884515e-09 1.45153982e-08 9.51884515e-09 9.62617902e-09 9.61884515e-09 1.40651079e-08 9.71884515e-09 1.00350389e-08 9.81884515e-09 1.36938755e-08 9.91884515e-09 1.03721003e-08
+ 1.00188451e-08 1.33878439e-08 1.01188451e-08 1.0649955e-08 1.02188451e-08 1.31355751e-08 1.03188451e-08 1.08789918e-08 1.04188451e-08 1.29276326e-08 1.05188451e-08 1.1067781e-08 1.06188451e-08 1.2756234e-08 1.07188451e-08 1.12233905e-08
+ 1.08188451e-08 1.26149608e-08 1.09188451e-08 1.13516473e-08 1.10188451e-08 1.2498521e-08 1.11188451e-08 1.14573578e-08 1.12188451e-08 1.24025519e-08 1.13188451e-08 1.15444831e-08 1.14188451e-08 1.23234558e-08 1.15188451e-08 1.16162896e-08
+ 1.16188451e-08 1.2258267e-08 1.17188451e-08 1.16754706e-08 1.18188451e-08 1.22045412e-08 1.19188451e-08 1.1724244e-08 1.20188451e-08 1.2160263e-08 1.21188451e-08 1.17644408e-08 1.22188451e-08 1.21237717e-08 1.23188451e-08 1.17975681e-08
+ 1.24188451e-08 1.2093698e-08 1.25188451e-08 1.18248696e-08 1.26188451e-08 1.20689136e-08 1.27188451e-08 1.18473697e-08 1.28188451e-08 1.20484878e-08 1.29188451e-08 1.18659123e-08 1.30188451e-08 1.20316546e-08 1.31188451e-08 1.18811934e-08
+ 1.32188451e-08 1.20177822e-08 1.33188451e-08 1.18937866e-08 1.34188451e-08 1.20063498e-08 1.35188451e-08 1.19041653e-08 1.36188451e-08 1.19969286e-08 1.37188451e-08 1.19127177e-08 1.38188451e-08 1.19891642e-08 1.39188451e-08 1.19197663e-08
+ 1.40188451e-08 1.19827653e-08 1.41188451e-08 1.19255752e-08 1.42188451e-08 1.19774923e-08 1.43188451e-08 1.19303619e-08 1.44188451e-08 1.19731467e-08 1.45188451e-08 1.19343068e-08 1.46188451e-08 1.19695658e-08 1.47188451e-08 1.19375577e-08
+ 1.48188451e-08 1.19666145e-08 1.49188451e-08 1.19402367e-08 1.50188451e-08 1.19641827e-08 1.51188451e-08 1.19424444e-08 1.52188451e-08 1.19621782e-08 1.53188451e-08 1.19442641e-08 1.54188451e-08 1.19605267e-08 1.55188451e-08 1.19457636e-08
+ 1.56188451e-08 1.1959165e-08 1.57188451e-08 1.19469991e-08 1.58188451e-08 1.19580437e-08 1.59188451e-08 1.19480176e-08 1.60188451e-08 1.19571193e-08 1.61188451e-08 1.19488567e-08 1.62188451e-08 1.19563575e-08 1.63188451e-08 1.19495481e-08
+ 1.64188451e-08 1.19557297e-08 1.65188451e-08 1.19501183e-08 1.66188451e-08 1.19552122e-08 1.67188451e-08 1.19505878e-08 1.68188451e-08 1.19547856e-08 1.69188451e-08 1.19509748e-08 1.70188451e-08 1.19544345e-08 1.71188451e-08 1.19512939e-08
+ 1.72188451e-08 1.19541446e-08 1.73188451e-08 1.19515569e-08 1.74188451e-08 1.19539062e-08 1.75188451e-08 1.19517733e-08 1.76188451e-08 1.19537095e-08 1.77188451e-08 1.19519517e-08 1.78188451e-08 1.19535477e-08 1.79188451e-08 1.19520987e-08
+ 1.80188451e-08 1.1953414e-08 1.81188451e-08 1.19522202e-08 1.82188451e-08 1.19533043e-08 1.83188451e-08 1.19523199e-08 1.84188451e-08 1.19532137e-08 1.85188451e-08 1.19524022e-08 1.86188451e-08 1.19531387e-08 1.87188451e-08 1.19524701e-08
+ 1.88188451e-08 1.19530771e-08 1.89188451e-08 1.19525261e-08 1.90188451e-08 1.19530263e-08 1.91188451e-08 1.19525723e-08 1.92188451e-08 1.19529845e-08 1.93188451e-08 1.19526101e-08 1.94188451e-08 1.195295e-08 1.95188451e-08 1.19526415e-08
+ 1.96188451e-08 1.19529215e-08 1.97188451e-08 1.19526673e-08 1.98188451e-08 1.1952898e-08 1.99188451e-08 1.19526885e-08 2e-08 1.19528767e-08 2.001e-08 3.86449984e-07 2.003e-08 -7.32508179e-07 2.007e-08 4.33825947e-09
+ 2.01e-08 1.15037632e-06 2.0108e-08 5.11179698e-06 2.0124e-08 8.89352763e-06 2.0156e-08 3.28123757e-07 2.02150599e-08 -1.37064563e-05 2.02823902e-08 9.68117413e-06 2.03483061e-08 -8.04395084e-06 2.04483061e-08 1.50420703e-05
+ 2.05483061e-08 -1.81591237e-05 2.06483061e-08 1.72259796e-05 2.07483061e-08 -1.59084351e-05 2.08483061e-08 1.45544798e-05 2.09483061e-08 -1.31529412e-05 2.10483061e-08 1.18735067e-05 2.11483061e-08 -1.06273411e-05 2.12483061e-08 9.53761307e-06
+ 2.13483061e-08 -8.49352239e-06 2.14483061e-08 7.60191331e-06 2.15483061e-08 -6.74784198e-06 2.16483061e-08 6.03193237e-06 2.17483061e-08 -5.34062261e-06 2.18483061e-08 4.77200309e-06 2.19483061e-08 -4.21510775e-06 2.20483061e-08 3.76689589e-06
+ 2.21483061e-08 -3.31909263e-06 2.22483061e-08 2.96809459e-06 2.23483061e-08 -2.60802067e-06 2.24483061e-08 2.33495561e-06 2.25483061e-08 -2.04503963e-06 2.26483061e-08 1.83417638e-06 2.27483061e-08 -1.60016532e-06 2.28483061e-08 1.43879842e-06
+ 2.29483061e-08 -1.24921924e-06 2.30483061e-08 1.1271487e-06 2.31483061e-08 -9.72810863e-07 2.32483061e-08 8.81880608e-07 2.33483061e-08 -7.55446402e-07 2.34483061e-08 6.89153224e-07 2.35483061e-08 -5.84778719e-07 2.36483061e-08 5.37948622e-07
+ 2.37483061e-08 -4.50988692e-07 2.38483061e-08 4.19512576e-07 2.39483061e-08 -3.46281091e-07 2.40483061e-08 3.26900628e-07 2.41483061e-08 -2.64476717e-07 2.42483061e-08 2.5461127e-07 2.43483061e-08 -2.00681834e-07 2.44483061e-08 1.98288955e-07
+ 2.45483061e-08 -1.51026451e-07 2.46483061e-08 1.54494925e-07 2.47483061e-08 -1.12458299e-07 2.48483061e-08 1.20517851e-07 2.49483061e-08 -8.25714142e-08 2.50483061e-08 9.42214333e-08 2.51483061e-08 -5.94699266e-08 2.52483061e-08 7.39209906e-08
+ 2.53483061e-08 -4.16603103e-08 2.54483061e-08 5.82936221e-08 2.55483061e-08 -2.79721057e-08 2.56483061e-08 4.63030894e-08 2.57483061e-08 -1.74885073e-08 2.58483061e-08 3.73635501e-08 2.59483061e-08 -9.37963068e-09 2.60483061e-08 3.03288909e-08
+ 2.61483061e-08 -3.34159528e-09 2.62483061e-08 2.50022764e-08 2.63483061e-08 1.21735225e-09 2.64483061e-08 2.10178148e-08 2.65483061e-08 4.61614585e-09 2.66483061e-08 1.80670574e-08 2.67483061e-08 7.12300333e-09 2.68483061e-08 1.59120002e-08
+ 2.69483061e-08 8.94344557e-09 2.70483061e-08 1.42640828e-08 2.71483061e-08 1.02348574e-08 2.72483061e-08 1.31728762e-08 2.73483061e-08 1.11482246e-08 2.74483061e-08 1.24127337e-08 2.75483061e-08 1.17765964e-08 2.76483061e-08 1.1897372e-08
+ 2.77483061e-08 1.21953285e-08 2.78483061e-08 1.15610448e-08 2.79483061e-08 1.24615614e-08 2.80483061e-08 1.13542415e-08 2.81483061e-08 1.26181253e-08 2.82483061e-08 1.12399789e-08 2.83483061e-08 1.26969505e-08 2.84483061e-08 1.11906641e-08
+ 2.85483061e-08 1.27218672e-08 2.86483061e-08 1.11857163e-08 2.87483061e-08 1.27105445e-08 2.88483061e-08 1.1210193e-08 2.89483061e-08 1.26757752e-08 2.90483061e-08 1.12528034e-08 2.91483061e-08 1.26272461e-08 2.92483061e-08 1.13056557e-08
+ 2.93483061e-08 1.25714118e-08 2.94483061e-08 1.13633543e-08 2.95483061e-08 1.2512622e-08 2.96483061e-08 1.14225253e-08 2.97483061e-08 1.24539498e-08 2.98483061e-08 1.14801615e-08 2.99483061e-08 1.23976145e-08 3.00483061e-08 1.15348899e-08
+ 3.01483061e-08 1.23447203e-08 3.02483061e-08 1.15857474e-08 3.03483061e-08 1.22960881e-08 3.04483061e-08 1.16320757e-08 3.05483061e-08 1.22520417e-08 3.06483061e-08 1.16738829e-08 3.07483061e-08 1.22124487e-08 3.08483061e-08 1.17112875e-08
+ 3.09483061e-08 1.21771885e-08 3.10483061e-08 1.17444609e-08 3.11483061e-08 1.21460337e-08 3.12483061e-08 1.17736726e-08 3.13483061e-08 1.21186849e-08 3.14483061e-08 1.1799242e-08 3.15483061e-08 1.20948098e-08 3.16483061e-08 1.18215075e-08
+ 3.17483061e-08 1.20740714e-08 3.18483061e-08 1.18408025e-08 3.19483061e-08 1.20561331e-08 3.20483061e-08 1.18574672e-08 3.21483061e-08 1.20406646e-08 3.22483061e-08 1.18718128e-08 3.23483061e-08 1.20273716e-08 3.24483061e-08 1.18841215e-08
+ 3.25483061e-08 1.20159826e-08 3.26483061e-08 1.18946532e-08 3.27483061e-08 1.20062486e-08 3.28483061e-08 1.19036447e-08 3.29483061e-08 1.1997948e-08 3.30483061e-08 1.19113023e-08 3.31483061e-08 1.19908877e-08 3.32483061e-08 1.19178091e-08
+ 3.33483061e-08 1.19848931e-08 3.34483061e-08 1.19233297e-08 3.35483061e-08 1.19798118e-08 3.36483061e-08 1.19280056e-08 3.37483061e-08 1.19755105e-08 3.38483061e-08 1.19319605e-08 3.39483061e-08 1.19718753e-08 3.40483061e-08 1.19353007e-08
+ 3.41483061e-08 1.19688067e-08 3.42483061e-08 1.19381186e-08 3.43483061e-08 1.19662197e-08 3.44483061e-08 1.19404925e-08 3.45483061e-08 1.19640415e-08 3.46483061e-08 1.19424911e-08 3.47483061e-08 1.19622088e-08 3.48483061e-08 1.19441713e-08
+ 3.49483061e-08 1.1960669e-08 3.50483061e-08 1.19455826e-08 3.51483061e-08 1.1959376e-08 3.52483061e-08 1.19467665e-08 3.53483061e-08 1.19582915e-08 3.54483061e-08 1.19477598e-08 3.55483061e-08 1.19573823e-08 3.56483061e-08 1.19485921e-08
+ 3.57483061e-08 1.19566207e-08 3.58483061e-08 1.19492889e-08 3.59483061e-08 1.19559832e-08 3.60483061e-08 1.19498719e-08 3.61483061e-08 1.19554499e-08 3.62483061e-08 1.19503596e-08 3.63483061e-08 1.1955004e-08 3.64483061e-08 1.1950767e-08
+ 3.65483061e-08 1.19546318e-08 3.66483061e-08 1.19511069e-08 3.67483061e-08 1.19543213e-08 3.68483061e-08 1.19513905e-08 3.69483061e-08 1.19540623e-08 3.70483061e-08 1.19516271e-08 3.71483061e-08 1.19538464e-08 3.72483061e-08 1.19518242e-08
+ 3.73483061e-08 1.19536668e-08 3.74483061e-08 1.19519881e-08 3.75483061e-08 1.19535172e-08 3.76483061e-08 1.19521246e-08 3.77483061e-08 1.19533926e-08 3.78483061e-08 1.19522378e-08 3.79483061e-08 1.19532894e-08 3.80483061e-08 1.19523321e-08
+ 3.81483061e-08 1.19532035e-08 3.82483061e-08 1.19524106e-08 3.83483061e-08 1.19531325e-08 3.84483061e-08 1.19524754e-08 3.85483061e-08 1.19530733e-08 3.86483061e-08 1.1952529e-08 3.87483061e-08 1.19530241e-08 3.88483061e-08 1.19525737e-08
+ 3.89483061e-08 1.19529835e-08 3.90483061e-08 1.19526107e-08 3.91483061e-08 1.19529498e-08 3.92483061e-08 1.19526414e-08 3.93483061e-08 1.1952922e-08 3.94483061e-08 1.19526666e-08 3.95483061e-08 1.19528989e-08 3.96483061e-08 1.19526875e-08
+ 3.97483061e-08 1.19528798e-08 3.98483061e-08 1.19527049e-08 3.99483061e-08 1.19528639e-08 4.00483061e-08 1.19527196e-08 4.01483061e-08 1.1952851e-08 4.02483061e-08 1.19527314e-08 4.03483061e-08 1.19528397e-08 4.04483061e-08 1.19527412e-08
+ 4.05483061e-08 1.19528308e-08 4.06483061e-08 1.19527495e-08 4.07483061e-08 1.19528237e-08 4.08483061e-08 1.19527564e-08 4.09483061e-08 1.19528174e-08 4.10483061e-08 1.19527618e-08 4.11483061e-08 1.19528125e-08 4.12483061e-08 1.19527665e-08
+ 4.13483061e-08 1.19528082e-08 4.14483061e-08 1.19527704e-08 4.15483061e-08 1.19528046e-08 4.16483061e-08 1.19527734e-08 4.17483061e-08 1.19528018e-08 4.18483061e-08 1.19527761e-08 4.19483061e-08 1.19527995e-08 4.20483061e-08 1.19527783e-08
+ 4.21483061e-08 1.19527973e-08 4.22483061e-08 1.195278e-08 4.23483061e-08 1.19527958e-08 4.24483061e-08 1.19527816e-08 4.25483061e-08 1.19527944e-08 4.26483061e-08 1.19527827e-08 4.27483061e-08 1.19527932e-08 4.28483061e-08 1.19527839e-08
+ 4.29483061e-08 1.19527924e-08 4.30483061e-08 1.19527848e-08 4.31483061e-08 1.19527921e-08 4.32483061e-08 1.1952785e-08 4.33483061e-08 1.19527912e-08 4.34483061e-08 1.19527857e-08 4.35483061e-08 1.19527906e-08 4.36483061e-08 1.19527861e-08
+ 4.37483061e-08 1.19527899e-08 4.38483061e-08 1.19527866e-08 4.39483061e-08 1.19527897e-08 4.40483061e-08 1.19527869e-08 4.41483061e-08 1.19527897e-08 4.42483061e-08 1.19527872e-08 4.43483061e-08 1.19527893e-08 4.44483061e-08 1.19527873e-08
+ 4.45483061e-08 1.19527893e-08 4.46483061e-08 1.19527872e-08 4.47483061e-08 1.19527894e-08 4.48483061e-08 1.19527875e-08 4.49483061e-08 1.19527891e-08 4.50483061e-08 1.19527874e-08 4.51483061e-08 1.1952789e-08 4.52483061e-08 1.19527877e-08
+ 4.53483061e-08 1.1952789e-08 4.54483061e-08 1.19527878e-08 4.55483061e-08 1.1952789e-08 4.56483061e-08 1.19527877e-08 4.57483061e-08 1.19527891e-08 4.58483061e-08 1.19527876e-08 4.59483061e-08 1.19527889e-08 4.60483061e-08 1.19527876e-08
+ 4.61483061e-08 1.19527886e-08 4.62483061e-08 1.1952788e-08 4.63483061e-08 1.19527886e-08 4.64483061e-08 1.19527881e-08 4.65483061e-08 1.19527888e-08 4.66483061e-08 1.19527881e-08 4.67483061e-08 1.19527887e-08 4.68483061e-08 1.1952788e-08
+ 4.69483061e-08 1.19527888e-08 4.70483061e-08 1.19527879e-08 4.71483061e-08 1.19527887e-08 4.72483061e-08 1.1952788e-08 4.73483061e-08 1.19527885e-08 4.74483061e-08 1.19527878e-08 4.75483061e-08 1.19527886e-08 4.76483061e-08 1.19527879e-08
+ 4.77483061e-08 1.19527888e-08 4.78483061e-08 1.19527878e-08 4.79483061e-08 1.19527886e-08 4.80483061e-08 1.19527879e-08 4.81483061e-08 1.19527889e-08 4.82483061e-08 1.19527878e-08 4.83483061e-08 1.19527888e-08 4.84483061e-08 1.1952788e-08
+ 4.85483061e-08 1.19527888e-08 4.86483061e-08 1.19527879e-08 4.87483061e-08 1.19527889e-08 4.88483061e-08 1.19527878e-08 4.89483061e-08 1.1952789e-08 4.90483061e-08 1.19527877e-08 4.91483061e-08 1.19527888e-08 4.92483061e-08 1.19527881e-08
+ 4.93483061e-08 1.19527886e-08 4.94483061e-08 1.19527881e-08 4.95483061e-08 1.19527888e-08 4.96483061e-08 1.19527879e-08 4.97483061e-08 1.19527886e-08 4.98483061e-08 1.19527881e-08 4.99483061e-08 1.19527886e-08 5.00483061e-08 1.19527882e-08
+ 5.01483061e-08 1.19527885e-08 5.02483061e-08 1.1952788e-08 5.03483061e-08 1.19527883e-08 5.04483061e-08 1.1952788e-08 5.05483061e-08 1.19527883e-08 5.06483061e-08 1.1952788e-08 5.07483061e-08 1.19527883e-08 5.08483061e-08 1.19527881e-08
+ 5.09483061e-08 1.19527883e-08 5.1e-08 1.19527879e-08 5.101e-08 1.19388703e-08 5.103e-08 1.20206012e-08 5.107e-08 1.18457672e-08 5.115e-08 1.20757645e-08 5.125e-08 1.1824367e-08 5.135e-08 1.20762619e-08
+ 5.145e-08 1.18443259e-08 5.155e-08 1.2038956e-08 5.165e-08 1.18919423e-08 5.175e-08 1.19848996e-08 5.185e-08 1.19539955e-08 5.19308282e-08 1.24465481e-07 5.2e-08 1.72241691e-06 5.20086083e-08 -4.61584982e-06
+ 5.2025825e-08 -7.81178603e-06 5.20602584e-08 1.16927987e-06 5.21061808e-08 1.10985042e-05 5.21500808e-08 -1.1940293e-05 5.21980262e-08 9.09814381e-06 5.22553803e-08 -8.63968124e-06 5.23120186e-08 6.70517737e-06 5.24042316e-08 -4.84128351e-06
+ 5.25042316e-08 3.27353005e-06 5.26042316e-08 -1.93156633e-06 5.27042316e-08 9.66792548e-07 5.28042316e-08 -1.39411115e-07 5.29042316e-08 -5.11143768e-07 5.30042316e-08 1.11061772e-06 5.31042316e-08 -1.58512576e-06 5.32042316e-08 2.03140601e-06
+ 5.33042316e-08 -2.36567644e-06 5.34042316e-08 2.68328844e-06 5.35042316e-08 -2.89776465e-06 5.36042316e-08 3.1061765e-06 5.37042316e-08 -3.22064693e-06 5.38042316e-08 3.33976795e-06 5.39042316e-08 -3.37423912e-06 5.40042316e-08 3.42349279e-06
+ 5.41042316e-08 -3.39673646e-06 5.42042316e-08 3.39370537e-06 5.43042316e-08 -3.32218859e-06 5.44042316e-08 3.2818823e-06 5.45042316e-08 -3.17933511e-06 5.46042316e-08 3.11401264e-06 5.47042316e-08 -2.99144427e-06 5.48042316e-08 2.91077283e-06
+ 5.49042316e-08 -2.77673027e-06 5.50042316e-08 2.68810303e-06 5.51042316e-08 -2.54902948e-06 5.52042316e-08 2.45794128e-06 5.53042316e-08 -2.31855258e-06 5.54042316e-08 2.22895839e-06 5.55042316e-08 -2.09258845e-06 5.56042316e-08 2.00722724e-06
+ 5.57042316e-08 -1.87612843e-06 5.58042316e-08 1.79679708e-06 5.59042316e-08 -1.67239441e-06 5.60042316e-08 1.60017616e-06 5.61042316e-08 -1.48327258e-06 5.62042316e-08 1.41871919e-06 5.63042316e-08 -1.30965968e-06 5.64042316e-08 1.2529363e-06
+ 5.65042316e-08 -1.15173689e-06 5.66042316e-08 1.10273487e-06 5.67042316e-08 -1.00918253e-06 5.68042316e-08 9.67606175e-07 5.69042316e-08 -8.8133448e-07 5.70042316e-08 8.46766002e-07 5.71042316e-08 -7.67312428e-07 5.72042316e-08 7.39262185e-07
+ 5.73042316e-08 -6.661121e-07 5.74042316e-08 6.4405523e-07 5.75042316e-08 -5.7667259e-07 5.76042316e-08 5.60075112e-07 5.77042316e-08 -4.9792477e-07 5.78042316e-08 4.86261632e-07 5.79042316e-08 -4.28824054e-07 5.80042316e-08 4.21591092e-07
+ 5.81042316e-08 -3.68372207e-07 5.82042316e-08 3.65094039e-07 5.83042316e-08 -3.15631469e-07 5.84042316e-08 3.15866178e-07 5.85042316e-08 -2.69732673e-07 5.86042316e-08 2.73074123e-07 5.87042316e-08 -2.29878557e-07 5.88042316e-08 2.35955165e-07
+ 5.89042316e-08 -1.9533981e-07 5.90042316e-08 2.03814114e-07 5.91042316e-08 -1.65458182e-07 5.92042316e-08 1.76030701e-07 5.93042316e-08 -1.3965074e-07 5.94042316e-08 1.52056661e-07 5.95042316e-08 -1.1740137e-07 5.96042316e-08 1.31405583e-07
+ 5.97042316e-08 -9.82519779e-08 5.98042316e-08 1.13646203e-07 5.99042316e-08 -8.17971039e-08 6.00042316e-08 9.83974839e-08 6.01042316e-08 -6.76791171e-08 6.02042316e-08 8.53238762e-08 6.03042316e-08 -5.55835805e-08 6.04042316e-08 7.41319191e-08
+ 6.05042316e-08 -4.52380916e-08 6.06042316e-08 6.45672094e-08 6.07042316e-08 -3.64036965e-08 6.08042316e-08 5.64051731e-08 6.09042316e-08 -2.88693529e-08 6.10042316e-08 4.94482737e-08 6.11042316e-08 -2.24511338e-08 6.12042316e-08 4.35252522e-08
+ 6.13042316e-08 -1.69897409e-08 6.14042316e-08 3.84879328e-08 6.15042316e-08 -1.23474838e-08 6.16042316e-08 3.42083642e-08 6.17042316e-08 -8.40557957e-09 6.18042316e-08 3.05762537e-08 6.19042316e-08 -5.0617289e-09 6.20042316e-08 2.74967836e-08
+ 6.21042316e-08 -2.22816141e-09 6.22042316e-08 2.48886164e-08 6.23042316e-08 1.69359748e-10 6.24042316e-08 2.26840074e-08 6.25042316e-08 2.18276033e-09 6.26042316e-08 2.08449579e-08 6.27042316e-08 3.86219992e-09 6.28042316e-08 1.93116058e-08
+ 6.29042316e-08 5.2618627e-09 6.30042316e-08 1.80342611e-08 6.31042316e-08 6.42731685e-09 6.32042316e-08 1.6971138e-08 6.33042316e-08 7.39687012e-09 6.34042316e-08 1.60871281e-08 6.35042316e-08 8.20268908e-09 6.36042316e-08 1.53527666e-08
+ 6.37042316e-08 8.87175813e-09 6.38042316e-08 1.47433459e-08 6.39042316e-08 9.4266977e-09 6.40042316e-08 1.42382001e-08 6.41042316e-08 9.88639348e-09 6.42042316e-08 1.38200885e-08 6.43042316e-08 1.02662796e-08 6.44042316e-08 1.34749875e-08
+ 6.45042316e-08 1.0580019e-08 6.46042316e-08 1.31896313e-08 6.47042316e-08 1.0839496e-08 6.48042316e-08 1.29538844e-08 6.49042316e-08 1.10535145e-08 6.50042316e-08 1.27597098e-08 6.51042316e-08 1.12295803e-08 6.52042316e-08 1.26001551e-08
+ 6.53042316e-08 1.13740932e-08 6.54042316e-08 1.24693366e-08 6.55042316e-08 1.14924754e-08 6.56042316e-08 1.23621976e-08 6.57042316e-08 1.15894158e-08 6.58042316e-08 1.2274617e-08 6.59042316e-08 1.16683967e-08 6.60042316e-08 1.22034577e-08
+ 6.61042316e-08 1.17324807e-08 6.62042316e-08 1.21457766e-08 6.63042316e-08 1.17843603e-08 6.64042316e-08 1.20991589e-08 6.65042316e-08 1.18262081e-08 6.66042316e-08 1.20616316e-08 6.67042316e-08 1.18598228e-08 6.68042316e-08 1.20314808e-08
+ 6.69042316e-08 1.18868204e-08 6.70042316e-08 1.20075228e-08 6.71042316e-08 1.19080438e-08 6.72042316e-08 1.19886447e-08 6.73042316e-08 1.19248248e-08 6.74042316e-08 1.19737601e-08 6.75042316e-08 1.1937991e-08 6.76042316e-08 1.1962149e-08
+ 6.77042316e-08 1.19481968e-08 6.78042316e-08 1.19532121e-08 6.79042316e-08 1.19559915e-08 6.80042316e-08 1.19464441e-08 6.81042316e-08 1.1961838e-08 6.82042316e-08 1.19414231e-08 6.83042316e-08 1.19661196e-08 6.84042316e-08 1.19378023e-08
+ 6.85042316e-08 1.19691669e-08 6.86042316e-08 1.19352478e-08 6.87042316e-08 1.19712532e-08 6.88042316e-08 1.19336179e-08 6.89042316e-08 1.19724877e-08 6.90042316e-08 1.19327113e-08 6.91042316e-08 1.19731116e-08 6.92042316e-08 1.19323329e-08
+ 6.93042316e-08 1.1973279e-08 6.94042316e-08 1.1932347e-08 6.95042316e-08 1.19731015e-08 6.96042316e-08 1.19326725e-08 6.97042316e-08 1.19726475e-08 6.98042316e-08 1.1933235e-08 6.99042316e-08 1.19719942e-08 7.00042316e-08 1.1933964e-08
+ 7.01042316e-08 1.19712032e-08 7.02042316e-08 1.19348057e-08 7.03042316e-08 1.19703205e-08 7.04042316e-08 1.19357198e-08 7.05042316e-08 1.1969383e-08 7.06042316e-08 1.1936674e-08 7.07042316e-08 1.19684178e-08 7.08042316e-08 1.19376446e-08
+ 7.09042316e-08 1.19674471e-08 7.10042316e-08 1.1938612e-08 7.11042316e-08 1.19664863e-08 7.12042316e-08 1.19395623e-08 7.13042316e-08 1.19655489e-08 7.14042316e-08 1.19404847e-08 7.15042316e-08 1.19646433e-08 7.16042316e-08 1.19413727e-08
+ 7.17042316e-08 1.19637745e-08 7.18042316e-08 1.19422209e-08 7.19042316e-08 1.19629479e-08 7.20042316e-08 1.19430255e-08 7.21042316e-08 1.1962165e-08 7.22042316e-08 1.19437859e-08 7.23042316e-08 1.19614279e-08 7.24042316e-08 1.19445e-08
+ 7.25042316e-08 1.19607366e-08 7.26042316e-08 1.19451685e-08 7.27042316e-08 1.19600904e-08 7.28042316e-08 1.19457929e-08 7.29042316e-08 1.19594879e-08 7.30042316e-08 1.19463736e-08 7.31042316e-08 1.19589283e-08 7.32042316e-08 1.19469127e-08
+ 7.33042316e-08 1.19584095e-08 7.34042316e-08 1.19474114e-08 7.35042316e-08 1.19579301e-08 7.36042316e-08 1.19478723e-08 7.37042316e-08 1.19574874e-08 7.38042316e-08 1.19482969e-08 7.39042316e-08 1.19570805e-08 7.40042316e-08 1.19486868e-08
+ 7.41042316e-08 1.19567067e-08 7.42042316e-08 1.19490445e-08 7.43042316e-08 1.19563644e-08 7.44042316e-08 1.19493724e-08 7.45042316e-08 1.19560506e-08 7.46042316e-08 1.19496726e-08 7.47042316e-08 1.19557634e-08 7.48042316e-08 1.19499474e-08
+ 7.49042316e-08 1.19555006e-08 7.50042316e-08 1.19501984e-08 7.51042316e-08 1.19552605e-08 7.52042316e-08 1.19504281e-08 7.53042316e-08 1.19550413e-08 7.54042316e-08 1.19506375e-08 7.55042316e-08 1.19548413e-08 7.56042316e-08 1.19508289e-08
+ 7.57042316e-08 1.19546578e-08 7.58042316e-08 1.19510047e-08 7.59042316e-08 1.19544901e-08 7.60042316e-08 1.19511647e-08 7.61042316e-08 1.19543372e-08 7.62042316e-08 1.19513105e-08 7.63042316e-08 1.19541985e-08 7.64042316e-08 1.19514424e-08
+ 7.65042316e-08 1.1954073e-08 7.66042316e-08 1.19515624e-08 7.67042316e-08 1.19539583e-08 7.68042316e-08 1.19516716e-08 7.69042316e-08 1.1953854e-08 7.70042316e-08 1.19517711e-08 7.71042316e-08 1.19537592e-08 7.72042316e-08 1.19518616e-08
+ 7.73042316e-08 1.19536728e-08 7.74042316e-08 1.19519439e-08 7.75042316e-08 1.19535941e-08 7.76042316e-08 1.1952019e-08 7.77042316e-08 1.19535226e-08 7.78042316e-08 1.19520871e-08 7.79042316e-08 1.19534575e-08 7.80042316e-08 1.19521492e-08
+ 7.81042316e-08 1.19533984e-08 7.82042316e-08 1.19522061e-08 7.83042316e-08 1.19533443e-08 7.84042316e-08 1.19522572e-08 7.85042316e-08 1.19532949e-08 7.86042316e-08 1.19523046e-08 7.87042316e-08 1.19532503e-08 7.88042316e-08 1.19523474e-08
+ 7.89042316e-08 1.19532093e-08 7.90042316e-08 1.19523862e-08 7.91042316e-08 1.19531719e-08 7.92042316e-08 1.19524222e-08 7.93042316e-08 1.1953138e-08 7.94042316e-08 1.19524546e-08 7.95042316e-08 1.19531066e-08 7.96042316e-08 1.19524845e-08
+ 7.97042316e-08 1.19530784e-08 7.98042316e-08 1.19525117e-08 7.99042316e-08 1.19530523e-08 8.00042316e-08 1.19525363e-08 8.01042316e-08 1.19530289e-08 8.02042316e-08 1.19525587e-08 8.03042316e-08 1.19530073e-08 8.04042316e-08 1.19525793e-08
+ 8.05042316e-08 1.19529879e-08 8.06042316e-08 1.19525978e-08 8.07042316e-08 1.19529701e-08 8.08042316e-08 1.19526149e-08 8.09042316e-08 1.19529537e-08 8.10042316e-08 1.19526306e-08 8.11042316e-08 1.19529387e-08 8.12042316e-08 1.19526447e-08
+ 8.13042316e-08 1.1952925e-08 8.14042316e-08 1.19526581e-08 8.15042316e-08 1.19529127e-08 8.16042316e-08 1.19526694e-08 8.17042316e-08 1.19529014e-08 8.18042316e-08 1.19526803e-08 8.19042316e-08 1.19528913e-08 8.20042316e-08 1.19526901e-08
+ 8.21042316e-08 1.19528823e-08 8.22042316e-08 1.1952699e-08 8.23042316e-08 1.19528734e-08 8.24042316e-08 1.1952707e-08 8.25042316e-08 1.19528658e-08 8.26042316e-08 1.19527145e-08 8.27042316e-08 1.19528588e-08 8.28042316e-08 1.19527213e-08
+ 8.29042316e-08 1.19528522e-08 8.30042316e-08 1.19527276e-08 8.31042316e-08 1.19528461e-08 8.32042316e-08 1.19527331e-08 8.33042316e-08 1.19528411e-08 8.34042316e-08 1.19527383e-08 8.35042316e-08 1.19528363e-08 8.36042316e-08 1.19527428e-08
+ 8.37042316e-08 1.19528318e-08 8.38042316e-08 1.19527467e-08 8.39042316e-08 1.19528277e-08 8.40042316e-08 1.19527505e-08 8.41042316e-08 1.1952824e-08 8.42042316e-08 1.19527542e-08 8.43042316e-08 1.19528209e-08 8.44042316e-08 1.19527572e-08
+ 8.45042316e-08 1.19528179e-08 8.46042316e-08 1.19527603e-08 8.47042316e-08 1.19528151e-08 8.48042316e-08 1.19527624e-08 8.49042316e-08 1.19528127e-08 8.50042316e-08 1.1952765e-08 8.51042316e-08 1.19528105e-08 8.52042316e-08 1.1952767e-08
+ 8.53042316e-08 1.19528085e-08 8.54042316e-08 1.19527692e-08 8.55042316e-08 1.19528065e-08 8.56042316e-08 1.19527708e-08 8.57042316e-08 1.19528048e-08 8.58042316e-08 1.19527724e-08 8.59042316e-08 1.19528035e-08 8.60042316e-08 1.19527738e-08
+ 8.61042316e-08 1.19528018e-08 8.62042316e-08 1.19527753e-08 8.63042316e-08 1.19528007e-08 8.64042316e-08 1.19527764e-08 8.65042316e-08 1.19527997e-08 8.66042316e-08 1.19527774e-08 8.67042316e-08 1.19527987e-08 8.68042316e-08 1.19527784e-08
+ 8.69042316e-08 1.19527975e-08 8.70042316e-08 1.19527795e-08 8.71042316e-08 1.19527966e-08 8.72042316e-08 1.19527804e-08 8.73042316e-08 1.19527957e-08 8.74042316e-08 1.19527812e-08 8.75042316e-08 1.19527949e-08 8.76042316e-08 1.19527822e-08
+ 8.77042316e-08 1.19527942e-08 8.78042316e-08 1.19527826e-08 8.79042316e-08 1.19527936e-08 8.80042316e-08 1.1952783e-08 8.81042316e-08 1.19527932e-08 8.82042316e-08 1.19527835e-08 8.83042316e-08 1.19527928e-08 8.84042316e-08 1.19527841e-08
+ 8.85042316e-08 1.19527922e-08 8.86042316e-08 1.19527847e-08 8.87042316e-08 1.19527919e-08 8.88042316e-08 1.19527848e-08 8.89042316e-08 1.19527917e-08 8.90042316e-08 1.19527851e-08 8.91042316e-08 1.19527915e-08 8.92042316e-08 1.19527853e-08
+ 8.93042316e-08 1.19527911e-08 8.94042316e-08 1.19527857e-08 8.95042316e-08 1.1952791e-08 8.96042316e-08 1.19527858e-08 8.97042316e-08 1.19527909e-08 8.98042316e-08 1.1952786e-08 8.99042316e-08 1.19527904e-08 9.00042316e-08 1.19527864e-08
+ 9.01042316e-08 1.19527901e-08 9.02042316e-08 1.19527866e-08 9.03042316e-08 1.195279e-08 9.04042316e-08 1.19527867e-08 9.05042316e-08 1.19527899e-08 9.06042316e-08 1.1952787e-08 9.07042316e-08 1.19527895e-08 9.08042316e-08 1.19527871e-08
+ 9.09042316e-08 1.19527896e-08 9.10042316e-08 1.1952787e-08 9.11042316e-08 1.19527893e-08 9.12042316e-08 1.19527871e-08 9.13042316e-08 1.19527894e-08 9.14042316e-08 1.1952787e-08 9.15042316e-08 1.19527894e-08 9.16042316e-08 1.19527871e-08
+ 9.17042316e-08 1.19527894e-08 9.18042316e-08 1.19527872e-08 9.19042316e-08 1.19527895e-08 9.20042316e-08 1.19527873e-08 9.21042316e-08 1.1952789e-08 9.22042316e-08 1.19527876e-08 9.23042316e-08 1.19527891e-08 9.24042316e-08 1.19527877e-08
+ 9.25042316e-08 1.19527889e-08 9.26042316e-08 1.19527878e-08 9.27042316e-08 1.19527891e-08 9.28042316e-08 1.19527877e-08 9.29042316e-08 1.19527891e-08 9.30042316e-08 1.19527878e-08 9.31042316e-08 1.19527891e-08 9.32042316e-08 1.19527878e-08
+ 9.33042316e-08 1.1952789e-08 9.34042316e-08 1.19527876e-08 9.35042316e-08 1.19527889e-08 9.36042316e-08 1.19527877e-08 9.37042316e-08 1.19527891e-08 9.38042316e-08 1.19527877e-08 9.39042316e-08 1.19527891e-08 9.40042316e-08 1.19527878e-08
+ 9.41042316e-08 1.1952789e-08 9.42042316e-08 1.19527877e-08 9.43042316e-08 1.19527891e-08 9.44042316e-08 1.19527877e-08 9.45042316e-08 1.19527891e-08 9.46042316e-08 1.19527877e-08 9.47042316e-08 1.19527891e-08 9.48042316e-08 1.19527877e-08
+ 9.49042316e-08 1.19527891e-08 9.50042316e-08 1.19527878e-08 9.51042316e-08 1.19527891e-08 9.52042316e-08 1.19527878e-08 9.53042316e-08 1.19527887e-08 9.54042316e-08 1.19527877e-08 9.55042316e-08 1.19527886e-08 9.56042316e-08 1.1952788e-08
+ 9.57042316e-08 1.19527886e-08 9.58042316e-08 1.19527882e-08 9.59042316e-08 1.19527886e-08 9.60042316e-08 1.19527883e-08 9.61042316e-08 1.19527886e-08 9.62042316e-08 1.19527881e-08 9.63042316e-08 1.19527886e-08 9.64042316e-08 1.1952788e-08
+ 9.65042316e-08 1.19527884e-08 9.66042316e-08 1.19527878e-08 9.67042316e-08 1.19527885e-08 9.68042316e-08 1.19527882e-08 9.69042316e-08 1.19527882e-08 9.70042316e-08 1.1952788e-08 9.71042316e-08 1.19527883e-08 9.72042316e-08 1.1952788e-08
+ 9.73042316e-08 1.19527883e-08 9.74042316e-08 1.1952788e-08 9.75042316e-08 1.19527883e-08 9.76042316e-08 1.19527881e-08 9.77042316e-08 1.19527883e-08 9.78042316e-08 1.19527881e-08 9.79042316e-08 1.19527883e-08 9.80042316e-08 1.1952788e-08
+ 9.81042316e-08 1.19527883e-08 9.82042316e-08 1.1952788e-08 9.83042316e-08 1.19527883e-08 9.84042316e-08 1.19527881e-08 9.85042316e-08 1.19527884e-08 9.86042316e-08 1.1952788e-08 9.87042316e-08 1.19527883e-08 9.88042316e-08 1.19527879e-08
+ 9.89042316e-08 1.19527883e-08 9.90042316e-08 1.1952788e-08 9.91042316e-08 1.19527883e-08 9.92042316e-08 1.1952788e-08 9.93042316e-08 1.19527883e-08 9.94042316e-08 1.1952788e-08 9.95042316e-08 1.19527883e-08 9.96042316e-08 1.19527879e-08
+ 9.97042316e-08 1.19527883e-08 9.98042316e-08 1.1952788e-08 9.99042316e-08 1.19527882e-08 1e-07 1.19527883e-08 1.0001e-07 1.19892439e-08 1.0003e-07 1.17769501e-08 1.0007e-07 1.22259536e-08 1.0015e-07 1.16459511e-08
+ 1.0025e-07 1.22666862e-08 1.0035e-07 1.16511428e-08 1.0045e-07 1.22243693e-08 1.0055e-07 1.17333459e-08 1.0065e-07 1.18158097e-08 1.0075e-07 2.88746968e-08 1.0085e-07 -5.4466577e-07 1.00932051e-07 7.37611719e-06
+ 1.01e-07 -4.67556033e-05 1.01008488e-07 -5.14147198e-05 1.01025463e-07 -3.72261328e-05 1.01059414e-07 -3.09370444e-05 1.0109062e-07 0.000250558184 1.0114347e-07 0.000494689166 1.01199151e-07 0.00157105355 1.01299151e-07 -0.0175443595
+ 1.01399151e-07 0.171698395 1.01499151e-07 4.36413971 1.01599151e-07 5.20247686 1.01699151e-07 4.88242009 1.01799151e-07 5.06727389 1.01893117e-07 4.95839538 1.01993117e-07 5.02693002 1.02093117e-07 4.98190659
+ 1.02193117e-07 5.012155 1.02293117e-07 4.99169062 1.02393117e-07 5.00564782 1.02493117e-07 4.9961172 1.02593117e-07 5.00264947 1.02693117e-07 4.99817488 1.02793117e-07 5.00124726 1.02893117e-07 4.99914008
+ 1.02993117e-07 5.00058802 1.03093117e-07 4.99959444 1.03193117e-07 5.00027735 1.03293117e-07 4.99980871 1.03393117e-07 5.00013073 1.03493117e-07 4.99990988 1.03593117e-07 5.00006148 1.03693117e-07 4.99995768
+ 1.03793117e-07 5.00002877 1.03893117e-07 4.99998025 1.03993117e-07 5.00001332 1.04093117e-07 4.9999909 1.04193117e-07 5.00000605 1.04293117e-07 4.99999589 1.04393117e-07 5.00000265 1.04493117e-07 4.99999822
+ 1.04593117e-07 5.00000108 1.04693117e-07 4.99999928 1.04793117e-07 5.00000037 1.04893117e-07 4.99999976 1.04993117e-07 5.00000007 1.05093117e-07 4.99999995 1.05193117e-07 4.99999995 1.05293117e-07 5.00000002
+ 1.05393117e-07 4.99999991 1.05493117e-07 5.00000004 1.05593117e-07 4.99999991 1.05693117e-07 5.00000003 1.05793117e-07 4.99999992 1.05893117e-07 5.00000002 1.05993117e-07 4.99999993 1.06093117e-07 5.0
+ 1.06193117e-07 4.99999995 1.06293117e-07 4.99999999 1.06393117e-07 4.99999996 1.06493117e-07 4.99999998 1.06593117e-07 4.99999997 1.06693117e-07 4.99999997 1.06793117e-07 4.99999997 1.06893117e-07 4.99999997
+ 1.06993117e-07 4.99999998 1.07093117e-07 4.99999997 1.07193117e-07 4.99999998 1.07293117e-07 4.99999996 1.07393117e-07 4.99999998 1.07493117e-07 4.99999996 1.07593117e-07 4.99999998 1.07693117e-07 4.99999996
+ 1.07793117e-07 4.99999998 1.07893117e-07 4.99999996 1.07993117e-07 4.99999998 1.08093117e-07 4.99999996 1.08193117e-07 4.99999998 1.08293117e-07 4.99999996 1.08393117e-07 4.99999998 1.08493117e-07 4.99999996
+ 1.08593117e-07 4.99999998 1.08693117e-07 4.99999996 1.08793117e-07 4.99999998 1.08893117e-07 4.99999996 1.08993117e-07 4.99999998 1.09093117e-07 4.99999996 1.09193117e-07 4.99999998 1.09293117e-07 4.99999997
+ 1.09393117e-07 4.99999998 1.09493117e-07 4.99999997 1.09593117e-07 4.99999998 1.09693117e-07 4.99999997 1.09793117e-07 4.99999998 1.09893117e-07 4.99999997 1.09993117e-07 4.99999998 1.10093117e-07 4.99999997
+ 1.10193117e-07 4.99999998 1.10293117e-07 4.99999997 1.10393117e-07 4.99999998 1.10493117e-07 4.99999997 1.10593117e-07 4.99999998 1.10693117e-07 4.99999997 1.10793117e-07 4.99999998 1.10893117e-07 4.99999997
+ 1.10993117e-07 4.99999997 1.11093117e-07 4.99999997 1.11193117e-07 4.99999997 1.11293117e-07 4.99999997 1.11393117e-07 4.99999997 1.11493117e-07 4.99999997 1.11593117e-07 4.99999997 1.11693117e-07 4.99999997
+ 1.11793117e-07 4.99999997 1.11893117e-07 4.99999997 1.11993117e-07 4.99999997 1.12093117e-07 4.99999997 1.12193117e-07 4.99999997 1.12293117e-07 4.99999997 1.12393117e-07 4.99999997 1.12493117e-07 4.99999997
+ 1.12593117e-07 4.99999997 1.12693117e-07 4.99999997 1.12793117e-07 4.99999997 1.12893117e-07 4.99999997 1.12993117e-07 4.99999997 1.13093117e-07 4.99999997 1.13193117e-07 4.99999997 1.13293117e-07 4.99999997
+ 1.13393117e-07 4.99999997 1.13493117e-07 4.99999997 1.13593117e-07 4.99999997 1.13693117e-07 4.99999997 1.13793117e-07 4.99999997 1.13893117e-07 4.99999997 1.13993117e-07 4.99999997 1.14093117e-07 4.99999997
+ 1.14193117e-07 4.99999997 1.14293117e-07 4.99999997 1.14393117e-07 4.99999997 1.14493117e-07 4.99999997 1.14593117e-07 4.99999997 1.14693117e-07 4.99999997 1.14793117e-07 4.99999997 1.14893117e-07 4.99999997
+ 1.14993117e-07 4.99999997 1.15093117e-07 4.99999997 1.15193117e-07 4.99999997 1.15293117e-07 4.99999997 1.15393117e-07 4.99999997 1.15493117e-07 4.99999997 1.15593117e-07 4.99999997 1.15693117e-07 4.99999997
+ 1.15793117e-07 4.99999997 1.15893117e-07 4.99999997 1.15993117e-07 4.99999997 1.16093117e-07 4.99999997 1.16193117e-07 4.99999997 1.16293117e-07 4.99999997 1.16393117e-07 4.99999997 1.16493117e-07 4.99999997
+ 1.16593117e-07 4.99999997 1.16693117e-07 4.99999997 1.16793117e-07 4.99999997 1.16893117e-07 4.99999997 1.16993117e-07 4.99999997 1.17093117e-07 4.99999997 1.17193117e-07 4.99999997 1.17293117e-07 4.99999997
+ 1.17393117e-07 4.99999997 1.17493117e-07 4.99999997 1.17593117e-07 4.99999997 1.17693117e-07 4.99999997 1.17793117e-07 4.99999997 1.17893117e-07 4.99999997 1.17993117e-07 4.99999997 1.18093117e-07 4.99999997
+ 1.18193117e-07 4.99999997 1.18293117e-07 4.99999997 1.18393117e-07 4.99999997 1.18493117e-07 4.99999997 1.18593117e-07 4.99999997 1.18693117e-07 4.99999997 1.18793117e-07 4.99999997 1.18893117e-07 4.99999997
+ 1.18993117e-07 4.99999997 1.19093117e-07 4.99999997 1.19193117e-07 4.99999997 1.19293117e-07 4.99999997 1.19393117e-07 4.99999997 1.19493117e-07 4.99999997 1.19593117e-07 4.99999997 1.19693117e-07 4.99999997
+ 1.19793117e-07 4.99999997 1.19893117e-07 4.99999997 1.19993117e-07 4.99999997 1.20093117e-07 4.99999997 1.20193117e-07 4.99999997 1.20293117e-07 4.99999997 1.20393117e-07 4.99999997 1.20493117e-07 4.99999997
+ 1.20593117e-07 4.99999997 1.20693117e-07 4.99999997 1.20793117e-07 4.99999997 1.20893117e-07 4.99999997 1.20993117e-07 4.99999997 1.21093117e-07 4.99999997 1.21193117e-07 4.99999997 1.21293117e-07 4.99999997
+ 1.21393117e-07 4.99999997 1.21493117e-07 4.99999997 1.21593117e-07 4.99999997 1.21693117e-07 4.99999997 1.21793117e-07 4.99999997 1.21893117e-07 4.99999997 1.21993117e-07 4.99999997 1.22093117e-07 4.99999997
+ 1.22193117e-07 4.99999997 1.22293117e-07 4.99999997 1.22393117e-07 4.99999997 1.22493117e-07 4.99999997 1.22593117e-07 4.99999997 1.22693117e-07 4.99999997 1.22793117e-07 4.99999997 1.22893117e-07 4.99999997
+ 1.22993117e-07 4.99999997 1.23093117e-07 4.99999997 1.23193117e-07 4.99999997 1.23293117e-07 4.99999997 1.23393117e-07 4.99999997 1.23493117e-07 4.99999997 1.23593117e-07 4.99999997 1.23693117e-07 4.99999997
+ 1.23793117e-07 4.99999997 1.23893117e-07 4.99999997 1.23993117e-07 4.99999997 1.24093117e-07 4.99999997 1.24193117e-07 4.99999997 1.24293117e-07 4.99999997 1.24393117e-07 4.99999997 1.24493117e-07 4.99999997
+ 1.24593117e-07 4.99999997 1.24693117e-07 4.99999997 1.24793117e-07 4.99999997 1.24893117e-07 4.99999997 1.24993117e-07 4.99999997 1.25093117e-07 4.99999997 1.25193117e-07 4.99999997 1.25293117e-07 4.99999997
+ 1.25393117e-07 4.99999997 1.25493117e-07 4.99999997 1.25593117e-07 4.99999997 1.25693117e-07 4.99999997 1.25793117e-07 4.99999997 1.25893117e-07 4.99999997 1.25993117e-07 4.99999997 1.26093117e-07 4.99999997
+ 1.26193117e-07 4.99999997 1.26293117e-07 4.99999997 1.26393117e-07 4.99999997 1.26493117e-07 4.99999997 1.26593117e-07 4.99999997 1.26693117e-07 4.99999997 1.26793117e-07 4.99999997 1.26893117e-07 4.99999997
+ 1.26993117e-07 4.99999997 1.27093117e-07 4.99999997 1.27193117e-07 4.99999997 1.27293117e-07 4.99999997 1.27393117e-07 4.99999997 1.27493117e-07 4.99999997 1.27593117e-07 4.99999997 1.27693117e-07 4.99999997
+ 1.27793117e-07 4.99999997 1.27893117e-07 4.99999997 1.27993117e-07 4.99999997 1.28093117e-07 4.99999997 1.28193117e-07 4.99999997 1.28293117e-07 4.99999997 1.28393117e-07 4.99999997 1.28493117e-07 4.99999997
+ 1.28593117e-07 4.99999997 1.28693117e-07 4.99999997 1.28793117e-07 4.99999997 1.28893117e-07 4.99999997 1.28993117e-07 4.99999997 1.29093117e-07 4.99999997 1.29193117e-07 4.99999997 1.29293117e-07 4.99999997
+ 1.29393117e-07 4.99999997 1.29493117e-07 4.99999997 1.29593117e-07 4.99999997 1.29693117e-07 4.99999997 1.29793117e-07 4.99999997 1.29893117e-07 4.99999997 1.29993117e-07 4.99999997 1.30093117e-07 4.99999997
+ 1.30193117e-07 4.99999997 1.30293117e-07 4.99999997 1.30393117e-07 4.99999997 1.30493117e-07 4.99999997 1.30593117e-07 4.99999997 1.30693117e-07 4.99999997 1.30793117e-07 4.99999997 1.30893117e-07 4.99999997
+ 1.30993117e-07 4.99999997 1.31093117e-07 4.99999997 1.31193117e-07 4.99999997 1.31293117e-07 4.99999997 1.31393117e-07 4.99999997 1.31493117e-07 4.99999997 1.31593117e-07 4.99999997 1.31693117e-07 4.99999997
+ 1.31793117e-07 4.99999997 1.31893117e-07 4.99999997 1.31993117e-07 4.99999997 1.32093117e-07 4.99999997 1.32193117e-07 4.99999997 1.32293117e-07 4.99999997 1.32393117e-07 4.99999997 1.32493117e-07 4.99999997
+ 1.32593117e-07 4.99999997 1.32693117e-07 4.99999997 1.32793117e-07 4.99999997 1.32893117e-07 4.99999997 1.32993117e-07 4.99999997 1.33093117e-07 4.99999997 1.33193117e-07 4.99999997 1.33293117e-07 4.99999997
+ 1.33393117e-07 4.99999997 1.33493117e-07 4.99999997 1.33593117e-07 4.99999997 1.33693117e-07 4.99999997 1.33793117e-07 4.99999997 1.33893117e-07 4.99999997 1.33993117e-07 4.99999997 1.34093117e-07 4.99999997
+ 1.34193117e-07 4.99999997 1.34293117e-07 4.99999997 1.34393117e-07 4.99999997 1.34493117e-07 4.99999997 1.34593117e-07 4.99999997 1.34693117e-07 4.99999997 1.34793117e-07 4.99999997 1.34893117e-07 4.99999997
+ 1.34993117e-07 4.99999997 1.35093117e-07 4.99999997 1.35193117e-07 4.99999997 1.35293117e-07 4.99999997 1.35393117e-07 4.99999997 1.35493117e-07 4.99999997 1.35593117e-07 4.99999997 1.35693117e-07 4.99999997
+ 1.35793117e-07 4.99999997 1.35893117e-07 4.99999997 1.35993117e-07 4.99999997 1.36093117e-07 4.99999997 1.36193117e-07 4.99999997 1.36293117e-07 4.99999997 1.36393117e-07 4.99999997 1.36493117e-07 4.99999997
+ 1.36593117e-07 4.99999997 1.36693117e-07 4.99999997 1.36793117e-07 4.99999997 1.36893117e-07 4.99999997 1.36993117e-07 4.99999997 1.37093117e-07 4.99999997 1.37193117e-07 4.99999997 1.37293117e-07 4.99999997
+ 1.37393117e-07 4.99999997 1.37493117e-07 4.99999997 1.37593117e-07 4.99999997 1.37693117e-07 4.99999997 1.37793117e-07 4.99999997 1.37893117e-07 4.99999997 1.37993117e-07 4.99999997 1.38093117e-07 4.99999997
+ 1.38193117e-07 4.99999997 1.38293117e-07 4.99999997 1.38393117e-07 4.99999997 1.38493117e-07 4.99999997 1.38593117e-07 4.99999997 1.38693117e-07 4.99999997 1.38793117e-07 4.99999997 1.38893117e-07 4.99999997
+ 1.38993117e-07 4.99999997 1.39093117e-07 4.99999997 1.39193117e-07 4.99999997 1.39293117e-07 4.99999997 1.39393117e-07 4.99999997 1.39493117e-07 4.99999997 1.39593117e-07 4.99999997 1.39693117e-07 4.99999997
+ 1.39793117e-07 4.99999997 1.39893117e-07 4.99999997 1.39993117e-07 4.99999997 1.40093117e-07 4.99999997 1.40193117e-07 4.99999997 1.40293117e-07 4.99999997 1.40393117e-07 4.99999997 1.40493117e-07 4.99999997
+ 1.40593117e-07 4.99999997 1.40693117e-07 4.99999997 1.40793117e-07 4.99999997 1.40893117e-07 4.99999997 1.40993117e-07 4.99999997 1.41093117e-07 4.99999997 1.41193117e-07 4.99999997 1.41293117e-07 4.99999997
+ 1.41393117e-07 4.99999997 1.41493117e-07 4.99999997 1.41593117e-07 4.99999997 1.41693117e-07 4.99999997 1.41793117e-07 4.99999997 1.41893117e-07 4.99999997 1.41993117e-07 4.99999997 1.42093117e-07 4.99999997
+ 1.42193117e-07 4.99999997 1.42293117e-07 4.99999997 1.42393117e-07 4.99999997 1.42493117e-07 4.99999997 1.42593117e-07 4.99999997 1.42693117e-07 4.99999997 1.42793117e-07 4.99999997 1.42893117e-07 4.99999997
+ 1.42993117e-07 4.99999997 1.43093117e-07 4.99999997 1.43193117e-07 4.99999997 1.43293117e-07 4.99999997 1.43393117e-07 4.99999997 1.43493117e-07 4.99999997 1.43593117e-07 4.99999997 1.43693117e-07 4.99999997
+ 1.43793117e-07 4.99999997 1.43893117e-07 4.99999997 1.43993117e-07 4.99999997 1.44093117e-07 4.99999997 1.44193117e-07 4.99999997 1.44293117e-07 4.99999997 1.44393117e-07 4.99999997 1.44493117e-07 4.99999997
+ 1.44593117e-07 4.99999997 1.44693117e-07 4.99999997 1.44793117e-07 4.99999997 1.44893117e-07 4.99999997 1.44993117e-07 4.99999997 1.45093117e-07 4.99999997 1.45193117e-07 4.99999997 1.45293117e-07 4.99999997
+ 1.45393117e-07 4.99999997 1.45493117e-07 4.99999997 1.45593117e-07 4.99999997 1.45693117e-07 4.99999997 1.45793117e-07 4.99999997 1.45893117e-07 4.99999997 1.45993117e-07 4.99999997 1.46093117e-07 4.99999997
+ 1.46193117e-07 4.99999997 1.46293117e-07 4.99999997 1.46393117e-07 4.99999997 1.46493117e-07 4.99999997 1.46593117e-07 4.99999997 1.46693117e-07 4.99999997 1.46793117e-07 4.99999997 1.46893117e-07 4.99999997
+ 1.46993117e-07 4.99999997 1.47093117e-07 4.99999997 1.47193117e-07 4.99999997 1.47293117e-07 4.99999997 1.47393117e-07 4.99999997 1.47493117e-07 4.99999997 1.47593117e-07 4.99999997 1.47693117e-07 4.99999997
+ 1.47793117e-07 4.99999997 1.47893117e-07 4.99999997 1.47993117e-07 4.99999997 1.48093117e-07 4.99999997 1.48193117e-07 4.99999997 1.48293117e-07 4.99999997 1.48393117e-07 4.99999997 1.48493117e-07 4.99999997
+ 1.48593117e-07 4.99999997 1.48693117e-07 4.99999997 1.48793117e-07 4.99999997 1.48893117e-07 4.99999997 1.48993117e-07 4.99999997 1.49093117e-07 4.99999997 1.49193117e-07 4.99999997 1.49293117e-07 4.99999997
+ 1.49393117e-07 4.99999997 1.49493117e-07 4.99999997 1.49593117e-07 4.99999997 1.49693117e-07 4.99999997 1.49793117e-07 4.99999997 1.49893117e-07 4.99999997 1.49993117e-07 4.99999997 1.50093117e-07 4.99999997
+ 1.50193117e-07 4.99999997 1.50293117e-07 4.99999997 1.50393117e-07 4.99999997 1.50493117e-07 4.99999997 1.50593117e-07 4.99999997 1.50693117e-07 4.99999997 1.50793117e-07 4.99999997 1.50893117e-07 4.99999997
+ 1.50993117e-07 4.99999997 1.51e-07 4.99999997 1.5101e-07 4.99999997 1.5103e-07 4.99999997 1.5107e-07 4.99999997 1.5115e-07 4.99999997 1.5125e-07 4.99999997 1.5135e-07 4.99999997
+ 1.5145e-07 4.99999997 1.5155e-07 4.99999997 1.5165e-07 4.99999997 1.5175e-07 4.99999997 1.5185e-07 4.99999997 1.51930828e-07 5.00000065 1.52e-07 5.00000149 1.52008608e-07 4.99999288
+ 1.52025825e-07 4.99997549 1.52060258e-07 4.99999257 1.52106188e-07 5.00004375 1.52150118e-07 5.00000856 1.5219811e-07 4.99994581 1.52255501e-07 5.00002983 1.52312176e-07 4.99999321 1.52404431e-07 5.00000355
+ 1.52490774e-07 5.00000011 1.52590774e-07 4.99999756 1.52690774e-07 5.00000329 1.52790774e-07 4.99999639 1.52890774e-07 5.0000034 1.52990774e-07 4.99999687 1.53090774e-07 5.00000266 1.53190774e-07 4.9999977
+ 1.53290774e-07 5.00000186 1.53390774e-07 4.99999842 1.53490774e-07 5.00000123 1.53590774e-07 4.99999895 1.53690774e-07 5.00000079 1.53790774e-07 4.99999931 1.53890774e-07 5.00000051 1.53990774e-07 4.99999954
+ 1.54090774e-07 5.00000033 1.54190774e-07 4.99999968 1.54290774e-07 5.00000021 1.54390774e-07 4.99999977 1.54490774e-07 5.00000014 1.54590774e-07 4.99999983 1.54690774e-07 5.00000009 1.54790774e-07 4.99999987
+ 1.54890774e-07 5.00000007 1.54990774e-07 4.99999989 1.55090774e-07 5.00000005 1.55190774e-07 4.99999991 1.55290774e-07 5.00000003 1.55390774e-07 4.99999992 1.55490774e-07 5.00000002 1.55590774e-07 4.99999993
+ 1.55690774e-07 5.00000001 1.55790774e-07 4.99999993 1.55890774e-07 5.00000001 1.55990774e-07 4.99999994 1.56090774e-07 5.0 1.56190774e-07 4.99999994 1.56290774e-07 5.0 1.56390774e-07 4.99999995
+ 1.56490774e-07 5.0 1.56590774e-07 4.99999995 1.56690774e-07 4.99999999 1.56790774e-07 4.99999995 1.56890774e-07 4.99999999 1.56990774e-07 4.99999996 1.57090774e-07 4.99999999 1.57190774e-07 4.99999996
+ 1.57290774e-07 4.99999999 1.57390774e-07 4.99999996 1.57490774e-07 4.99999998 1.57590774e-07 4.99999996 1.57690774e-07 4.99999998 1.57790774e-07 4.99999996 1.57890774e-07 4.99999998 1.57990774e-07 4.99999996
+ 1.58090774e-07 4.99999998 1.58190774e-07 4.99999997 1.58290774e-07 4.99999998 1.58390774e-07 4.99999997 1.58490774e-07 4.99999998 1.58590774e-07 4.99999997 1.58690774e-07 4.99999998 1.58790774e-07 4.99999997
+ 1.58890774e-07 4.99999998 1.58990774e-07 4.99999997 1.59090774e-07 4.99999998 1.59190774e-07 4.99999997 1.59290774e-07 4.99999997 1.59390774e-07 4.99999997 1.59490774e-07 4.99999997 1.59590774e-07 4.99999997
+ 1.59690774e-07 4.99999997 1.59790774e-07 4.99999997 1.59890774e-07 4.99999997 1.59990774e-07 4.99999997 1.60090774e-07 4.99999997 1.60190774e-07 4.99999997 1.60290774e-07 4.99999997 1.60390774e-07 4.99999997
+ 1.60490774e-07 4.99999997 1.60590774e-07 4.99999997 1.60690774e-07 4.99999997 1.60790774e-07 4.99999997 1.60890774e-07 4.99999997 1.60990774e-07 4.99999997 1.61090774e-07 4.99999997 1.61190774e-07 4.99999997
+ 1.61290774e-07 4.99999997 1.61390774e-07 4.99999997 1.61490774e-07 4.99999997 1.61590774e-07 4.99999997 1.61690774e-07 4.99999997 1.61790774e-07 4.99999997 1.61890774e-07 4.99999997 1.61990774e-07 4.99999997
+ 1.62090774e-07 4.99999997 1.62190774e-07 4.99999997 1.62290774e-07 4.99999997 1.62390774e-07 4.99999997 1.62490774e-07 4.99999997 1.62590774e-07 4.99999997 1.62690774e-07 4.99999997 1.62790774e-07 4.99999997
+ 1.62890774e-07 4.99999997 1.62990774e-07 4.99999997 1.63090774e-07 4.99999997 1.63190774e-07 4.99999997 1.63290774e-07 4.99999997 1.63390774e-07 4.99999997 1.63490774e-07 4.99999997 1.63590774e-07 4.99999997
+ 1.63690774e-07 4.99999997 1.63790774e-07 4.99999997 1.63890774e-07 4.99999997 1.63990774e-07 4.99999997 1.64090774e-07 4.99999997 1.64190774e-07 4.99999997 1.64290774e-07 4.99999997 1.64390774e-07 4.99999997
+ 1.64490774e-07 4.99999997 1.64590774e-07 4.99999997 1.64690774e-07 4.99999997 1.64790774e-07 4.99999997 1.64890774e-07 4.99999997 1.64990774e-07 4.99999997 1.65090774e-07 4.99999997 1.65190774e-07 4.99999997
+ 1.65290774e-07 4.99999997 1.65390774e-07 4.99999997 1.65490774e-07 4.99999997 1.65590774e-07 4.99999997 1.65690774e-07 4.99999997 1.65790774e-07 4.99999997 1.65890774e-07 4.99999997 1.65990774e-07 4.99999997
+ 1.66090774e-07 4.99999997 1.66190774e-07 4.99999997 1.66290774e-07 4.99999997 1.66390774e-07 4.99999997 1.66490774e-07 4.99999997 1.66590774e-07 4.99999997 1.66690774e-07 4.99999997 1.66790774e-07 4.99999997
+ 1.66890774e-07 4.99999997 1.66990774e-07 4.99999997 1.67090774e-07 4.99999997 1.67190774e-07 4.99999997 1.67290774e-07 4.99999997 1.67390774e-07 4.99999997 1.67490774e-07 4.99999997 1.67590774e-07 4.99999997
+ 1.67690774e-07 4.99999997 1.67790774e-07 4.99999997 1.67890774e-07 4.99999997 1.67990774e-07 4.99999997 1.68090774e-07 4.99999997 1.68190774e-07 4.99999997 1.68290774e-07 4.99999997 1.68390774e-07 4.99999997
+ 1.68490774e-07 4.99999997 1.68590774e-07 4.99999997 1.68690774e-07 4.99999997 1.68790774e-07 4.99999997 1.68890774e-07 4.99999997 1.68990774e-07 4.99999997 1.69090774e-07 4.99999997 1.69190774e-07 4.99999997
+ 1.69290774e-07 4.99999997 1.69390774e-07 4.99999997 1.69490774e-07 4.99999997 1.69590774e-07 4.99999997 1.69690774e-07 4.99999997 1.69790774e-07 4.99999997 1.69890774e-07 4.99999997 1.69990774e-07 4.99999997
+ 1.70090774e-07 4.99999997 1.70190774e-07 4.99999997 1.70290774e-07 4.99999997 1.70390774e-07 4.99999997 1.70490774e-07 4.99999997 1.70590774e-07 4.99999997 1.70690774e-07 4.99999997 1.70790774e-07 4.99999997
+ 1.70890774e-07 4.99999997 1.70990774e-07 4.99999997 1.71090774e-07 4.99999997 1.71190774e-07 4.99999997 1.71290774e-07 4.99999997 1.71390774e-07 4.99999997 1.71490774e-07 4.99999997 1.71590774e-07 4.99999997
+ 1.71690774e-07 4.99999997 1.71790774e-07 4.99999997 1.71890774e-07 4.99999997 1.71990774e-07 4.99999997 1.72090774e-07 4.99999997 1.72190774e-07 4.99999997 1.72290774e-07 4.99999997 1.72390774e-07 4.99999997
+ 1.72490774e-07 4.99999997 1.72590774e-07 4.99999997 1.72690774e-07 4.99999997 1.72790774e-07 4.99999997 1.72890774e-07 4.99999997 1.72990774e-07 4.99999997 1.73090774e-07 4.99999997 1.73190774e-07 4.99999997
+ 1.73290774e-07 4.99999997 1.73390774e-07 4.99999997 1.73490774e-07 4.99999997 1.73590774e-07 4.99999997 1.73690774e-07 4.99999997 1.73790774e-07 4.99999997 1.73890774e-07 4.99999997 1.73990774e-07 4.99999997
+ 1.74090774e-07 4.99999997 1.74190774e-07 4.99999997 1.74290774e-07 4.99999997 1.74390774e-07 4.99999997 1.74490774e-07 4.99999997 1.74590774e-07 4.99999997 1.74690774e-07 4.99999997 1.74790774e-07 4.99999997
+ 1.74890774e-07 4.99999997 1.74990774e-07 4.99999997 1.75090774e-07 4.99999997 1.75190774e-07 4.99999997 1.75290774e-07 4.99999997 1.75390774e-07 4.99999997 1.75490774e-07 4.99999997 1.75590774e-07 4.99999997
+ 1.75690774e-07 4.99999997 1.75790774e-07 4.99999997 1.75890774e-07 4.99999997 1.75990774e-07 4.99999997 1.76090774e-07 4.99999997 1.76190774e-07 4.99999997 1.76290774e-07 4.99999997 1.76390774e-07 4.99999997
+ 1.76490774e-07 4.99999997 1.76590774e-07 4.99999997 1.76690774e-07 4.99999997 1.76790774e-07 4.99999997 1.76890774e-07 4.99999997 1.76990774e-07 4.99999997 1.77090774e-07 4.99999997 1.77190774e-07 4.99999997
+ 1.77290774e-07 4.99999997 1.77390774e-07 4.99999997 1.77490774e-07 4.99999997 1.77590774e-07 4.99999997 1.77690774e-07 4.99999997 1.77790774e-07 4.99999997 1.77890774e-07 4.99999997 1.77990774e-07 4.99999997
+ 1.78090774e-07 4.99999997 1.78190774e-07 4.99999997 1.78290774e-07 4.99999997 1.78390774e-07 4.99999997 1.78490774e-07 4.99999997 1.78590774e-07 4.99999997 1.78690774e-07 4.99999997 1.78790774e-07 4.99999997
+ 1.78890774e-07 4.99999997 1.78990774e-07 4.99999997 1.79090774e-07 4.99999997 1.79190774e-07 4.99999997 1.79290774e-07 4.99999997 1.79390774e-07 4.99999997 1.79490774e-07 4.99999997 1.79590774e-07 4.99999997
+ 1.79690774e-07 4.99999997 1.79790774e-07 4.99999997 1.79890774e-07 4.99999997 1.79990774e-07 4.99999997 1.80090774e-07 4.99999997 1.80190774e-07 4.99999997 1.80290774e-07 4.99999997 1.80390774e-07 4.99999997
+ 1.80490774e-07 4.99999997 1.80590774e-07 4.99999997 1.80690774e-07 4.99999997 1.80790774e-07 4.99999997 1.80890774e-07 4.99999997 1.80990774e-07 4.99999997 1.81090774e-07 4.99999997 1.81190774e-07 4.99999997
+ 1.81290774e-07 4.99999997 1.81390774e-07 4.99999997 1.81490774e-07 4.99999997 1.81590774e-07 4.99999997 1.81690774e-07 4.99999997 1.81790774e-07 4.99999997 1.81890774e-07 4.99999997 1.81990774e-07 4.99999997
+ 1.82090774e-07 4.99999997 1.82190774e-07 4.99999997 1.82290774e-07 4.99999997 1.82390774e-07 4.99999997 1.82490774e-07 4.99999997 1.82590774e-07 4.99999997 1.82690774e-07 4.99999997 1.82790774e-07 4.99999997
+ 1.82890774e-07 4.99999997 1.82990774e-07 4.99999997 1.83090774e-07 4.99999997 1.83190774e-07 4.99999997 1.83290774e-07 4.99999997 1.83390774e-07 4.99999997 1.83490774e-07 4.99999997 1.83590774e-07 4.99999997
+ 1.83690774e-07 4.99999997 1.83790774e-07 4.99999997 1.83890774e-07 4.99999997 1.83990774e-07 4.99999997 1.84090774e-07 4.99999997 1.84190774e-07 4.99999997 1.84290774e-07 4.99999997 1.84390774e-07 4.99999997
+ 1.84490774e-07 4.99999997 1.84590774e-07 4.99999997 1.84690774e-07 4.99999997 1.84790774e-07 4.99999997 1.84890774e-07 4.99999997 1.84990774e-07 4.99999997 1.85090774e-07 4.99999997 1.85190774e-07 4.99999997
+ 1.85290774e-07 4.99999997 1.85390774e-07 4.99999997 1.85490774e-07 4.99999997 1.85590774e-07 4.99999997 1.85690774e-07 4.99999997 1.85790774e-07 4.99999997 1.85890774e-07 4.99999997 1.85990774e-07 4.99999997
+ 1.86090774e-07 4.99999997 1.86190774e-07 4.99999997 1.86290774e-07 4.99999997 1.86390774e-07 4.99999997 1.86490774e-07 4.99999997 1.86590774e-07 4.99999997 1.86690774e-07 4.99999997 1.86790774e-07 4.99999997
+ 1.86890774e-07 4.99999997 1.86990774e-07 4.99999997 1.87090774e-07 4.99999997 1.87190774e-07 4.99999997 1.87290774e-07 4.99999997 1.87390774e-07 4.99999997 1.87490774e-07 4.99999997 1.87590774e-07 4.99999997
+ 1.87690774e-07 4.99999997 1.87790774e-07 4.99999997 1.87890774e-07 4.99999997 1.87990774e-07 4.99999997 1.88090774e-07 4.99999997 1.88190774e-07 4.99999997 1.88290774e-07 4.99999997 1.88390774e-07 4.99999997
+ 1.88490774e-07 4.99999997 1.88590774e-07 4.99999997 1.88690774e-07 4.99999997 1.88790774e-07 4.99999997 1.88890774e-07 4.99999997 1.88990774e-07 4.99999997 1.89090774e-07 4.99999997 1.89190774e-07 4.99999997
+ 1.89290774e-07 4.99999997 1.89390774e-07 4.99999997 1.89490774e-07 4.99999997 1.89590774e-07 4.99999997 1.89690774e-07 4.99999997 1.89790774e-07 4.99999997 1.89890774e-07 4.99999997 1.89990774e-07 4.99999997
+ 1.90090774e-07 4.99999997 1.90190774e-07 4.99999997 1.90290774e-07 4.99999997 1.90390774e-07 4.99999997 1.90490774e-07 4.99999997 1.90590774e-07 4.99999997 1.90690774e-07 4.99999997 1.90790774e-07 4.99999997
+ 1.90890774e-07 4.99999997 1.90990774e-07 4.99999997 1.91090774e-07 4.99999997 1.91190774e-07 4.99999997 1.91290774e-07 4.99999997 1.91390774e-07 4.99999997 1.91490774e-07 4.99999997 1.91590774e-07 4.99999997
+ 1.91690774e-07 4.99999997 1.91790774e-07 4.99999997 1.91890774e-07 4.99999997 1.91990774e-07 4.99999997 1.92090774e-07 4.99999997 1.92190774e-07 4.99999997 1.92290774e-07 4.99999997 1.92390774e-07 4.99999997
+ 1.92490774e-07 4.99999997 1.92590774e-07 4.99999997 1.92690774e-07 4.99999997 1.92790774e-07 4.99999997 1.92890774e-07 4.99999997 1.92990774e-07 4.99999997 1.93090774e-07 4.99999997 1.93190774e-07 4.99999997
+ 1.93290774e-07 4.99999997 1.93390774e-07 4.99999997 1.93490774e-07 4.99999997 1.93590774e-07 4.99999997 1.93690774e-07 4.99999997 1.93790774e-07 4.99999997 1.93890774e-07 4.99999997 1.93990774e-07 4.99999997
+ 1.94090774e-07 4.99999997 1.94190774e-07 4.99999997 1.94290774e-07 4.99999997 1.94390774e-07 4.99999997 1.94490774e-07 4.99999997 1.94590774e-07 4.99999997 1.94690774e-07 4.99999997 1.94790774e-07 4.99999997
+ 1.94890774e-07 4.99999997 1.94990774e-07 4.99999997 1.95090774e-07 4.99999997 1.95190774e-07 4.99999997 1.95290774e-07 4.99999997 1.95390774e-07 4.99999997 1.95490774e-07 4.99999997 1.95590774e-07 4.99999997
+ 1.95690774e-07 4.99999997 1.95790774e-07 4.99999997 1.95890774e-07 4.99999997 1.95990774e-07 4.99999997 1.96090774e-07 4.99999997 1.96190774e-07 4.99999997 1.96290774e-07 4.99999997 1.96390774e-07 4.99999997
+ 1.96490774e-07 4.99999997 1.96590774e-07 4.99999997 1.96690774e-07 4.99999997 1.96790774e-07 4.99999997 1.96890774e-07 4.99999997 1.96990774e-07 4.99999997 1.97090774e-07 4.99999997 1.97190774e-07 4.99999997
+ 1.97290774e-07 4.99999997 1.97390774e-07 4.99999997 1.97490774e-07 4.99999997 1.97590774e-07 4.99999997 1.97690774e-07 4.99999997 1.97790774e-07 4.99999997 1.97890774e-07 4.99999997 1.97990774e-07 4.99999997
+ 1.98090774e-07 4.99999997 1.98190774e-07 4.99999997 1.98290774e-07 4.99999997 1.98390774e-07 4.99999997 1.98490774e-07 4.99999997 1.98590774e-07 4.99999997 1.98690774e-07 4.99999997 1.98790774e-07 4.99999997
+ 1.98890774e-07 4.99999997 1.98990774e-07 4.99999997 1.99090774e-07 4.99999997 1.99190774e-07 4.99999997 1.99290774e-07 4.99999997 1.99390774e-07 4.99999997 1.99490774e-07 4.99999997 1.99590774e-07 4.99999997
+ 1.99690774e-07 4.99999997 1.99790774e-07 4.99999997 1.99890774e-07 4.99999997 1.99990774e-07 4.99999997 2e-07 4.99999997 2.0001e-07 4.99999997 2.0003e-07 4.99999997 2.0007e-07 4.99999997
+ 2.0015e-07 4.99999997 2.0025e-07 4.99999997 2.0035e-07 4.99999997 2.0045e-07 4.99999997 2.0055e-07 4.99999997 2.0065e-07 4.99999997 2.0075e-07 5.00000001 2.0085e-07 4.99999718
+ 2.00932239e-07 5.00000338 2.01e-07 5.00008492 2.01008502e-07 5.000115 2.01025505e-07 5.00022464 2.01059511e-07 4.99960722 2.01090728e-07 4.99799758 2.01143656e-07 4.99699984 2.01199398e-07 5.02510852
+ 2.01276452e-07 4.95223975 2.01342062e-07 2.70342682 2.01411951e-07 0.0431011932 2.01487979e-07 0.0413288898 2.01566956e-07 -0.0198570509 2.01643585e-07 0.0200526747 2.01743585e-07 -0.0178801195 2.01843585e-07 0.0163673972
+ 2.01943585e-07 -0.0148974057 2.02043585e-07 0.0136306143 2.02143585e-07 -0.0124132097 2.02243585e-07 0.0113552946 2.02343585e-07 -0.0103461822 2.02443585e-07 0.0094630689 2.02543585e-07 -0.00862578629 2.02643585e-07 0.00788868402
+ 2.02743585e-07 -0.00719330222 2.02843585e-07 0.00657807192 2.02943585e-07 -0.006000042 2.03043585e-07 0.00548651241 2.03143585e-07 -0.00500567123 2.03243585e-07 0.00457700773 2.03343585e-07 -0.00417676053 2.03443585e-07 0.00381891884
+ 2.03543585e-07 -0.0034855792 2.03643585e-07 0.00318684373 2.03743585e-07 -0.00290910243 2.03843585e-07 0.00265969964 2.03943585e-07 -0.00242819624 2.04043585e-07 0.00221997183 2.04143585e-07 -0.00202694784 2.04243585e-07 0.00185309768
+ 2.04343585e-07 -0.00169211461 2.04443585e-07 0.00154696059 2.04543585e-07 -0.00141266991 2.04643585e-07 0.00129147307 2.04743585e-07 -0.00117942793 2.04843585e-07 0.00107823278 2.04943585e-07 -0.000984733296 2.05043585e-07 0.000900238043
+ 2.05143585e-07 -0.000822203994 2.05243585e-07 0.000751652326 2.05343585e-07 -0.000684967497 2.05443585e-07 0.000628009411 2.05543585e-07 -0.000573313512 2.05643585e-07 0.000524119197 2.05743585e-07 -0.000478719923 2.05843585e-07 0.000437643874
+ 2.05943585e-07 -0.000399739745 2.06043585e-07 0.000365442996 2.06143585e-07 -0.000333794097 2.06243585e-07 0.00030515815 2.06343585e-07 -0.000278730355 2.06443585e-07 0.000254821376 2.06543585e-07 -0.00023159652 2.06643585e-07 0.000212980054
+ 2.06743585e-07 -0.000193420857 2.06843585e-07 0.000177921478 2.06943585e-07 -0.000161548089 2.07043585e-07 0.000149658205 2.07143585e-07 -0.000134776618 2.07243585e-07 0.000124935858 2.07343585e-07 -0.000112502013 2.07443585e-07 0.00010430023
+ 2.07543585e-07 -9.39128182e-05 2.07643585e-07 8.7076031e-05 2.07743585e-07 -7.83977713e-05 2.07843585e-07 7.26984165e-05 2.07943585e-07 -6.54475826e-05 2.08043585e-07 6.06963617e-05 2.08143585e-07 -5.46376243e-05 2.08243585e-07 5.06769633e-05
+ 2.08343585e-07 -4.56137591e-05 2.08443585e-07 4.23124246e-05 2.08543585e-07 -3.80805791e-05 2.08643585e-07 3.53292281e-05 2.08743585e-07 -3.1791625e-05 2.08843585e-07 2.9499122e-05 2.08943585e-07 -2.65412486e-05 2.09043585e-07 2.46316109e-05
+ 2.09143585e-07 -2.21578353e-05 2.09243585e-07 2.05676984e-05 2.09343585e-07 -1.84981586e-05 2.09443585e-07 1.71746699e-05 2.09543585e-07 -1.5442675e-05 2.09643585e-07 1.43417422e-05 2.09743585e-07 -1.28916015e-05 2.09843585e-07 1.19764355e-05
+ 2.09943585e-07 -1.07616446e-05 2.10043585e-07 1.00015461e-05 2.10143585e-07 -8.98327234e-06 2.10243585e-07 8.35262224e-06 2.10343585e-07 -7.49844226e-06 2.10443585e-07 6.97585964e-06 2.10543585e-07 -6.25869755e-06 2.10643585e-07 5.82633423e-06
+ 2.10743585e-07 -5.22358013e-06 2.10843585e-07 4.86653702e-06 2.10943585e-07 -4.35931147e-06 2.11043585e-07 4.06515128e-06 2.11143585e-07 -3.63768999e-06 2.11243585e-07 3.39603008e-06 2.11343585e-07 -3.03517004e-06 2.11443585e-07 2.8373427e-06
+ 2.11543585e-07 -2.53209303e-06 2.11643585e-07 2.37085708e-06 2.11743585e-07 -2.11203389e-06 2.11843585e-07 1.98135588e-06 2.11943585e-07 -1.76130989e-06 2.12043585e-07 1.65614584e-06 2.12143585e-07 -1.46847298e-06 2.12243585e-07 1.38460953e-06
+ 2.12343585e-07 -1.22396639e-06 2.12443585e-07 1.15788736e-06 2.12543585e-07 -1.01981312e-06 2.12643585e-07 9.68583023e-07 2.12743585e-07 -8.49353045e-07 2.12843585e-07 8.10520995e-07 2.12943585e-07 -7.07025356e-07 2.13043585e-07 6.78545058e-07
+ 2.13143585e-07 -5.88187152e-07 2.13243585e-07 5.68350126e-07 2.13343585e-07 -4.88961596e-07 2.13443585e-07 4.76341167e-07 2.13543585e-07 -4.06111844e-07 2.13643585e-07 3.9951709e-07 2.13743585e-07 -3.3693541e-07 2.13843585e-07 3.35371832e-07
+ 2.13943585e-07 -2.79175661e-07 2.14043585e-07 2.81812899e-07 2.14143585e-07 -2.30948406e-07 2.14243585e-07 2.37093158e-07 2.14343585e-07 -1.90680431e-07 2.14443585e-07 1.99753818e-07 2.14543585e-07 -1.57058162e-07 2.14643585e-07 1.68576846e-07
+ 2.14743585e-07 -1.28984815e-07 2.14843585e-07 1.42545229e-07 2.14943585e-07 -1.05544617e-07 2.15043585e-07 1.208098e-07 2.15143585e-07 -8.59729298e-08 2.15243585e-07 1.0266153e-07 2.15343585e-07 -6.96340728e-08 2.15443585e-07 8.7513677e-08
+ 2.15543585e-07 -5.59972484e-08 2.15643585e-07 7.48717104e-08 2.15743585e-07 -4.46163243e-08 2.15843585e-07 6.43210657e-08 2.15943585e-07 -3.51181101e-08 2.16043585e-07 5.55157795e-08 2.16143585e-07 -2.71911566e-08 2.16243585e-07 4.81671261e-08
+ 2.16343585e-07 -2.05755378e-08 2.16443585e-07 4.20341418e-08 2.16543585e-07 -1.50403404e-08 2.16643585e-07 3.69030002e-08 2.16743585e-07 -1.04355915e-08 2.16843585e-07 3.26339483e-08 2.16943585e-07 -6.59228291e-09 2.17043585e-07 2.90710202e-08
+ 2.17143585e-07 -3.38468492e-09 2.17243585e-07 2.60974319e-08 2.17343585e-07 -7.07656128e-10 2.17443585e-07 2.36157067e-08 2.17543585e-07 1.52656177e-09 2.17643585e-07 2.15643594e-08 2.17743585e-07 3.37429304e-09 2.17843585e-07 1.98754834e-08
+ 2.17943585e-07 4.89591356e-09 2.18043585e-07 1.84846787e-08 2.18143585e-07 6.14898474e-09 2.18243585e-07 1.73393341e-08 2.18343585e-07 7.18090426e-09 2.18443585e-07 1.63961289e-08 2.18543585e-07 8.03070199e-09 2.18643585e-07 1.56193891e-08
+ 2.18743585e-07 8.73051897e-09 2.18843585e-07 1.48828709e-08 2.18943585e-07 9.2930609e-09 2.19043585e-07 1.43671893e-08 2.19143585e-07 9.76114548e-09 2.19243585e-07 1.39422635e-08 2.19343585e-07 1.01468813e-08 2.19443585e-07 1.35921051e-08
+ 2.19543585e-07 1.04647401e-08 2.19643585e-07 1.33035664e-08 2.19743585e-07 1.07266619e-08 2.19843585e-07 1.30658054e-08 2.19943585e-07 1.0942489e-08 2.20043585e-07 1.28698879e-08 2.20143585e-07 1.11203326e-08 2.20243585e-07 1.27084502e-08
+ 2.20343585e-07 1.12668763e-08 2.20443585e-07 1.25754253e-08 2.20543585e-07 1.13876288e-08 2.20643585e-07 1.24658124e-08 2.20743585e-07 1.14871286e-08 2.20843585e-07 1.23754919e-08 2.20943585e-07 1.15691153e-08 2.21043585e-07 1.2301069e-08
+ 2.21143585e-07 1.16366711e-08 2.21243585e-07 1.22397455e-08 2.21343585e-07 1.16923362e-08 2.21443585e-07 1.21892161e-08 2.21543585e-07 1.17382027e-08 2.21643585e-07 1.21475811e-08 2.21743585e-07 1.17759955e-08 2.21843585e-07 1.21132755e-08
+ 2.21943585e-07 1.18071349e-08 2.22043585e-07 1.20850087e-08 2.22143585e-07 1.18327928e-08 2.22243585e-07 1.20617189e-08 2.22343585e-07 1.18539328e-08 2.22443585e-07 1.20425292e-08 2.22543585e-07 1.18713514e-08 2.22643585e-07 1.20267178e-08
+ 2.22743585e-07 1.1885703e-08 2.22843585e-07 1.20136909e-08 2.22943585e-07 1.18975271e-08 2.23043585e-07 1.20029578e-08 2.23143585e-07 1.1907269e-08 2.23243585e-07 1.19941146e-08 2.23343585e-07 1.19152953e-08 2.23443585e-07 1.19868293e-08
+ 2.23543585e-07 1.19219077e-08 2.23643585e-07 1.19808266e-08 2.23743585e-07 1.19273557e-08 2.23843585e-07 1.19758821e-08 2.23943585e-07 1.19318434e-08 2.24043585e-07 1.19718082e-08 2.24143585e-07 1.19355402e-08 2.24243585e-07 1.19684525e-08
+ 2.24343585e-07 1.19385861e-08 2.24443585e-07 1.19656879e-08 2.24543585e-07 1.19410951e-08 2.24643585e-07 1.19634105e-08 2.24743585e-07 1.19431615e-08 2.24843585e-07 1.19615347e-08 2.24943585e-07 1.19448637e-08 2.25043585e-07 1.19599898e-08
+ 2.25143585e-07 1.19462654e-08 2.25243585e-07 1.19587167e-08 2.25343585e-07 1.19474204e-08 2.25443585e-07 1.19576687e-08 2.25543585e-07 1.19483713e-08 2.25643585e-07 1.19568055e-08 2.25743585e-07 1.19491542e-08 2.25843585e-07 1.19560949e-08
+ 2.25943585e-07 1.19497993e-08 2.26043585e-07 1.19555094e-08 2.26143585e-07 1.19503303e-08 2.26243585e-07 1.19550274e-08 2.26343585e-07 1.19507672e-08 2.26443585e-07 1.19546309e-08 2.26543585e-07 1.19511272e-08 2.26643585e-07 1.19543036e-08
+ 2.26743585e-07 1.19514236e-08 2.26843585e-07 1.1954035e-08 2.26943585e-07 1.19516674e-08 2.27043585e-07 1.19538137e-08 2.27143585e-07 1.19518677e-08 2.27243585e-07 1.19536313e-08 2.27343585e-07 1.19520331e-08 2.27443585e-07 1.19534814e-08
+ 2.27543585e-07 1.19521688e-08 2.27643585e-07 1.19533582e-08 2.27743585e-07 1.19522802e-08 2.27843585e-07 1.19532564e-08 2.27943585e-07 1.19523724e-08 2.28043585e-07 1.19531732e-08 2.28143585e-07 1.19524476e-08 2.28243585e-07 1.19531045e-08
+ 2.28343585e-07 1.19525098e-08 2.28443585e-07 1.19530484e-08 2.28543585e-07 1.19525608e-08 2.28643585e-07 1.19530015e-08 2.28743585e-07 1.19526027e-08 2.28843585e-07 1.19529636e-08 2.28943585e-07 1.1952637e-08 2.29043585e-07 1.19529323e-08
+ 2.29143585e-07 1.19526655e-08 2.29243585e-07 1.19529064e-08 2.29343585e-07 1.19526888e-08 2.29443585e-07 1.19528851e-08 2.29543585e-07 1.19527077e-08 2.29643585e-07 1.19528681e-08 2.29743585e-07 1.19527232e-08 2.29843585e-07 1.19528539e-08
+ 2.29943585e-07 1.19527359e-08 2.30043585e-07 1.19528422e-08 2.30143585e-07 1.19527462e-08 2.30243585e-07 1.19528327e-08 2.30343585e-07 1.19527548e-08 2.30443585e-07 1.19528248e-08 2.30543585e-07 1.19527616e-08 2.30643585e-07 1.19528183e-08
+ 2.30743585e-07 1.19527674e-08 2.30843585e-07 1.19528133e-08 2.30943585e-07 1.19527717e-08 2.31043585e-07 1.1952809e-08 2.31143585e-07 1.1952776e-08 2.31243585e-07 1.19528054e-08 2.31343585e-07 1.19527788e-08 2.31443585e-07 1.19528025e-08
+ 2.31543585e-07 1.19527814e-08 2.31643585e-07 1.19528002e-08 2.31743585e-07 1.19527834e-08 2.31843585e-07 1.19527982e-08 2.31943585e-07 1.19527851e-08 2.32043585e-07 1.19527966e-08 2.32143585e-07 1.19527862e-08 2.32243585e-07 1.19527955e-08
+ 2.32343585e-07 1.19527874e-08 2.32443585e-07 1.19527944e-08 2.32543585e-07 1.19527881e-08 2.32643585e-07 1.19527938e-08 2.32743585e-07 1.19527885e-08 2.32843585e-07 1.19527929e-08 2.32943585e-07 1.19527892e-08 2.33043585e-07 1.19527924e-08
+ 2.33143585e-07 1.19527897e-08 2.33243585e-07 1.19527916e-08 2.33343585e-07 1.19527899e-08 2.33443585e-07 1.19527915e-08 2.33543585e-07 1.19527903e-08 2.33643585e-07 1.19527911e-08 2.33743585e-07 1.19527903e-08 2.33843585e-07 1.19527909e-08
+ 2.33943585e-07 1.19527906e-08 2.34043585e-07 1.1952791e-08 2.34143585e-07 1.19527905e-08 2.34243585e-07 1.19527908e-08 2.34343585e-07 1.19527905e-08 2.34443585e-07 1.19527908e-08 2.34543585e-07 1.19527905e-08 2.34643585e-07 1.19527907e-08
+ 2.34743585e-07 1.19527906e-08 2.34843585e-07 1.19527905e-08 2.34943585e-07 1.19527903e-08 2.35043585e-07 1.19527905e-08 2.35143585e-07 1.19527907e-08 2.35243585e-07 1.19527902e-08 2.35343585e-07 1.19527905e-08 2.35443585e-07 1.19527902e-08
+ 2.35543585e-07 1.19527905e-08 2.35643585e-07 1.19527902e-08 2.35743585e-07 1.19527906e-08 2.35843585e-07 1.19527902e-08 2.35943585e-07 1.19527903e-08 2.36043585e-07 1.19527901e-08 2.36143585e-07 1.19527903e-08 2.36243585e-07 1.19527904e-08
+ 2.36343585e-07 1.19527902e-08 2.36443585e-07 1.195279e-08 2.36543585e-07 1.19527905e-08 2.36643585e-07 1.19527901e-08 2.36743585e-07 1.195279e-08 2.36843585e-07 1.19527903e-08 2.36943585e-07 1.19527901e-08 2.37043585e-07 1.19527902e-08
+ 2.37143585e-07 1.19527901e-08 2.37243585e-07 1.19527901e-08 2.37343585e-07 1.19527903e-08 2.37443585e-07 1.19527899e-08 2.37543585e-07 1.19527903e-08 2.37643585e-07 1.195279e-08 2.37743585e-07 1.19527902e-08 2.37843585e-07 1.19527901e-08
+ 2.37943585e-07 1.19527901e-08 2.38043585e-07 1.19527898e-08 2.38143585e-07 1.19527901e-08 2.38243585e-07 1.195279e-08 2.38343585e-07 1.19527901e-08 2.38443585e-07 1.195279e-08 2.38543585e-07 1.195279e-08 2.38643585e-07 1.195279e-08
+ 2.38743585e-07 1.195279e-08 2.38843585e-07 1.195279e-08 2.38943585e-07 1.19527899e-08 2.39043585e-07 1.195279e-08 2.39143585e-07 1.19527898e-08 2.39243585e-07 1.19527898e-08 2.39343585e-07 1.19527897e-08 2.39443585e-07 1.19527901e-08
+ 2.39543585e-07 1.19527897e-08 2.39643585e-07 1.19527898e-08 2.39743585e-07 1.19527896e-08 2.39843585e-07 1.195279e-08 2.39943585e-07 1.19527894e-08 2.40043585e-07 1.19527897e-08 2.40143585e-07 1.19527898e-08 2.40243585e-07 1.19527895e-08
+ 2.40343585e-07 1.19527898e-08 2.40443585e-07 1.19527896e-08 2.40543585e-07 1.19527897e-08 2.40643585e-07 1.19527897e-08 2.40743585e-07 1.19527899e-08 2.40843585e-07 1.19527898e-08 2.40943585e-07 1.19527896e-08 2.41043585e-07 1.19527895e-08
+ 2.41143585e-07 1.19527897e-08 2.41243585e-07 1.19527896e-08 2.41343585e-07 1.19527898e-08 2.41443585e-07 1.19527896e-08 2.41543585e-07 1.19527897e-08 2.41643585e-07 1.19527897e-08 2.41743585e-07 1.19527895e-08 2.41843585e-07 1.19527896e-08
+ 2.41943585e-07 1.19527896e-08 2.42043585e-07 1.19527898e-08 2.42143585e-07 1.19527895e-08 2.42243585e-07 1.19527897e-08 2.42343585e-07 1.19527895e-08 2.42443585e-07 1.19527898e-08 2.42543585e-07 1.19527893e-08 2.42643585e-07 1.19527894e-08
+ 2.42743585e-07 1.19527892e-08 2.42843585e-07 1.19527898e-08 2.42943585e-07 1.19527893e-08 2.43043585e-07 1.19527898e-08 2.43143585e-07 1.19527893e-08 2.43243585e-07 1.19527895e-08 2.43343585e-07 1.19527894e-08 2.43443585e-07 1.19527896e-08
+ 2.43543585e-07 1.19527895e-08 2.43643585e-07 1.19527896e-08 2.43743585e-07 1.19527891e-08 2.43843585e-07 1.19527892e-08 2.43943585e-07 1.19527891e-08 2.44043585e-07 1.19527896e-08 2.44143585e-07 1.19527892e-08 2.44243585e-07 1.19527897e-08
+ 2.44343585e-07 1.1952789e-08 2.44443585e-07 1.19527895e-08 2.44543585e-07 1.19527892e-08 2.44643585e-07 1.19527894e-08 2.44743585e-07 1.19527891e-08 2.44843585e-07 1.19527895e-08 2.44943585e-07 1.1952789e-08 2.45043585e-07 1.19527893e-08
+ 2.45143585e-07 1.1952789e-08 2.45243585e-07 1.19527893e-08 2.45343585e-07 1.19527893e-08 2.45443585e-07 1.19527893e-08 2.45543585e-07 1.19527891e-08 2.45643585e-07 1.19527891e-08 2.45743585e-07 1.19527896e-08 2.45843585e-07 1.19527892e-08
+ 2.45943585e-07 1.19527895e-08 2.46043585e-07 1.19527893e-08 2.46143585e-07 1.1952789e-08 2.46243585e-07 1.19527891e-08 2.46343585e-07 1.1952789e-08 2.46443585e-07 1.19527893e-08 2.46543585e-07 1.19527894e-08 2.46643585e-07 1.1952789e-08
+ 2.46743585e-07 1.19527894e-08 2.46843585e-07 1.1952789e-08 2.46943585e-07 1.19527893e-08 2.47043585e-07 1.1952789e-08 2.47143585e-07 1.19527892e-08 2.47243585e-07 1.19527893e-08 2.47343585e-07 1.19527891e-08 2.47443585e-07 1.19527893e-08
+ 2.47543585e-07 1.19527891e-08 2.47643585e-07 1.1952789e-08 2.47743585e-07 1.19527892e-08 2.47843585e-07 1.19527891e-08 2.47943585e-07 1.19527891e-08 2.48043585e-07 1.19527891e-08 2.48143585e-07 1.19527891e-08 2.48243585e-07 1.19527892e-08
+ 2.48343585e-07 1.1952789e-08 2.48443585e-07 1.19527894e-08 2.48543585e-07 1.19527889e-08 2.48643585e-07 1.19527893e-08 2.48743585e-07 1.19527888e-08 2.48843585e-07 1.19527892e-08 2.48943585e-07 1.19527891e-08 2.49043585e-07 1.19527892e-08
+ 2.49143585e-07 1.19527891e-08 2.49243585e-07 1.19527893e-08 2.49343585e-07 1.19527887e-08 2.49443585e-07 1.19527889e-08 2.49543585e-07 1.19527889e-08 2.49643585e-07 1.19527892e-08 2.49743585e-07 1.19527891e-08 2.49843585e-07 1.19527893e-08
+ 2.49943585e-07 1.1952789e-08 2.50043585e-07 1.19527893e-08 2.50143585e-07 1.1952789e-08 2.50243585e-07 1.19527893e-08 2.50343585e-07 1.1952789e-08 2.50443585e-07 1.19527887e-08 2.50543585e-07 1.19527891e-08 2.50643585e-07 1.1952789e-08
+ 2.50743585e-07 1.19527892e-08 2.50843585e-07 1.19527889e-08 2.50943585e-07 1.19527892e-08 2.51e-07 1.19527886e-08 2.5101e-07 1.19387336e-08 2.5103e-07 1.20209579e-08 2.5107e-07 1.1845657e-08 2.5115e-07 1.20751984e-08
+ 2.5125e-07 1.1825728e-08 2.5135e-07 1.20743629e-08 2.5145e-07 1.18466581e-08 2.5155e-07 1.20361451e-08 2.5165e-07 1.1895076e-08 2.5175e-07 1.19816164e-08 2.5185e-07 1.19573519e-08 2.51930828e-07 1.29898242e-07
+ 2.52e-07 1.68693818e-06 2.52008608e-07 -4.63455704e-06 2.52025825e-07 -7.9808205e-06 2.52060258e-07 1.5061975e-06 2.52106181e-07 1.0973022e-05 2.52150081e-07 -1.19545368e-05 2.52198026e-07 8.69407647e-06 2.5225538e-07 -7.92726691e-06
+ 2.52312019e-07 6.0886179e-06 2.52404231e-07 -4.35191802e-06 2.52504231e-07 2.87067141e-06 2.52604231e-07 -1.60647351e-06 2.52704231e-07 7.09383149e-07 2.52804231e-07 6.21050557e-08 2.52904231e-07 -6.67617034e-07 2.53004231e-07 1.2280794e-06
+ 2.53104231e-07 -1.66857258e-06 2.53204231e-07 2.08522619e-06 2.53304231e-07 -2.39320129e-06 2.53404231e-07 2.68781493e-06 2.53504231e-07 -2.88197065e-06 2.53604231e-07 3.07280994e-06 2.53704231e-07 -3.17200642e-06 2.53804231e-07 3.2781936e-06
+ 2.53904231e-07 -3.30170758e-06 2.54004231e-07 3.34196797e-06 2.54104231e-07 -3.30788027e-06 2.54204231e-07 3.2991216e-06 2.54304231e-07 -3.2232367e-06 2.54404231e-07 3.17983294e-06 2.54504231e-07 -3.07526771e-06 2.54604231e-07 3.00890095e-06
+ 2.54704231e-07 -2.88611918e-06 2.54804231e-07 2.80595288e-06 2.54904231e-07 -2.67303462e-06 2.55004231e-07 2.58603942e-06 2.55104231e-07 -2.44904115e-06 2.55204231e-07 2.36036454e-06 2.55304231e-07 -2.22368841e-06 2.55404231e-07 2.13700757e-06
+ 2.55504231e-07 -2.00373963e-06 2.55604231e-07 1.92157875e-06 2.55704231e-07 -1.79378453e-06 2.55804231e-07 1.71778029e-06 2.55904231e-07 -1.59674487e-06 2.56004231e-07 1.52786046e-06 2.56104231e-07 -1.41428355e-06 2.56204231e-07 1.3529841e-06
+ 2.56304231e-07 -1.24713754e-06 2.56404231e-07 1.19352802e-06 2.56504231e-07 -1.09537836e-06 2.56604231e-07 1.04931085e-06 2.56704231e-07 -9.58614229e-07 2.56804231e-07 9.1976977e-07 2.56904231e-07 -8.36142431e-07 2.57004231e-07 8.04091186e-07
+ 2.57104231e-07 -7.27063187e-07 2.57204231e-07 7.01312281e-07 2.57304231e-07 -6.30369486e-07 2.57404231e-07 6.10398102e-07 2.57504231e-07 -5.45011509e-07 2.57604231e-07 5.30294844e-07 2.57704231e-07 -4.69940202e-07 2.57804231e-07 4.59965237e-07
+ 2.57904231e-07 -4.04136037e-07 2.58004231e-07 3.98412181e-07 2.58104231e-07 -3.46628439e-07 2.58204231e-07 3.44694536e-07 2.58304231e-07 -2.96508307e-07 2.58404231e-07 2.97936752e-07 2.58504231e-07 -2.52935085e-07 2.58604231e-07 2.57333733e-07
+ 2.58704231e-07 -2.1513933e-07 2.58804231e-07 2.22150053e-07 2.58904231e-07 -1.82418412e-07 2.59004231e-07 1.91716469e-07 2.59104231e-07 -1.54139153e-07 2.59204231e-07 1.65436835e-07 2.59304231e-07 -1.29741724e-07 2.59404231e-07 1.42784958e-07
+ 2.59504231e-07 -1.08731077e-07 2.59604231e-07 1.23294537e-07 2.59704231e-07 -9.06683014e-08 2.59804231e-07 1.06552593e-07 2.59904231e-07 -7.5165328e-08 2.60004231e-07 9.21946308e-08 2.60104231e-07 -6.1880455e-08 2.60204231e-07 7.9901253e-08
+ 2.60304231e-07 -5.05158949e-08 2.60404231e-07 6.93947394e-08 2.60504231e-07 -4.08130819e-08 2.60604231e-07 6.04320325e-08 2.60704231e-07 -3.25414545e-08 2.60804231e-07 5.2796264e-08 2.60904231e-07 -2.54989314e-08 2.61004231e-07 4.6299143e-08
+ 2.61104231e-07 -1.95102627e-08 2.61204231e-07 4.07775695e-08 2.61304231e-07 -1.44238234e-08 2.61404231e-07 3.60905903e-08 2.61504231e-07 -1.01087192e-08 2.61604231e-07 3.21166455e-08 2.61704231e-07 -6.45216364e-09 2.61804231e-07 2.87510622e-08
+ 2.61904231e-07 -3.35709149e-09 2.62004231e-07 2.59038327e-08 2.62104231e-07 -7.40147277e-10 2.62204231e-07 2.34977895e-08 2.62304231e-07 1.46047893e-09 2.62404231e-07 2.14846642e-08 2.62504231e-07 3.29716074e-09 2.62604231e-07 1.98091944e-08
+ 2.62704231e-07 4.82515078e-09 2.62804231e-07 1.84160882e-08 2.62904231e-07 6.09492229e-09 2.63004231e-07 1.72590652e-08 2.63104231e-07 7.1488967e-09 2.63204231e-07 1.62992531e-08 2.63304231e-07 8.02268585e-09 2.63404231e-07 1.55040344e-08
+ 2.63504231e-07 8.74615708e-09 2.63604231e-07 1.4846065e-08 2.63704231e-07 9.34433927e-09 2.63804231e-07 1.43024405e-08 2.63904231e-07 9.83818957e-09 2.64004231e-07 1.38540379e-08 2.64104231e-07 1.0245185e-08 2.64204231e-07 1.34848203e-08
+ 2.64304231e-07 1.05797129e-08 2.64404231e-07 1.31818536e-08 2.64504231e-07 1.08542378e-08 2.64604231e-07 1.29330901e-08 2.64704231e-07 1.10795437e-08 2.64804231e-07 1.27292158e-08 2.64904231e-07 1.12638395e-08 2.65004231e-07 1.25627462e-08
+ 2.65104231e-07 1.1414136e-08 2.65204231e-07 1.24270859e-08 2.65304231e-07 1.15365051e-08 2.65404231e-07 1.23168961e-08 2.65504231e-07 1.1635532e-08 2.65604231e-07 1.22280073e-08 2.65704231e-07 1.171526e-08 2.65804231e-07 1.21565573e-08
+ 2.65904231e-07 1.17792246e-08 2.66004231e-07 1.2099364e-08 2.66104231e-07 1.18302939e-08 2.66204231e-07 1.20538321e-08 2.66304231e-07 1.18708183e-08 2.66404231e-07 1.20178359e-08 2.66504231e-07 1.19027241e-08 2.66604231e-07 1.19896193e-08
+ 2.66704231e-07 1.19276162e-08 2.66804231e-07 1.1967644e-08 2.66904231e-07 1.1946949e-08 2.67004231e-07 1.19508729e-08 2.67104231e-07 1.19614317e-08 2.67204231e-07 1.19383219e-08 2.67304231e-07 1.19722687e-08 2.67404231e-07 1.19290235e-08
+ 2.67504231e-07 1.19801837e-08 2.67604231e-07 1.19223498e-08 2.67704231e-07 1.1985747e-08 2.67804231e-07 1.19177779e-08 2.67904231e-07 1.19894367e-08 2.68004231e-07 1.19148712e-08 2.68104231e-07 1.19916496e-08 2.68204231e-07 1.19132703e-08
+ 2.68304231e-07 1.19927118e-08 2.68404231e-07 1.19126811e-08 2.68504231e-07 1.19929031e-08 2.68604231e-07 1.19128184e-08 2.68704231e-07 1.19924516e-08 2.68804231e-07 1.19135801e-08 2.68904231e-07 1.19914318e-08 2.69004231e-07 1.19147993e-08
+ 2.69104231e-07 1.19900505e-08 2.69204231e-07 1.19163129e-08 2.69304231e-07 1.19884327e-08 2.69404231e-07 1.19180125e-08 2.69504231e-07 1.19866635e-08 2.69604231e-07 1.19198409e-08 2.69704231e-07 1.19847905e-08 2.69804231e-07 1.19217441e-08
+ 2.69904231e-07 1.19828699e-08 2.70004231e-07 1.19236704e-08 2.70104231e-07 1.19809475e-08 2.70204231e-07 1.19255817e-08 2.70304231e-07 1.1979054e-08 2.70404231e-07 1.19274516e-08 2.70504231e-07 1.19772123e-08 2.70604231e-07 1.19292608e-08
+ 2.70704231e-07 1.19754388e-08 2.70804231e-07 1.19309963e-08 2.70904231e-07 1.19737436e-08 2.71004231e-07 1.19326491e-08 2.71104231e-07 1.19721346e-08 2.71204231e-07 1.19342135e-08 2.71304231e-07 1.19706149e-08 2.71404231e-07 1.19356876e-08
+ 2.71504231e-07 1.19691865e-08 2.71604231e-07 1.19370709e-08 2.71704231e-07 1.19678489e-08 2.71804231e-07 1.1938363e-08 2.71904231e-07 1.19666017e-08 2.72004231e-07 1.1939566e-08 2.72104231e-07 1.19654423e-08 2.72204231e-07 1.19406826e-08
+ 2.72304231e-07 1.19643671e-08 2.72404231e-07 1.19417169e-08 2.72504231e-07 1.19633726e-08 2.72604231e-07 1.19426724e-08 2.72704231e-07 1.19624554e-08 2.72804231e-07 1.19435533e-08 2.72904231e-07 1.19616099e-08 2.73004231e-07 1.1944364e-08
+ 2.73104231e-07 1.19608332e-08 2.73204231e-07 1.19451074e-08 2.73304231e-07 1.19601217e-08 2.73404231e-07 1.19457901e-08 2.73504231e-07 1.19594656e-08 2.73604231e-07 1.19464194e-08 2.73704231e-07 1.19588637e-08 2.73804231e-07 1.19469943e-08
+ 2.73904231e-07 1.19583143e-08 2.74004231e-07 1.19475187e-08 2.74104231e-07 1.19578139e-08 2.74204231e-07 1.19479968e-08 2.74304231e-07 1.19573574e-08 2.74404231e-07 1.19484326e-08 2.74504231e-07 1.19569411e-08 2.74604231e-07 1.19488295e-08
+ 2.74704231e-07 1.19565625e-08 2.74804231e-07 1.19491911e-08 2.74904231e-07 1.19562177e-08 2.75004231e-07 1.19495198e-08 2.75104231e-07 1.19559041e-08 2.75204231e-07 1.1949819e-08 2.75304231e-07 1.19556191e-08 2.75404231e-07 1.19500907e-08
+ 2.75504231e-07 1.19553598e-08 2.75604231e-07 1.19503385e-08 2.75704231e-07 1.19551227e-08 2.75804231e-07 1.19505643e-08 2.75904231e-07 1.19549074e-08 2.76004231e-07 1.19507698e-08 2.76104231e-07 1.19547122e-08 2.76204231e-07 1.19509557e-08
+ 2.76304231e-07 1.19545349e-08 2.76404231e-07 1.19511244e-08 2.76504231e-07 1.19543742e-08 2.76604231e-07 1.19512773e-08 2.76704231e-07 1.19542286e-08 2.76804231e-07 1.19514159e-08 2.76904231e-07 1.19540967e-08 2.77004231e-07 1.19515417e-08
+ 2.77104231e-07 1.19539768e-08 2.77204231e-07 1.19516557e-08 2.77304231e-07 1.1953868e-08 2.77404231e-07 1.19517596e-08 2.77504231e-07 1.19537691e-08 2.77604231e-07 1.19518537e-08 2.77704231e-07 1.19536793e-08 2.77804231e-07 1.19519392e-08
+ 2.77904231e-07 1.19535979e-08 2.78004231e-07 1.19520171e-08 2.78104231e-07 1.19535237e-08 2.78204231e-07 1.19520876e-08 2.78304231e-07 1.19534564e-08 2.78404231e-07 1.19521517e-08 2.78504231e-07 1.19533954e-08 2.78604231e-07 1.19522099e-08
+ 2.78704231e-07 1.19533396e-08 2.78804231e-07 1.19522632e-08 2.78904231e-07 1.19532892e-08 2.79004231e-07 1.19523111e-08 2.79104231e-07 1.19532434e-08 2.79204231e-07 1.19523551e-08 2.79304231e-07 1.19532014e-08 2.79404231e-07 1.19523949e-08
+ 2.79504231e-07 1.19531635e-08 2.79604231e-07 1.1952431e-08 2.79704231e-07 1.19531292e-08 2.79804231e-07 1.19524637e-08 2.79904231e-07 1.19530979e-08 2.80004231e-07 1.19524935e-08 2.80104231e-07 1.19530695e-08 2.80204231e-07 1.19525208e-08
+ 2.80304231e-07 1.19530436e-08 2.80404231e-07 1.19525451e-08 2.80504231e-07 1.195302e-08 2.80604231e-07 1.1952568e-08 2.80704231e-07 1.19529988e-08 2.80804231e-07 1.19525882e-08 2.80904231e-07 1.19529793e-08 2.81004231e-07 1.19526065e-08
+ 2.81104231e-07 1.19529619e-08 2.81204231e-07 1.19526234e-08 2.81304231e-07 1.19529459e-08 2.81404231e-07 1.19526387e-08 2.81504231e-07 1.19529313e-08 2.81604231e-07 1.19526526e-08 2.81704231e-07 1.1952918e-08 2.81804231e-07 1.19526652e-08
+ 2.81904231e-07 1.19529059e-08 2.82004231e-07 1.19526767e-08 2.82104231e-07 1.1952895e-08 2.82204231e-07 1.19526866e-08 2.82304231e-07 1.19528852e-08 2.82404231e-07 1.19526961e-08 2.82504231e-07 1.19528764e-08 2.82604231e-07 1.1952705e-08
+ 2.82704231e-07 1.19528683e-08 2.82804231e-07 1.19527123e-08 2.82904231e-07 1.19528606e-08 2.83004231e-07 1.19527198e-08 2.83104231e-07 1.19528535e-08 2.83204231e-07 1.19527264e-08 2.83304231e-07 1.19528479e-08 2.83404231e-07 1.1952732e-08
+ 2.83504231e-07 1.19528422e-08 2.83604231e-07 1.19527371e-08 2.83704231e-07 1.19528371e-08 2.83804231e-07 1.19527419e-08 2.83904231e-07 1.19528328e-08 2.84004231e-07 1.19527464e-08 2.84104231e-07 1.19528285e-08 2.84204231e-07 1.19527503e-08
+ 2.84304231e-07 1.19528247e-08 2.84404231e-07 1.19527538e-08 2.84504231e-07 1.19528215e-08 2.84604231e-07 1.19527571e-08 2.84704231e-07 1.19528183e-08 2.84804231e-07 1.195276e-08 2.84904231e-07 1.19528156e-08 2.85004231e-07 1.19527629e-08
+ 2.85104231e-07 1.19528129e-08 2.85204231e-07 1.19527654e-08 2.85304231e-07 1.19528105e-08 2.85404231e-07 1.19527673e-08 2.85504231e-07 1.19528085e-08 2.85604231e-07 1.19527695e-08 2.85704231e-07 1.19528064e-08 2.85804231e-07 1.19527716e-08
+ 2.85904231e-07 1.19528049e-08 2.86004231e-07 1.1952773e-08 2.86104231e-07 1.19528032e-08 2.86204231e-07 1.19527744e-08 2.86304231e-07 1.19528017e-08 2.86404231e-07 1.19527758e-08 2.86504231e-07 1.19528007e-08 2.86604231e-07 1.19527767e-08
+ 2.86704231e-07 1.19527995e-08 2.86804231e-07 1.1952778e-08 2.86904231e-07 1.19527984e-08 2.87004231e-07 1.19527789e-08 2.87104231e-07 1.19527974e-08 2.87204231e-07 1.19527799e-08 2.87304231e-07 1.19527964e-08 2.87404231e-07 1.19527808e-08
+ 2.87504231e-07 1.19527958e-08 2.87604231e-07 1.19527814e-08 2.87704231e-07 1.1952795e-08 2.87804231e-07 1.19527823e-08 2.87904231e-07 1.19527944e-08 2.88004231e-07 1.19527826e-08 2.88104231e-07 1.19527938e-08 2.88204231e-07 1.19527831e-08
+ 2.88304231e-07 1.19527934e-08 2.88404231e-07 1.19527836e-08 2.88504231e-07 1.19527928e-08 2.88604231e-07 1.19527842e-08 2.88704231e-07 1.19527926e-08 2.88804231e-07 1.19527843e-08 2.88904231e-07 1.19527923e-08 2.89004231e-07 1.19527848e-08
+ 2.89104231e-07 1.19527923e-08 2.89204231e-07 1.19527851e-08 2.89304231e-07 1.19527917e-08 2.89404231e-07 1.19527854e-08 2.89504231e-07 1.19527914e-08 2.89604231e-07 1.19527857e-08 2.89704231e-07 1.19527908e-08 2.89804231e-07 1.1952786e-08
+ 2.89904231e-07 1.19527909e-08 2.90004231e-07 1.19527862e-08 2.90104231e-07 1.19527904e-08 2.90204231e-07 1.19527865e-08 2.90304231e-07 1.19527901e-08 2.90404231e-07 1.19527867e-08 2.90504231e-07 1.19527898e-08 2.90604231e-07 1.19527868e-08
+ 2.90704231e-07 1.19527896e-08 2.90804231e-07 1.19527872e-08 2.90904231e-07 1.19527897e-08 2.91004231e-07 1.19527873e-08 2.91104231e-07 1.19527897e-08 2.91204231e-07 1.19527875e-08 2.91304231e-07 1.19527894e-08 2.91404231e-07 1.19527875e-08
+ 2.91504231e-07 1.19527894e-08 2.91604231e-07 1.19527875e-08 2.91704231e-07 1.19527891e-08 2.91804231e-07 1.19527877e-08 2.91904231e-07 1.19527891e-08 2.92004231e-07 1.19527876e-08 2.92104231e-07 1.19527892e-08 2.92204231e-07 1.19527876e-08
+ 2.92304231e-07 1.19527892e-08 2.92404231e-07 1.19527877e-08 2.92504231e-07 1.19527892e-08 2.92604231e-07 1.19527878e-08 2.92704231e-07 1.1952789e-08 2.92804231e-07 1.19527879e-08 2.92904231e-07 1.19527892e-08 2.93004231e-07 1.19527877e-08
+ 2.93104231e-07 1.1952789e-08 2.93204231e-07 1.19527879e-08 2.93304231e-07 1.19527887e-08 2.93404231e-07 1.19527881e-08 2.93504231e-07 1.19527889e-08 2.93604231e-07 1.19527881e-08 2.93704231e-07 1.19527886e-08 2.93804231e-07 1.1952788e-08
+ 2.93904231e-07 1.19527889e-08 2.94004231e-07 1.19527882e-08 2.94104231e-07 1.19527888e-08 2.94204231e-07 1.19527882e-08 2.94304231e-07 1.19527886e-08 2.94404231e-07 1.19527884e-08 2.94504231e-07 1.19527883e-08 2.94604231e-07 1.19527884e-08
+ 2.94704231e-07 1.19527883e-08 2.94804231e-07 1.19527884e-08 2.94904231e-07 1.19527884e-08 2.95004231e-07 1.19527883e-08 2.95104231e-07 1.19527884e-08 2.95204231e-07 1.19527885e-08 2.95304231e-07 1.19527884e-08 2.95404231e-07 1.19527885e-08
+ 2.95504231e-07 1.19527884e-08 2.95604231e-07 1.19527886e-08 2.95704231e-07 1.19527884e-08 2.95804231e-07 1.19527886e-08 2.95904231e-07 1.19527884e-08 2.96004231e-07 1.19527886e-08 2.96104231e-07 1.19527884e-08 2.96204231e-07 1.19527884e-08
+ 2.96304231e-07 1.19527883e-08 2.96404231e-07 1.19527887e-08 2.96504231e-07 1.19527883e-08 2.96604231e-07 1.19527887e-08 2.96704231e-07 1.19527885e-08 2.96804231e-07 1.19527885e-08 2.96904231e-07 1.19527884e-08 2.97004231e-07 1.19527885e-08
+ 2.97104231e-07 1.19527885e-08 2.97204231e-07 1.19527885e-08 2.97304231e-07 1.19527885e-08 2.97404231e-07 1.19527885e-08 2.97504231e-07 1.19527884e-08 2.97604231e-07 1.19527886e-08 2.97704231e-07 1.19527885e-08 2.97804231e-07 1.19527884e-08
+ 2.97904231e-07 1.19527884e-08 2.98004231e-07 1.19527885e-08 2.98104231e-07 1.19527881e-08 2.98204231e-07 1.19527885e-08 2.98304231e-07 1.19527882e-08 2.98404231e-07 1.19527885e-08 2.98504231e-07 1.19527883e-08 2.98604231e-07 1.19527885e-08
+ 2.98704231e-07 1.19527884e-08 2.98804231e-07 1.19527884e-08 2.98904231e-07 1.19527883e-08 2.99004231e-07 1.19527885e-08 2.99104231e-07 1.19527885e-08 2.99204231e-07 1.19527883e-08 2.99304231e-07 1.19527885e-08 2.99404231e-07 1.19527885e-08
+ 2.99504231e-07 1.19527884e-08 2.99604231e-07 1.19527884e-08 2.99704231e-07 1.19527885e-08 2.99804231e-07 1.19527884e-08 2.99904231e-07 1.19527884e-08 3e-07 1.19527883e-08 3.0001e-07 1.19885671e-08 3.0003e-07 1.17808827e-08
+ 3.0007e-07 1.22180336e-08 3.0015e-07 1.1655688e-08 3.0025e-07 1.22568031e-08 3.0035e-07 1.16606775e-08 3.0045e-07 1.22151902e-08 3.0055e-07 1.17418278e-08 3.0065e-07 1.18107334e-08 3.0075e-07 2.87697417e-08
+ 3.0085e-07 -5.432075e-07 3.00931988e-07 7.32055252e-06 3.01e-07 -4.5908469e-05 3.01008484e-07 -5.04559152e-05 3.01025451e-07 -3.69618015e-05 3.01059385e-07 -3.09903885e-05 3.01090588e-07 0.000242070373 3.01143428e-07 0.000483109234
+ 3.011991e-07 0.00152689372 3.012991e-07 -0.0155867066 3.013991e-07 0.117270425 3.014991e-07 4.30152836 3.01578678e-07 5.13555996 3.01663998e-07 4.92548528 3.01763998e-07 5.04581425 3.01858547e-07 4.97061047
+ 3.01958547e-07 5.01945309 3.02058547e-07 4.98680161 3.02158547e-07 5.00891418 3.02258547e-07 4.99390118 3.02358547e-07 5.00413809 3.02458547e-07 4.99716775 3.02558547e-07 5.00191851 3.02658547e-07 4.99869244
+ 3.02758547e-07 5.00087968 3.02858547e-07 4.99940653 3.02958547e-07 5.00039318 3.03058547e-07 4.99974055 3.03158547e-07 5.0001661 3.03258547e-07 4.9998959 3.03358547e-07 5.00006105 3.03458547e-07 4.99996722
+ 3.03558547e-07 5.00001337 3.03658547e-07 4.99999907 3.03758547e-07 4.99999272 3.03858547e-07 5.00001245 3.03958547e-07 4.99998442 3.04058547e-07 5.00001725 3.04158547e-07 4.99998194 3.04258547e-07 5.00001816
+ 3.04358547e-07 4.99998204 3.04458547e-07 5.00001738 3.04558547e-07 4.99998323 3.04658547e-07 5.00001594 3.04758547e-07 4.9999848 3.04858547e-07 5.00001432 3.04958547e-07 4.99998643 3.05058547e-07 5.00001272
+ 3.05158547e-07 4.99998798 3.05258547e-07 5.00001123 3.05358547e-07 4.9999894 3.05458547e-07 5.00000988 3.05558547e-07 4.99999068 3.05658547e-07 5.00000868 3.05758547e-07 4.99999181 3.05858547e-07 5.00000762
+ 3.05958547e-07 4.99999281 3.06058547e-07 5.00000668 3.06158547e-07 4.99999369 3.06258547e-07 5.00000585 3.06358547e-07 4.99999446 3.06458547e-07 5.00000513 3.06558547e-07 4.99999514 3.06658547e-07 5.00000449
+ 3.06758547e-07 4.99999573 3.06858547e-07 5.00000394 3.06958547e-07 4.99999626 3.07058547e-07 5.00000345 3.07158547e-07 4.99999671 3.07258547e-07 5.00000302 3.07358547e-07 4.99999712 3.07458547e-07 5.00000264
+ 3.07558547e-07 4.99999747 3.07658547e-07 5.00000231 3.07758547e-07 4.99999778 3.07858547e-07 5.00000203 3.07958547e-07 4.99999805 3.08058547e-07 5.00000177 3.08158547e-07 4.99999828 3.08258547e-07 5.00000155
+ 3.08358547e-07 4.99999849 3.08458547e-07 5.00000136 3.08558547e-07 4.99999868 3.08658547e-07 5.00000119 3.08758547e-07 4.99999884 3.08858547e-07 5.00000104 3.08958547e-07 4.99999898 3.09058547e-07 5.0000009
+ 3.09158547e-07 4.9999991 3.09258547e-07 5.00000079 3.09358547e-07 4.99999921 3.09458547e-07 5.00000069 3.09558547e-07 4.9999993 3.09658547e-07 5.0000006 3.09758547e-07 4.99999938 3.09858547e-07 5.00000052
+ 3.09958547e-07 4.99999946 3.10058547e-07 5.00000045 3.10158547e-07 4.99999952 3.10258547e-07 5.0000004 3.10358547e-07 4.99999958 3.10458547e-07 5.00000034 3.10558547e-07 4.99999962 3.10658547e-07 5.0000003
+ 3.10758547e-07 4.99999967 3.10858547e-07 5.00000026 3.10958547e-07 4.99999971 3.11058547e-07 5.00000022 3.11158547e-07 4.99999973 3.11258547e-07 5.00000019 3.11358547e-07 4.99999976 3.11458547e-07 5.00000016
+ 3.11558547e-07 4.99999979 3.11658547e-07 5.00000014 3.11758547e-07 4.99999981 3.11858547e-07 5.00000012 3.11958547e-07 4.99999983 3.12058547e-07 5.0000001 3.12158547e-07 4.99999985 3.12258547e-07 5.00000008
+ 3.12358547e-07 4.99999986 3.12458547e-07 5.00000007 3.12558547e-07 4.99999988 3.12658547e-07 5.00000006 3.12758547e-07 4.99999989 3.12858547e-07 5.00000005 3.12958547e-07 4.9999999 3.13058547e-07 5.00000004
+ 3.13158547e-07 4.99999991 3.13258547e-07 5.00000003 3.13358547e-07 4.99999992 3.13458547e-07 5.00000002 3.13558547e-07 4.99999992 3.13658547e-07 5.00000002 3.13758547e-07 4.99999993 3.13858547e-07 5.00000001
+ 3.13958547e-07 4.99999994 3.14058547e-07 5.0 3.14158547e-07 4.99999994 3.14258547e-07 5.0 3.14358547e-07 4.99999994 3.14458547e-07 5.0 3.14558547e-07 4.99999995 3.14658547e-07 4.99999999
+ 3.14758547e-07 4.99999995 3.14858547e-07 4.99999999 3.14958547e-07 4.99999995 3.15058547e-07 4.99999999 3.15158547e-07 4.99999996 3.15258547e-07 4.99999999 3.15358547e-07 4.99999996 3.15458547e-07 4.99999998
+ 3.15558547e-07 4.99999996 3.15658547e-07 4.99999998 3.15758547e-07 4.99999996 3.15858547e-07 4.99999998 3.15958547e-07 4.99999996 3.16058547e-07 4.99999998 3.16158547e-07 4.99999996 3.16258547e-07 4.99999998
+ 3.16358547e-07 4.99999997 3.16458547e-07 4.99999998 3.16558547e-07 4.99999997 3.16658547e-07 4.99999998 3.16758547e-07 4.99999997 3.16858547e-07 4.99999998 3.16958547e-07 4.99999997 3.17058547e-07 4.99999998
+ 3.17158547e-07 4.99999997 3.17258547e-07 4.99999998 3.17358547e-07 4.99999997 3.17458547e-07 4.99999998 3.17558547e-07 4.99999997 3.17658547e-07 4.99999998 3.17758547e-07 4.99999997 3.17858547e-07 4.99999997
+ 3.17958547e-07 4.99999997 3.18058547e-07 4.99999997 3.18158547e-07 4.99999997 3.18258547e-07 4.99999997 3.18358547e-07 4.99999997 3.18458547e-07 4.99999997 3.18558547e-07 4.99999997 3.18658547e-07 4.99999997
+ 3.18758547e-07 4.99999997 3.18858547e-07 4.99999997 3.18958547e-07 4.99999997 3.19058547e-07 4.99999997 3.19158547e-07 4.99999997 3.19258547e-07 4.99999997 3.19358547e-07 4.99999997 3.19458547e-07 4.99999997
+ 3.19558547e-07 4.99999997 3.19658547e-07 4.99999997 3.19758547e-07 4.99999997 3.19858547e-07 4.99999997 3.19958547e-07 4.99999997 3.20058547e-07 4.99999997 3.20158547e-07 4.99999997 3.20258547e-07 4.99999997
+ 3.20358547e-07 4.99999997 3.20458547e-07 4.99999997 3.20558547e-07 4.99999997 3.20658547e-07 4.99999997 3.20758547e-07 4.99999997 3.20858547e-07 4.99999997 3.20958547e-07 4.99999997 3.21058547e-07 4.99999997
+ 3.21158547e-07 4.99999997 3.21258547e-07 4.99999997 3.21358547e-07 4.99999997 3.21458547e-07 4.99999997 3.21558547e-07 4.99999997 3.21658547e-07 4.99999997 3.21758547e-07 4.99999997 3.21858547e-07 4.99999997
+ 3.21958547e-07 4.99999997 3.22058547e-07 4.99999997 3.22158547e-07 4.99999997 3.22258547e-07 4.99999997 3.22358547e-07 4.99999997 3.22458547e-07 4.99999997 3.22558547e-07 4.99999997 3.22658547e-07 4.99999997
+ 3.22758547e-07 4.99999997 3.22858547e-07 4.99999997 3.22958547e-07 4.99999997 3.23058547e-07 4.99999997 3.23158547e-07 4.99999997 3.23258547e-07 4.99999997 3.23358547e-07 4.99999997 3.23458547e-07 4.99999997
+ 3.23558547e-07 4.99999997 3.23658547e-07 4.99999997 3.23758547e-07 4.99999997 3.23858547e-07 4.99999997 3.23958547e-07 4.99999997 3.24058547e-07 4.99999997 3.24158547e-07 4.99999997 3.24258547e-07 4.99999997
+ 3.24358547e-07 4.99999997 3.24458547e-07 4.99999997 3.24558547e-07 4.99999997 3.24658547e-07 4.99999997 3.24758547e-07 4.99999997 3.24858547e-07 4.99999997 3.24958547e-07 4.99999997 3.25058547e-07 4.99999997
+ 3.25158547e-07 4.99999997 3.25258547e-07 4.99999997 3.25358547e-07 4.99999997 3.25458547e-07 4.99999997 3.25558547e-07 4.99999997 3.25658547e-07 4.99999997 3.25758547e-07 4.99999997 3.25858547e-07 4.99999997
+ 3.25958547e-07 4.99999997 3.26058547e-07 4.99999997 3.26158547e-07 4.99999997 3.26258547e-07 4.99999997 3.26358547e-07 4.99999997 3.26458547e-07 4.99999997 3.26558547e-07 4.99999997 3.26658547e-07 4.99999997
+ 3.26758547e-07 4.99999997 3.26858547e-07 4.99999997 3.26958547e-07 4.99999997 3.27058547e-07 4.99999997 3.27158547e-07 4.99999997 3.27258547e-07 4.99999997 3.27358547e-07 4.99999997 3.27458547e-07 4.99999997
+ 3.27558547e-07 4.99999997 3.27658547e-07 4.99999997 3.27758547e-07 4.99999997 3.27858547e-07 4.99999997 3.27958547e-07 4.99999997 3.28058547e-07 4.99999997 3.28158547e-07 4.99999997 3.28258547e-07 4.99999997
+ 3.28358547e-07 4.99999997 3.28458547e-07 4.99999997 3.28558547e-07 4.99999997 3.28658547e-07 4.99999997 3.28758547e-07 4.99999997 3.28858547e-07 4.99999997 3.28958547e-07 4.99999997 3.29058547e-07 4.99999997
+ 3.29158547e-07 4.99999997 3.29258547e-07 4.99999997 3.29358547e-07 4.99999997 3.29458547e-07 4.99999997 3.29558547e-07 4.99999997 3.29658547e-07 4.99999997 3.29758547e-07 4.99999997 3.29858547e-07 4.99999997
+ 3.29958547e-07 4.99999997 3.30058547e-07 4.99999997 3.30158547e-07 4.99999997 3.30258547e-07 4.99999997 3.30358547e-07 4.99999997 3.30458547e-07 4.99999997 3.30558547e-07 4.99999997 3.30658547e-07 4.99999997
+ 3.30758547e-07 4.99999997 3.30858547e-07 4.99999997 3.30958547e-07 4.99999997 3.31058547e-07 4.99999997 3.31158547e-07 4.99999997 3.31258547e-07 4.99999997 3.31358547e-07 4.99999997 3.31458547e-07 4.99999997
+ 3.31558547e-07 4.99999997 3.31658547e-07 4.99999997 3.31758547e-07 4.99999997 3.31858547e-07 4.99999997 3.31958547e-07 4.99999997 3.32058547e-07 4.99999997 3.32158547e-07 4.99999997 3.32258547e-07 4.99999997
+ 3.32358547e-07 4.99999997 3.32458547e-07 4.99999997 3.32558547e-07 4.99999997 3.32658547e-07 4.99999997 3.32758547e-07 4.99999997 3.32858547e-07 4.99999997 3.32958547e-07 4.99999997 3.33058547e-07 4.99999997
+ 3.33158547e-07 4.99999997 3.33258547e-07 4.99999997 3.33358547e-07 4.99999997 3.33458547e-07 4.99999997 3.33558547e-07 4.99999997 3.33658547e-07 4.99999997 3.33758547e-07 4.99999997 3.33858547e-07 4.99999997
+ 3.33958547e-07 4.99999997 3.34058547e-07 4.99999997 3.34158547e-07 4.99999997 3.34258547e-07 4.99999997 3.34358547e-07 4.99999997 3.34458547e-07 4.99999997 3.34558547e-07 4.99999997 3.34658547e-07 4.99999997
+ 3.34758547e-07 4.99999997 3.34858547e-07 4.99999997 3.34958547e-07 4.99999997 3.35058547e-07 4.99999997 3.35158547e-07 4.99999997 3.35258547e-07 4.99999997 3.35358547e-07 4.99999997 3.35458547e-07 4.99999997
+ 3.35558547e-07 4.99999997 3.35658547e-07 4.99999997 3.35758547e-07 4.99999997 3.35858547e-07 4.99999997 3.35958547e-07 4.99999997 3.36058547e-07 4.99999997 3.36158547e-07 4.99999997 3.36258547e-07 4.99999997
+ 3.36358547e-07 4.99999997 3.36458547e-07 4.99999997 3.36558547e-07 4.99999997 3.36658547e-07 4.99999997 3.36758547e-07 4.99999997 3.36858547e-07 4.99999997 3.36958547e-07 4.99999997 3.37058547e-07 4.99999997
+ 3.37158547e-07 4.99999997 3.37258547e-07 4.99999997 3.37358547e-07 4.99999997 3.37458547e-07 4.99999997 3.37558547e-07 4.99999997 3.37658547e-07 4.99999997 3.37758547e-07 4.99999997 3.37858547e-07 4.99999997
+ 3.37958547e-07 4.99999997 3.38058547e-07 4.99999997 3.38158547e-07 4.99999997 3.38258547e-07 4.99999997 3.38358547e-07 4.99999997 3.38458547e-07 4.99999997 3.38558547e-07 4.99999997 3.38658547e-07 4.99999997
+ 3.38758547e-07 4.99999997 3.38858547e-07 4.99999997 3.38958547e-07 4.99999997 3.39058547e-07 4.99999997 3.39158547e-07 4.99999997 3.39258547e-07 4.99999997 3.39358547e-07 4.99999997 3.39458547e-07 4.99999997
+ 3.39558547e-07 4.99999997 3.39658547e-07 4.99999997 3.39758547e-07 4.99999997 3.39858547e-07 4.99999997 3.39958547e-07 4.99999997 3.40058547e-07 4.99999997 3.40158547e-07 4.99999997 3.40258547e-07 4.99999997
+ 3.40358547e-07 4.99999997 3.40458547e-07 4.99999997 3.40558547e-07 4.99999997 3.40658547e-07 4.99999997 3.40758547e-07 4.99999997 3.40858547e-07 4.99999997 3.40958547e-07 4.99999997 3.41058547e-07 4.99999997
+ 3.41158547e-07 4.99999997 3.41258547e-07 4.99999997 3.41358547e-07 4.99999997 3.41458547e-07 4.99999997 3.41558547e-07 4.99999997 3.41658547e-07 4.99999997 3.41758547e-07 4.99999997 3.41858547e-07 4.99999997
+ 3.41958547e-07 4.99999997 3.42058547e-07 4.99999997 3.42158547e-07 4.99999997 3.42258547e-07 4.99999997 3.42358547e-07 4.99999997 3.42458547e-07 4.99999997 3.42558547e-07 4.99999997 3.42658547e-07 4.99999997
+ 3.42758547e-07 4.99999997 3.42858547e-07 4.99999997 3.42958547e-07 4.99999997 3.43058547e-07 4.99999997 3.43158547e-07 4.99999997 3.43258547e-07 4.99999997 3.43358547e-07 4.99999997 3.43458547e-07 4.99999997
+ 3.43558547e-07 4.99999997 3.43658547e-07 4.99999997 3.43758547e-07 4.99999997 3.43858547e-07 4.99999997 3.43958547e-07 4.99999997 3.44058547e-07 4.99999997 3.44158547e-07 4.99999997 3.44258547e-07 4.99999997
+ 3.44358547e-07 4.99999997 3.44458547e-07 4.99999997 3.44558547e-07 4.99999997 3.44658547e-07 4.99999997 3.44758547e-07 4.99999997 3.44858547e-07 4.99999997 3.44958547e-07 4.99999997 3.45058547e-07 4.99999997
+ 3.45158547e-07 4.99999997 3.45258547e-07 4.99999997 3.45358547e-07 4.99999997 3.45458547e-07 4.99999997 3.45558547e-07 4.99999997 3.45658547e-07 4.99999997 3.45758547e-07 4.99999997 3.45858547e-07 4.99999997
+ 3.45958547e-07 4.99999997 3.46058547e-07 4.99999997 3.46158547e-07 4.99999997 3.46258547e-07 4.99999997 3.46358547e-07 4.99999997 3.46458547e-07 4.99999997 3.46558547e-07 4.99999997 3.46658547e-07 4.99999997
+ 3.46758547e-07 4.99999997 3.46858547e-07 4.99999997 3.46958547e-07 4.99999997 3.47058547e-07 4.99999997 3.47158547e-07 4.99999997 3.47258547e-07 4.99999997 3.47358547e-07 4.99999997 3.47458547e-07 4.99999997
+ 3.47558547e-07 4.99999997 3.47658547e-07 4.99999997 3.47758547e-07 4.99999997 3.47858547e-07 4.99999997 3.47958547e-07 4.99999997 3.48058547e-07 4.99999997 3.48158547e-07 4.99999997 3.48258547e-07 4.99999997
+ 3.48358547e-07 4.99999997 3.48458547e-07 4.99999997 3.48558547e-07 4.99999997 3.48658547e-07 4.99999997 3.48758547e-07 4.99999997 3.48858547e-07 4.99999997 3.48958547e-07 4.99999997 3.49058547e-07 4.99999997
+ 3.49158547e-07 4.99999997 3.49258547e-07 4.99999997 3.49358547e-07 4.99999997 3.49458547e-07 4.99999997 3.49558547e-07 4.99999997 3.49658547e-07 4.99999997 3.49758547e-07 4.99999997 3.49858547e-07 4.99999997
+ 3.49958547e-07 4.99999997 3.50058547e-07 4.99999997 3.50158547e-07 4.99999997 3.50258547e-07 4.99999997 3.50358547e-07 4.99999997 3.50458547e-07 4.99999997 3.50558547e-07 4.99999997 3.50658547e-07 4.99999997
+ 3.50758547e-07 4.99999997 3.50858547e-07 4.99999997 3.50958547e-07 4.99999997 3.51e-07 4.99999997 3.5101e-07 4.99999997 3.5103e-07 4.99999997 3.5107e-07 4.99999997 3.5115e-07 4.99999997
+ 3.5125e-07 4.99999997 3.5135e-07 4.99999997 3.5145e-07 4.99999997 3.5155e-07 4.99999997 3.5165e-07 4.99999997 3.5175e-07 4.99999997 3.5185e-07 4.99999997 3.51930828e-07 5.00000066
+ 3.52e-07 5.00000151 3.52008608e-07 4.9999927 3.52025825e-07 4.99997482 3.52060258e-07 4.99999285 3.52106188e-07 5.00004461 3.52150118e-07 5.00000795 3.5219811e-07 4.99994547 3.522555e-07 5.00002987
+ 3.52312176e-07 4.9999935 3.52404431e-07 5.0000036 3.52490759e-07 4.99999971 3.52590759e-07 4.99999801 3.52690759e-07 5.00000291 3.52790759e-07 4.99999668 3.52890759e-07 5.00000318 3.52990759e-07 4.99999704
+ 3.53090759e-07 5.00000252 3.53190759e-07 4.99999781 3.53290759e-07 5.00000177 3.53390759e-07 4.9999985 3.53490759e-07 5.00000116 3.53590759e-07 4.99999902 3.53690759e-07 5.00000073 3.53790759e-07 4.99999937
+ 3.53890759e-07 5.00000045 3.53990759e-07 4.99999959 3.54090759e-07 5.00000027 3.54190759e-07 4.99999973 3.54290759e-07 5.00000017 3.54390759e-07 4.99999981 3.54490759e-07 5.0000001 3.54590759e-07 4.99999986
+ 3.54690759e-07 5.00000006 3.54790759e-07 4.99999989 3.54890759e-07 5.00000004 3.54990759e-07 4.99999991 3.55090759e-07 5.00000002 3.55190759e-07 4.99999992 3.55290759e-07 5.00000002 3.55390759e-07 4.99999993
+ 3.55490759e-07 5.00000001 3.55590759e-07 4.99999994 3.55690759e-07 5.0 3.55790759e-07 4.99999994 3.55890759e-07 5.0 3.55990759e-07 4.99999994 3.56090759e-07 5.0 3.56190759e-07 4.99999995
+ 3.56290759e-07 5.0 3.56390759e-07 4.99999995 3.56490759e-07 4.99999999 3.56590759e-07 4.99999995 3.56690759e-07 4.99999999 3.56790759e-07 4.99999995 3.56890759e-07 4.99999999 3.56990759e-07 4.99999995
+ 3.57090759e-07 4.99999999 3.57190759e-07 4.99999996 3.57290759e-07 4.99999999 3.57390759e-07 4.99999996 3.57490759e-07 4.99999999 3.57590759e-07 4.99999996 3.57690759e-07 4.99999998 3.57790759e-07 4.99999996
+ 3.57890759e-07 4.99999998 3.57990759e-07 4.99999996 3.58090759e-07 4.99999998 3.58190759e-07 4.99999996 3.58290759e-07 4.99999998 3.58390759e-07 4.99999996 3.58490759e-07 4.99999998 3.58590759e-07 4.99999997
+ 3.58690759e-07 4.99999998 3.58790759e-07 4.99999997 3.58890759e-07 4.99999998 3.58990759e-07 4.99999997 3.59090759e-07 4.99999998 3.59190759e-07 4.99999997 3.59290759e-07 4.99999998 3.59390759e-07 4.99999997
+ 3.59490759e-07 4.99999998 3.59590759e-07 4.99999997 3.59690759e-07 4.99999998 3.59790759e-07 4.99999997 3.59890759e-07 4.99999998 3.59990759e-07 4.99999997 3.60090759e-07 4.99999997 3.60190759e-07 4.99999997
+ 3.60290759e-07 4.99999997 3.60390759e-07 4.99999997 3.60490759e-07 4.99999997 3.60590759e-07 4.99999997 3.60690759e-07 4.99999997 3.60790759e-07 4.99999997 3.60890759e-07 4.99999997 3.60990759e-07 4.99999997
+ 3.61090759e-07 4.99999997 3.61190759e-07 4.99999997 3.61290759e-07 4.99999997 3.61390759e-07 4.99999997 3.61490759e-07 4.99999997 3.61590759e-07 4.99999997 3.61690759e-07 4.99999997 3.61790759e-07 4.99999997
+ 3.61890759e-07 4.99999997 3.61990759e-07 4.99999997 3.62090759e-07 4.99999997 3.62190759e-07 4.99999997 3.62290759e-07 4.99999997 3.62390759e-07 4.99999997 3.62490759e-07 4.99999997 3.62590759e-07 4.99999997
+ 3.62690759e-07 4.99999997 3.62790759e-07 4.99999997 3.62890759e-07 4.99999997 3.62990759e-07 4.99999997 3.63090759e-07 4.99999997 3.63190759e-07 4.99999997 3.63290759e-07 4.99999997 3.63390759e-07 4.99999997
+ 3.63490759e-07 4.99999997 3.63590759e-07 4.99999997 3.63690759e-07 4.99999997 3.63790759e-07 4.99999997 3.63890759e-07 4.99999997 3.63990759e-07 4.99999997 3.64090759e-07 4.99999997 3.64190759e-07 4.99999997
+ 3.64290759e-07 4.99999997 3.64390759e-07 4.99999997 3.64490759e-07 4.99999997 3.64590759e-07 4.99999997 3.64690759e-07 4.99999997 3.64790759e-07 4.99999997 3.64890759e-07 4.99999997 3.64990759e-07 4.99999997
+ 3.65090759e-07 4.99999997 3.65190759e-07 4.99999997 3.65290759e-07 4.99999997 3.65390759e-07 4.99999997 3.65490759e-07 4.99999997 3.65590759e-07 4.99999997 3.65690759e-07 4.99999997 3.65790759e-07 4.99999997
+ 3.65890759e-07 4.99999997 3.65990759e-07 4.99999997 3.66090759e-07 4.99999997 3.66190759e-07 4.99999997 3.66290759e-07 4.99999997 3.66390759e-07 4.99999997 3.66490759e-07 4.99999997 3.66590759e-07 4.99999997
+ 3.66690759e-07 4.99999997 3.66790759e-07 4.99999997 3.66890759e-07 4.99999997 3.66990759e-07 4.99999997 3.67090759e-07 4.99999997 3.67190759e-07 4.99999997 3.67290759e-07 4.99999997 3.67390759e-07 4.99999997
+ 3.67490759e-07 4.99999997 3.67590759e-07 4.99999997 3.67690759e-07 4.99999997 3.67790759e-07 4.99999997 3.67890759e-07 4.99999997 3.67990759e-07 4.99999997 3.68090759e-07 4.99999997 3.68190759e-07 4.99999997
+ 3.68290759e-07 4.99999997 3.68390759e-07 4.99999997 3.68490759e-07 4.99999997 3.68590759e-07 4.99999997 3.68690759e-07 4.99999997 3.68790759e-07 4.99999997 3.68890759e-07 4.99999997 3.68990759e-07 4.99999997
+ 3.69090759e-07 4.99999997 3.69190759e-07 4.99999997 3.69290759e-07 4.99999997 3.69390759e-07 4.99999997 3.69490759e-07 4.99999997 3.69590759e-07 4.99999997 3.69690759e-07 4.99999997 3.69790759e-07 4.99999997
+ 3.69890759e-07 4.99999997 3.69990759e-07 4.99999997 3.70090759e-07 4.99999997 3.70190759e-07 4.99999997 3.70290759e-07 4.99999997 3.70390759e-07 4.99999997 3.70490759e-07 4.99999997 3.70590759e-07 4.99999997
+ 3.70690759e-07 4.99999997 3.70790759e-07 4.99999997 3.70890759e-07 4.99999997 3.70990759e-07 4.99999997 3.71090759e-07 4.99999997 3.71190759e-07 4.99999997 3.71290759e-07 4.99999997 3.71390759e-07 4.99999997
+ 3.71490759e-07 4.99999997 3.71590759e-07 4.99999997 3.71690759e-07 4.99999997 3.71790759e-07 4.99999997 3.71890759e-07 4.99999997 3.71990759e-07 4.99999997 3.72090759e-07 4.99999997 3.72190759e-07 4.99999997
+ 3.72290759e-07 4.99999997 3.72390759e-07 4.99999997 3.72490759e-07 4.99999997 3.72590759e-07 4.99999997 3.72690759e-07 4.99999997 3.72790759e-07 4.99999997 3.72890759e-07 4.99999997 3.72990759e-07 4.99999997
+ 3.73090759e-07 4.99999997 3.73190759e-07 4.99999997 3.73290759e-07 4.99999997 3.73390759e-07 4.99999997 3.73490759e-07 4.99999997 3.73590759e-07 4.99999997 3.73690759e-07 4.99999997 3.73790759e-07 4.99999997
+ 3.73890759e-07 4.99999997 3.73990759e-07 4.99999997 3.74090759e-07 4.99999997 3.74190759e-07 4.99999997 3.74290759e-07 4.99999997 3.74390759e-07 4.99999997 3.74490759e-07 4.99999997 3.74590759e-07 4.99999997
+ 3.74690759e-07 4.99999997 3.74790759e-07 4.99999997 3.74890759e-07 4.99999997 3.74990759e-07 4.99999997 3.75090759e-07 4.99999997 3.75190759e-07 4.99999997 3.75290759e-07 4.99999997 3.75390759e-07 4.99999997
+ 3.75490759e-07 4.99999997 3.75590759e-07 4.99999997 3.75690759e-07 4.99999997 3.75790759e-07 4.99999997 3.75890759e-07 4.99999997 3.75990759e-07 4.99999997 3.76090759e-07 4.99999997 3.76190759e-07 4.99999997
+ 3.76290759e-07 4.99999997 3.76390759e-07 4.99999997 3.76490759e-07 4.99999997 3.76590759e-07 4.99999997 3.76690759e-07 4.99999997 3.76790759e-07 4.99999997 3.76890759e-07 4.99999997 3.76990759e-07 4.99999997
+ 3.77090759e-07 4.99999997 3.77190759e-07 4.99999997 3.77290759e-07 4.99999997 3.77390759e-07 4.99999997 3.77490759e-07 4.99999997 3.77590759e-07 4.99999997 3.77690759e-07 4.99999997 3.77790759e-07 4.99999997
+ 3.77890759e-07 4.99999997 3.77990759e-07 4.99999997 3.78090759e-07 4.99999997 3.78190759e-07 4.99999997 3.78290759e-07 4.99999997 3.78390759e-07 4.99999997 3.78490759e-07 4.99999997 3.78590759e-07 4.99999997
+ 3.78690759e-07 4.99999997 3.78790759e-07 4.99999997 3.78890759e-07 4.99999997 3.78990759e-07 4.99999997 3.79090759e-07 4.99999997 3.79190759e-07 4.99999997 3.79290759e-07 4.99999997 3.79390759e-07 4.99999997
+ 3.79490759e-07 4.99999997 3.79590759e-07 4.99999997 3.79690759e-07 4.99999997 3.79790759e-07 4.99999997 3.79890759e-07 4.99999997 3.79990759e-07 4.99999997 3.80090759e-07 4.99999997 3.80190759e-07 4.99999997
+ 3.80290759e-07 4.99999997 3.80390759e-07 4.99999997 3.80490759e-07 4.99999997 3.80590759e-07 4.99999997 3.80690759e-07 4.99999997 3.80790759e-07 4.99999997 3.80890759e-07 4.99999997 3.80990759e-07 4.99999997
+ 3.81090759e-07 4.99999997 3.81190759e-07 4.99999997 3.81290759e-07 4.99999997 3.81390759e-07 4.99999997 3.81490759e-07 4.99999997 3.81590759e-07 4.99999997 3.81690759e-07 4.99999997 3.81790759e-07 4.99999997
+ 3.81890759e-07 4.99999997 3.81990759e-07 4.99999997 3.82090759e-07 4.99999997 3.82190759e-07 4.99999997 3.82290759e-07 4.99999997 3.82390759e-07 4.99999997 3.82490759e-07 4.99999997 3.82590759e-07 4.99999997
+ 3.82690759e-07 4.99999997 3.82790759e-07 4.99999997 3.82890759e-07 4.99999997 3.82990759e-07 4.99999997 3.83090759e-07 4.99999997 3.83190759e-07 4.99999997 3.83290759e-07 4.99999997 3.83390759e-07 4.99999997
+ 3.83490759e-07 4.99999997 3.83590759e-07 4.99999997 3.83690759e-07 4.99999997 3.83790759e-07 4.99999997 3.83890759e-07 4.99999997 3.83990759e-07 4.99999997 3.84090759e-07 4.99999997 3.84190759e-07 4.99999997
+ 3.84290759e-07 4.99999997 3.84390759e-07 4.99999997 3.84490759e-07 4.99999997 3.84590759e-07 4.99999997 3.84690759e-07 4.99999997 3.84790759e-07 4.99999997 3.84890759e-07 4.99999997 3.84990759e-07 4.99999997
+ 3.85090759e-07 4.99999997 3.85190759e-07 4.99999997 3.85290759e-07 4.99999997 3.85390759e-07 4.99999997 3.85490759e-07 4.99999997 3.85590759e-07 4.99999997 3.85690759e-07 4.99999997 3.85790759e-07 4.99999997
+ 3.85890759e-07 4.99999997 3.85990759e-07 4.99999997 3.86090759e-07 4.99999997 3.86190759e-07 4.99999997 3.86290759e-07 4.99999997 3.86390759e-07 4.99999997 3.86490759e-07 4.99999997 3.86590759e-07 4.99999997
+ 3.86690759e-07 4.99999997 3.86790759e-07 4.99999997 3.86890759e-07 4.99999997 3.86990759e-07 4.99999997 3.87090759e-07 4.99999997 3.87190759e-07 4.99999997 3.87290759e-07 4.99999997 3.87390759e-07 4.99999997
+ 3.87490759e-07 4.99999997 3.87590759e-07 4.99999997 3.87690759e-07 4.99999997 3.87790759e-07 4.99999997 3.87890759e-07 4.99999997 3.87990759e-07 4.99999997 3.88090759e-07 4.99999997 3.88190759e-07 4.99999997
+ 3.88290759e-07 4.99999997 3.88390759e-07 4.99999997 3.88490759e-07 4.99999997 3.88590759e-07 4.99999997 3.88690759e-07 4.99999997 3.88790759e-07 4.99999997 3.88890759e-07 4.99999997 3.88990759e-07 4.99999997
+ 3.89090759e-07 4.99999997 3.89190759e-07 4.99999997 3.89290759e-07 4.99999997 3.89390759e-07 4.99999997 3.89490759e-07 4.99999997 3.89590759e-07 4.99999997 3.89690759e-07 4.99999997 3.89790759e-07 4.99999997
+ 3.89890759e-07 4.99999997 3.89990759e-07 4.99999997 3.90090759e-07 4.99999997 3.90190759e-07 4.99999997 3.90290759e-07 4.99999997 3.90390759e-07 4.99999997 3.90490759e-07 4.99999997 3.90590759e-07 4.99999997
+ 3.90690759e-07 4.99999997 3.90790759e-07 4.99999997 3.90890759e-07 4.99999997 3.90990759e-07 4.99999997 3.91090759e-07 4.99999997 3.91190759e-07 4.99999997 3.91290759e-07 4.99999997 3.91390759e-07 4.99999997
+ 3.91490759e-07 4.99999997 3.91590759e-07 4.99999997 3.91690759e-07 4.99999997 3.91790759e-07 4.99999997 3.91890759e-07 4.99999997 3.91990759e-07 4.99999997 3.92090759e-07 4.99999997 3.92190759e-07 4.99999997
+ 3.92290759e-07 4.99999997 3.92390759e-07 4.99999997 3.92490759e-07 4.99999997 3.92590759e-07 4.99999997 3.92690759e-07 4.99999997 3.92790759e-07 4.99999997 3.92890759e-07 4.99999997 3.92990759e-07 4.99999997
+ 3.93090759e-07 4.99999997 3.93190759e-07 4.99999997 3.93290759e-07 4.99999997 3.93390759e-07 4.99999997 3.93490759e-07 4.99999997 3.93590759e-07 4.99999997 3.93690759e-07 4.99999997 3.93790759e-07 4.99999997
+ 3.93890759e-07 4.99999997 3.93990759e-07 4.99999997 3.94090759e-07 4.99999997 3.94190759e-07 4.99999997 3.94290759e-07 4.99999997 3.94390759e-07 4.99999997 3.94490759e-07 4.99999997 3.94590759e-07 4.99999997
+ 3.94690759e-07 4.99999997 3.94790759e-07 4.99999997 3.94890759e-07 4.99999997 3.94990759e-07 4.99999997 3.95090759e-07 4.99999997 3.95190759e-07 4.99999997 3.95290759e-07 4.99999997 3.95390759e-07 4.99999997
+ 3.95490759e-07 4.99999997 3.95590759e-07 4.99999997 3.95690759e-07 4.99999997 3.95790759e-07 4.99999997 3.95890759e-07 4.99999997 3.95990759e-07 4.99999997 3.96090759e-07 4.99999997 3.96190759e-07 4.99999997
+ 3.96290759e-07 4.99999997 3.96390759e-07 4.99999997 3.96490759e-07 4.99999997 3.96590759e-07 4.99999997 3.96690759e-07 4.99999997 3.96790759e-07 4.99999997 3.96890759e-07 4.99999997 3.96990759e-07 4.99999997
+ 3.97090759e-07 4.99999997 3.97190759e-07 4.99999997 3.97290759e-07 4.99999997 3.97390759e-07 4.99999997 3.97490759e-07 4.99999997 3.97590759e-07 4.99999997 3.97690759e-07 4.99999997 3.97790759e-07 4.99999997
+ 3.97890759e-07 4.99999997 3.97990759e-07 4.99999997 3.98090759e-07 4.99999997 3.98190759e-07 4.99999997 3.98290759e-07 4.99999997 3.98390759e-07 4.99999997 3.98490759e-07 4.99999997 3.98590759e-07 4.99999997
+ 3.98690759e-07 4.99999997 3.98790759e-07 4.99999997 3.98890759e-07 4.99999997 3.98990759e-07 4.99999997 3.99090759e-07 4.99999997 3.99190759e-07 4.99999997 3.99290759e-07 4.99999997 3.99390759e-07 4.99999997
+ 3.99490759e-07 4.99999997 3.99590759e-07 4.99999997 3.99690759e-07 4.99999997 3.99790759e-07 4.99999997 3.99890759e-07 4.99999997 3.99990759e-07 4.99999997 4e-07 4.99999997 4.0001e-07 4.99999997
+ 4.0003e-07 4.99999997 4.0007e-07 4.99999997 4.0015e-07 4.99999997 4.0025e-07 4.99999997 4.0035e-07 4.99999997 4.0045e-07 4.99999997 4.0055e-07 4.99999997 4.0065e-07 4.99999997
+ 4.0075e-07 5.00000001 4.0085e-07 4.99999717 4.00931913e-07 5.00000328 4.01e-07 5.00008601 4.01008477e-07 5.00011635 4.01025432e-07 5.00022698 4.01059342e-07 4.99960029 4.01090545e-07 4.99796703
+ 4.01143412e-07 4.99703072 4.01199108e-07 5.02828621 4.01266691e-07 4.9918975 4.01329415e-07 3.49023986 4.01394829e-07 0.154819829 4.01464618e-07 -0.00376126514 4.01533535e-07 0.0257937047 4.01610366e-07 -0.0174819665
+ 4.01709241e-07 0.0166256226 4.01809241e-07 -0.0151036136 4.01909241e-07 0.0138168911 4.02009241e-07 -0.0125784687 4.02109241e-07 0.011505171 4.02209241e-07 -0.010481817 4.02309241e-07 0.00958739706 4.02409241e-07 -0.00873958877
+ 4.02509241e-07 0.00799375037 4.02609241e-07 -0.00729006223 4.02709241e-07 0.00666768862 4.02809241e-07 -0.00608276976 4.02909241e-07 0.00556317247 4.03009241e-07 -0.00507645127 4.03109241e-07 0.00464253506 4.03209241e-07 -0.00423720493
+ 4.03309241e-07 0.00387478758 4.03409241e-07 -0.00353704076 4.03509241e-07 0.00323432261 4.03609241e-07 -0.00295276769 4.03709241e-07 0.00269991248 4.03809241e-07 -0.00246512287 4.03909241e-07 0.00225392144 4.04009241e-07 -0.00205807943
+ 4.04109241e-07 0.00188167602 4.04209241e-07 -0.00171828798 4.04309241e-07 0.00157095524 4.04409241e-07 -0.00143462118 4.04509241e-07 0.00131157363 4.04609241e-07 -0.00119779915 4.04709241e-07 0.00109503818 4.04809241e-07 -0.00100008016
+ 4.04909241e-07 0.000914264687 4.05009241e-07 -0.000835004145 4.05109241e-07 0.000763342619 4.05209241e-07 -0.00069717962 4.05309241e-07 0.000637339801 4.05409241e-07 -0.000582106412 4.05509241e-07 0.000532139928 4.05609241e-07 -0.000486027981
+ 4.05709241e-07 0.000444307246 4.05809241e-07 -0.000405808347 4.05909241e-07 0.000370973849 4.06009241e-07 -0.000338829481 4.06109241e-07 0.000309745686 4.06209241e-07 -0.000282905677 4.06309241e-07 0.000258624171 4.06409241e-07 -0.000236212099
+ 4.06509241e-07 0.000215940793 4.06609241e-07 -0.000197225188 4.06709241e-07 0.000180302581 4.06809241e-07 -0.000164672908 4.06909241e-07 0.000151581252 4.07009241e-07 -0.000137330071 4.07109241e-07 0.000125617353 4.07209241e-07 -0.000114721651
+ 4.07309241e-07 0.000104886816 4.07409241e-07 -9.57863029e-05 4.07509241e-07 8.75782273e-05 4.07609241e-07 -7.99758898e-05 4.07709241e-07 7.31262283e-05 4.07809241e-07 -6.67747637e-05 4.07909241e-07 6.14617377e-05 4.08009241e-07 -5.56877955e-05
+ 4.08109241e-07 5.12854283e-05 4.08209241e-07 -4.64651204e-05 4.08309241e-07 4.27945085e-05 4.08409241e-07 -3.85326677e-05 4.08509241e-07 3.57459199e-05 4.08609241e-07 -3.21645777e-05 4.08709241e-07 2.98427245e-05 4.08809241e-07 -2.68487335e-05
+ 4.08909241e-07 2.49148683e-05 4.09009241e-07 -2.24112808e-05 4.09109241e-07 2.08011545e-05 4.09209241e-07 -1.87070504e-05 4.09309241e-07 1.73671183e-05 4.09409241e-07 -1.56148482e-05 4.09509241e-07 1.45003217e-05 4.09609241e-07 -1.30334472e-05
+ 4.09709241e-07 1.2107067e-05 4.09809241e-07 -1.08784781e-05 4.09909241e-07 1.01091346e-05 4.10009241e-07 -9.07948871e-06 4.10109241e-07 8.44121874e-06 4.10209241e-07 -7.57766587e-06 4.10309241e-07 7.04880191e-06 4.10409241e-07 -6.3239152e-06
+ 4.10509241e-07 5.8863742e-06 4.10609241e-07 -5.27725522e-06 4.10709241e-07 4.91594507e-06 4.10809241e-07 -4.40347637e-06 4.10909241e-07 4.10580046e-06 4.11009241e-07 -3.67402123e-06 4.11109241e-07 3.42946531e-06 4.11209241e-07 -3.06505021e-06
+ 4.11309241e-07 2.8648379e-06 4.11409241e-07 -2.55666197e-06 4.11509241e-07 2.39346732e-06 4.11609241e-07 -2.13224273e-06 4.11709241e-07 1.99995037e-06 4.11809241e-07 -1.77792302e-06 4.11909241e-07 1.67142791e-06 4.12009241e-07 -1.48212383e-06
+ 4.12109241e-07 1.39716414e-06 4.12209241e-07 -1.23517925e-06 4.12309241e-07 1.16819841e-06 4.12409241e-07 -1.0290213e-06 4.12509241e-07 9.77049652e-07 4.12609241e-07 -8.56913387e-07 4.12709241e-07 8.17471684e-07 4.12809241e-07 -7.13231541e-07
+ 4.12909241e-07 6.84250153e-07 4.13009241e-07 -5.93280523e-07 4.13109241e-07 5.73031515e-07 4.13209241e-07 -4.93140772e-07 4.13309241e-07 4.80181928e-07 4.13409241e-07 -4.09540301e-07 4.13509241e-07 4.026675e-07 4.13609241e-07 -3.39747396e-07
+ 4.13709241e-07 3.37955415e-07 4.13809241e-07 -2.81481545e-07 4.13909241e-07 2.83931201e-07 4.14009241e-07 -2.32838909e-07 4.14109241e-07 2.38829636e-07 4.14209241e-07 -1.92230101e-07 4.14309241e-07 2.01177043e-07 4.14409241e-07 -1.58328245e-07
+ 4.14509241e-07 1.69743148e-07 4.14609241e-07 -1.30025615e-07 4.14709241e-07 1.43500864e-07 4.14809241e-07 -1.06397437e-07 4.14909241e-07 1.21592743e-07 4.15009241e-07 -8.66716733e-08 4.15109241e-07 1.03302951e-07 4.15209241e-07 -7.02059616e-08
+ 4.15309241e-07 8.80380009e-08 4.15409241e-07 -5.64647246e-08 4.15509241e-07 7.53001778e-08 4.15609241e-07 -4.49983215e-08 4.15709241e-07 6.46710725e-08 4.15809241e-07 -3.54301523e-08 4.15909241e-07 5.58015891e-08 4.16009241e-07 -2.74459686e-08
+ 4.16109241e-07 4.84004265e-08 4.16209241e-07 -2.07835452e-08 4.16309241e-07 4.22245086e-08 4.16409241e-07 -1.5210292e-08 4.16509241e-07 3.70584685e-08 4.16609241e-07 -1.05742364e-08 4.16709241e-07 3.27607129e-08 4.16809241e-07 -6.70534928e-09
+ 4.16909241e-07 2.91743373e-08 4.17009241e-07 -3.47686144e-09 4.17109241e-07 2.61816051e-08 4.17209241e-07 -7.8277887e-10 4.17309241e-07 2.36842578e-08 4.17409241e-07 1.4653537e-09 4.17509241e-07 2.16193713e-08 4.17609241e-07 3.3251118e-09
+ 4.17709241e-07 1.99196335e-08 4.17809241e-07 4.85641724e-09 4.17909241e-07 1.85200862e-08 4.18009241e-07 6.11728246e-09 4.18109241e-07 1.73677097e-08 4.18209241e-07 7.1554718e-09 4.18309241e-07 1.64188499e-08 4.18409241e-07 8.0103093e-09
+ 4.18509241e-07 1.5637569e-08 4.18609241e-07 8.71417213e-09 4.18709241e-07 1.4897315e-08 4.18809241e-07 9.2799454e-09 4.18909241e-07 1.43787411e-08 4.19009241e-07 9.75062575e-09 4.19109241e-07 1.39514975e-08 4.19209241e-07 1.01384436e-08
+ 4.19309241e-07 1.35994825e-08 4.19409241e-07 1.04579695e-08 4.19509241e-07 1.33094586e-08 4.19609241e-07 1.07212252e-08 4.19709241e-07 1.30705115e-08 4.19809241e-07 1.09381179e-08 4.19909241e-07 1.28736474e-08 4.20009241e-07 1.1116812e-08
+ 4.20109241e-07 1.2711455e-08 4.20209241e-07 1.12640354e-08 4.20309241e-07 1.25778278e-08 4.20409241e-07 1.13853302e-08 4.20509241e-07 1.24677353e-08 4.20609241e-07 1.14852628e-08 4.20709241e-07 1.23770332e-08 4.20809241e-07 1.15675951e-08
+ 4.20909241e-07 1.2302306e-08 4.21009241e-07 1.1635427e-08 4.21109241e-07 1.22407403e-08 4.21209241e-07 1.16913122e-08 4.21309241e-07 1.2190018e-08 4.21409241e-07 1.17373553e-08 4.21509241e-07 1.21482294e-08 4.21609241e-07 1.17752894e-08
+ 4.21709241e-07 1.21138008e-08 4.21809241e-07 1.18065427e-08 4.21909241e-07 1.2085436e-08 4.22009241e-07 1.18322917e-08 4.22109241e-07 1.20620667e-08 4.22209241e-07 1.18535065e-08 4.22309241e-07 1.20428135e-08 4.22409241e-07 1.1870985e-08
+ 4.22509241e-07 1.20269515e-08 4.22609241e-07 1.18853856e-08 4.22709241e-07 1.20138832e-08 4.22809241e-07 1.18972499e-08 4.22909241e-07 1.20031167e-08 4.23009241e-07 1.19070249e-08 4.23109241e-07 1.19942465e-08 4.23209241e-07 1.19150785e-08
+ 4.23309241e-07 1.19869386e-08 4.23409241e-07 1.19217136e-08 4.23509241e-07 1.19809182e-08 4.23609241e-07 1.19271808e-08 4.23709241e-07 1.19759583e-08 4.23809241e-07 1.19316851e-08 4.23909241e-07 1.1971872e-08 4.24009241e-07 1.19353963e-08
+ 4.24109241e-07 1.19685052e-08 4.24209241e-07 1.19384543e-08 4.24309241e-07 1.19657318e-08 4.24409241e-07 1.19409732e-08 4.24509241e-07 1.19634471e-08 4.24609241e-07 1.19430491e-08 4.24709241e-07 1.19615647e-08 4.24809241e-07 1.19447594e-08
+ 4.24909241e-07 1.1960014e-08 4.25009241e-07 1.19461686e-08 4.25109241e-07 1.19587366e-08 4.25209241e-07 1.19473297e-08 4.25309241e-07 1.19576844e-08 4.25409241e-07 1.19482863e-08 4.25509241e-07 1.19568176e-08 4.25609241e-07 1.1949075e-08
+ 4.25709241e-07 1.19561031e-08 4.25809241e-07 1.19497245e-08 4.25909241e-07 1.1955515e-08 4.26009241e-07 1.19502597e-08 4.26109241e-07 1.19550307e-08 4.26209241e-07 1.1950701e-08 4.26309241e-07 1.19546316e-08 4.26409241e-07 1.19510642e-08
+ 4.26509241e-07 1.19543032e-08 4.26609241e-07 1.19513639e-08 4.26709241e-07 1.19540323e-08 4.26809241e-07 1.19516108e-08 4.26909241e-07 1.19538091e-08 4.27009241e-07 1.19518146e-08 4.27109241e-07 1.1953626e-08 4.27209241e-07 1.19519825e-08
+ 4.27309241e-07 1.19534745e-08 4.27409241e-07 1.19521204e-08 4.27509241e-07 1.19533501e-08 4.27609241e-07 1.19522348e-08 4.27709241e-07 1.19532475e-08 4.27809241e-07 1.19523286e-08 4.27909241e-07 1.19531632e-08 4.28009241e-07 1.19524063e-08
+ 4.28109241e-07 1.19530938e-08 4.28209241e-07 1.19524702e-08 4.28309241e-07 1.19530371e-08 4.28409241e-07 1.1952523e-08 4.28509241e-07 1.19529899e-08 4.28609241e-07 1.19525668e-08 4.28709241e-07 1.19529514e-08 4.28809241e-07 1.19526025e-08
+ 4.28909241e-07 1.19529195e-08 4.29009241e-07 1.19526321e-08 4.29109241e-07 1.19528933e-08 4.29209241e-07 1.19526568e-08 4.29309241e-07 1.19528723e-08 4.29409241e-07 1.1952677e-08 4.29509241e-07 1.19528543e-08 4.29609241e-07 1.19526941e-08
+ 4.29709241e-07 1.19528396e-08 4.29809241e-07 1.19527081e-08 4.29909241e-07 1.1952828e-08 4.30009241e-07 1.19527194e-08 4.30109241e-07 1.19528185e-08 4.30209241e-07 1.19527286e-08 4.30309241e-07 1.19528105e-08 4.30409241e-07 1.19527364e-08
+ 4.30509241e-07 1.1952804e-08 4.30609241e-07 1.19527431e-08 4.30709241e-07 1.19527989e-08 4.30809241e-07 1.19527485e-08 4.30909241e-07 1.19527944e-08 4.31009241e-07 1.19527532e-08 4.31109241e-07 1.19527912e-08 4.31209241e-07 1.1952757e-08
+ 4.31309241e-07 1.19527881e-08 4.31409241e-07 1.19527601e-08 4.31509241e-07 1.19527858e-08 4.31609241e-07 1.19527629e-08 4.31709241e-07 1.19527839e-08 4.31809241e-07 1.19527652e-08 4.31909241e-07 1.19527821e-08 4.32009241e-07 1.1952767e-08
+ 4.32109241e-07 1.19527813e-08 4.32209241e-07 1.19527684e-08 4.32309241e-07 1.19527804e-08 4.32409241e-07 1.19527696e-08 4.32509241e-07 1.195278e-08 4.32609241e-07 1.19527711e-08 4.32709241e-07 1.19527794e-08 4.32809241e-07 1.19527717e-08
+ 4.32909241e-07 1.1952779e-08 4.33009241e-07 1.1952773e-08 4.33109241e-07 1.19527787e-08 4.33209241e-07 1.19527737e-08 4.33309241e-07 1.19527785e-08 4.33409241e-07 1.19527741e-08 4.33509241e-07 1.19527783e-08 4.33609241e-07 1.1952775e-08
+ 4.33709241e-07 1.19527779e-08 4.33809241e-07 1.19527756e-08 4.33909241e-07 1.19527777e-08 4.34009241e-07 1.19527762e-08 4.34109241e-07 1.19527781e-08 4.34209241e-07 1.19527767e-08 4.34309241e-07 1.19527777e-08 4.34409241e-07 1.19527769e-08
+ 4.34509241e-07 1.19527778e-08 4.34609241e-07 1.19527773e-08 4.34709241e-07 1.19527782e-08 4.34809241e-07 1.19527776e-08 4.34909241e-07 1.19527785e-08 4.35009241e-07 1.19527776e-08 4.35109241e-07 1.19527782e-08 4.35209241e-07 1.19527781e-08
+ 4.35309241e-07 1.19527784e-08 4.35409241e-07 1.19527782e-08 4.35509241e-07 1.19527786e-08 4.35609241e-07 1.19527783e-08 4.35709241e-07 1.1952779e-08 4.35809241e-07 1.19527786e-08 4.35909241e-07 1.1952779e-08 4.36009241e-07 1.1952779e-08
+ 4.36109241e-07 1.1952779e-08 4.36209241e-07 1.19527789e-08 4.36309241e-07 1.19527792e-08 4.36409241e-07 1.19527791e-08 4.36509241e-07 1.19527795e-08 4.36609241e-07 1.19527795e-08 4.36709241e-07 1.19527793e-08 4.36809241e-07 1.19527795e-08
+ 4.36909241e-07 1.19527798e-08 4.37009241e-07 1.19527797e-08 4.37109241e-07 1.19527799e-08 4.37209241e-07 1.195278e-08 4.37309241e-07 1.19527797e-08 4.37409241e-07 1.19527801e-08 4.37509241e-07 1.19527797e-08 4.37609241e-07 1.19527805e-08
+ 4.37709241e-07 1.19527799e-08 4.37809241e-07 1.19527805e-08 4.37909241e-07 1.195278e-08 4.38009241e-07 1.1952781e-08 4.38109241e-07 1.19527803e-08 4.38209241e-07 1.19527807e-08 4.38309241e-07 1.19527805e-08 4.38409241e-07 1.19527808e-08
+ 4.38509241e-07 1.19527809e-08 4.38609241e-07 1.1952781e-08 4.38709241e-07 1.1952781e-08 4.38809241e-07 1.19527808e-08 4.38909241e-07 1.19527812e-08 4.39009241e-07 1.1952781e-08 4.39109241e-07 1.19527813e-08 4.39209241e-07 1.1952781e-08
+ 4.39309241e-07 1.19527815e-08 4.39409241e-07 1.19527813e-08 4.39509241e-07 1.19527817e-08 4.39609241e-07 1.19527811e-08 4.39709241e-07 1.19527816e-08 4.39809241e-07 1.19527815e-08 4.39909241e-07 1.1952782e-08 4.40009241e-07 1.19527815e-08
+ 4.40109241e-07 1.19527822e-08 4.40209241e-07 1.19527815e-08 4.40309241e-07 1.19527821e-08 4.40409241e-07 1.19527813e-08 4.40509241e-07 1.19527824e-08 4.40609241e-07 1.19527815e-08 4.40709241e-07 1.19527823e-08 4.40809241e-07 1.19527816e-08
+ 4.40909241e-07 1.19527827e-08 4.41009241e-07 1.1952782e-08 4.41109241e-07 1.19527822e-08 4.41209241e-07 1.19527821e-08 4.41309241e-07 1.19527824e-08 4.41409241e-07 1.1952782e-08 4.41509241e-07 1.19527825e-08 4.41609241e-07 1.19527825e-08
+ 4.41709241e-07 1.19527828e-08 4.41809241e-07 1.19527825e-08 4.41909241e-07 1.1952783e-08 4.42009241e-07 1.19527822e-08 4.42109241e-07 1.19527829e-08 4.42209241e-07 1.19527824e-08 4.42309241e-07 1.19527829e-08 4.42409241e-07 1.19527827e-08
+ 4.42509241e-07 1.19527827e-08 4.42609241e-07 1.1952783e-08 4.42709241e-07 1.19527829e-08 4.42809241e-07 1.19527831e-08 4.42909241e-07 1.19527828e-08 4.43009241e-07 1.19527832e-08 4.43109241e-07 1.1952783e-08 4.43209241e-07 1.19527833e-08
+ 4.43309241e-07 1.19527829e-08 4.43409241e-07 1.1952783e-08 4.43509241e-07 1.19527832e-08 4.43609241e-07 1.19527833e-08 4.43709241e-07 1.19527834e-08 4.43809241e-07 1.19527835e-08 4.43909241e-07 1.19527833e-08 4.44009241e-07 1.19527833e-08
+ 4.44109241e-07 1.19527836e-08 4.44209241e-07 1.19527835e-08 4.44309241e-07 1.19527835e-08 4.44409241e-07 1.19527837e-08 4.44509241e-07 1.19527833e-08 4.44609241e-07 1.19527838e-08 4.44709241e-07 1.19527838e-08 4.44809241e-07 1.19527835e-08
+ 4.44909241e-07 1.19527836e-08 4.45009241e-07 1.19527838e-08 4.45109241e-07 1.19527836e-08 4.45209241e-07 1.19527836e-08 4.45309241e-07 1.19527841e-08 4.45409241e-07 1.1952784e-08 4.45509241e-07 1.19527839e-08 4.45609241e-07 1.19527839e-08
+ 4.45709241e-07 1.19527839e-08 4.45809241e-07 1.19527838e-08 4.45909241e-07 1.19527842e-08 4.46009241e-07 1.1952784e-08 4.46109241e-07 1.19527838e-08 4.46209241e-07 1.19527843e-08 4.46309241e-07 1.19527841e-08 4.46409241e-07 1.19527842e-08
+ 4.46509241e-07 1.19527844e-08 4.46609241e-07 1.19527844e-08 4.46709241e-07 1.1952784e-08 4.46809241e-07 1.19527844e-08 4.46909241e-07 1.19527842e-08 4.47009241e-07 1.19527845e-08 4.47109241e-07 1.19527843e-08 4.47209241e-07 1.19527844e-08
+ 4.47309241e-07 1.19527845e-08 4.47409241e-07 1.19527845e-08 4.47509241e-07 1.19527846e-08 4.47609241e-07 1.19527842e-08 4.47709241e-07 1.19527848e-08 4.47809241e-07 1.19527843e-08 4.47909241e-07 1.19527848e-08 4.48009241e-07 1.19527845e-08
+ 4.48109241e-07 1.1952785e-08 4.48209241e-07 1.19527842e-08 4.48309241e-07 1.1952785e-08 4.48409241e-07 1.19527846e-08 4.48509241e-07 1.19527849e-08 4.48609241e-07 1.19527846e-08 4.48709241e-07 1.19527849e-08 4.48809241e-07 1.19527843e-08
+ 4.48909241e-07 1.19527852e-08 4.49009241e-07 1.19527847e-08 4.49109241e-07 1.19527852e-08 4.49209241e-07 1.1952785e-08 4.49309241e-07 1.19527848e-08 4.49409241e-07 1.19527849e-08 4.49509241e-07 1.19527848e-08 4.49609241e-07 1.19527849e-08
+ 4.49709241e-07 1.19527848e-08 4.49809241e-07 1.19527852e-08 4.49909241e-07 1.19527849e-08 4.50009241e-07 1.1952785e-08 4.50109241e-07 1.19527854e-08 4.50209241e-07 1.19527848e-08 4.50309241e-07 1.19527853e-08 4.50409241e-07 1.19527853e-08
+ 4.50509241e-07 1.19527851e-08 4.50609241e-07 1.1952785e-08 4.50709241e-07 1.19527854e-08 4.50809241e-07 1.1952785e-08 4.50909241e-07 1.19527855e-08 4.51e-07 1.19527851e-08 4.5101e-07 1.19386921e-08 4.5103e-07 1.20215821e-08
+ 4.5107e-07 1.18440783e-08 4.5115e-07 1.20775721e-08 4.5125e-07 1.18225586e-08 4.5135e-07 1.20783145e-08 4.5145e-07 1.18420541e-08 4.5155e-07 1.20411273e-08 4.5165e-07 1.18900525e-08 4.5175e-07 1.19863693e-08
+ 4.5185e-07 1.19530396e-08 4.51930828e-07 1.24467922e-07 4.52e-07 1.72239017e-06 4.52008608e-07 -4.6155889e-06 4.52025825e-07 -7.7865531e-06 4.52060258e-07 1.13509844e-06 4.52106181e-07 1.11144542e-05 4.52150081e-07 -1.1934542e-05
+ 4.52198026e-07 9.08990105e-06 4.5225538e-07 -8.63563247e-06 4.52312019e-07 6.70440666e-06 4.52404232e-07 -4.84172578e-06 4.52504232e-07 3.27464683e-06 4.52604232e-07 -1.93327282e-06 4.52704232e-07 9.69006195e-07 4.52804232e-07 -1.42030635e-07
+ 4.52904232e-07 -5.08190821e-07 4.53004232e-07 1.1074106e-06 4.53104232e-07 -1.58170361e-06 4.53204232e-07 2.02780267e-06 4.53304232e-07 -2.36191986e-06 4.53404232e-07 2.67940834e-06 4.53504232e-07 -2.89378902e-06 4.53604232e-07 3.10213512e-06
+ 4.53704232e-07 -3.21656805e-06 4.53804232e-07 3.33567977e-06 4.53904232e-07 -3.37016818e-06 4.54004232e-07 3.41946247e-06 4.54104232e-07 -3.39276677e-06 4.54204232e-07 3.38981241e-06 4.54304232e-07 -3.31838696e-06 4.54404232e-07 3.27818282e-06
+ 4.54504232e-07 -3.175748e-06 4.54604232e-07 3.11054471e-06 4.54704232e-07 -2.98810251e-06 4.54804232e-07 2.90756109e-06 4.54904232e-07 -2.77365299e-06 4.55004232e-07 2.68516151e-06 4.55104232e-07 -2.54622598e-06 4.55204232e-07 2.45527496e-06
+ 4.55304232e-07 -2.31602352e-06 4.55404232e-07 2.22656391e-06 4.55504232e-07 -2.0903272e-06 4.55604232e-07 2.00509543e-06 4.55704232e-07 -1.87412373e-06 4.55804232e-07 1.79491502e-06 4.55904232e-07 -1.67063204e-06 4.56004232e-07 1.59852859e-06
+ 4.56104232e-07 -1.48173646e-06 4.56204232e-07 1.4172895e-06 4.56304232e-07 -1.30833291e-06 4.56404232e-07 1.25170759e-06 4.56504232e-07 -1.15060305e-06 4.56604232e-07 1.10169152e-06 4.56704232e-07 -1.0082267e-06 4.56804232e-07 9.66733687e-07
+ 4.56904232e-07 -8.80542186e-07 4.57004232e-07 8.46049289e-07 4.57104232e-07 -7.6666751e-07 4.57204232e-07 7.3868397e-07 4.57304232e-07 -6.65596517e-07 4.57404232e-07 6.43597459e-07 4.57504232e-07 -5.76268889e-07 4.57604232e-07 5.59721194e-07
+ 4.57704232e-07 -4.97617339e-07 4.57804232e-07 4.85996962e-07 4.57904232e-07 -4.28599301e-07 4.58004232e-07 4.21403053e-07 4.58104232e-07 -3.68218431e-07 4.58204232e-07 3.64971765e-07 4.58304232e-07 -3.15538581e-07 4.58404232e-07 3.15800292e-07
+ 4.58504232e-07 -2.69691964e-07 4.58604232e-07 2.73056533e-07 4.58704232e-07 -2.2988251e-07 4.58804232e-07 2.35978874e-07 4.58904232e-07 -1.95381872e-07 4.59004232e-07 2.03872939e-07 4.59104232e-07 -1.65532531e-07 4.59204232e-07 1.76119001e-07
+ 4.59304232e-07 -1.39751474e-07 4.59404232e-07 1.52167858e-07 4.59504232e-07 -1.1752094e-07 4.59604232e-07 1.3153135e-07 4.59704232e-07 -9.83820627e-08 4.59804232e-07 1.13778877e-07 4.59904232e-07 -8.19309295e-08 4.60004232e-07 9.85312138e-08
+ 4.60104232e-07 -6.78117255e-08 4.60204232e-07 8.54545179e-08 4.60304232e-07 -5.57115593e-08 4.60404232e-07 7.42566393e-08 4.60504232e-07 -4.53590549e-08 4.60604232e-07 6.46841333e-08 4.60704232e-07 -3.65163433e-08 4.60804232e-07 5.65134236e-08
+ 4.60904232e-07 -2.89731027e-08 4.61004232e-07 4.95475204e-08 4.61104232e-07 -2.25458683e-08 4.61204232e-07 4.3615552e-08 4.61304232e-07 -1.70756622e-08 4.61404232e-07 3.85696048e-08 4.61504232e-07 -1.24250062e-08 4.61604232e-07 3.42818965e-08
+ 4.61704232e-07 -8.47524873e-09 4.61804232e-07 3.06422353e-08 4.61904232e-07 -5.12413284e-09 4.62004232e-07 2.75557193e-08 4.62104232e-07 -2.28369371e-09 4.62204232e-07 2.49408499e-08 4.62304232e-07 1.20663202e-10 4.62404232e-07 2.27293332e-08
+ 4.62504232e-07 2.14064186e-09 4.62604232e-07 2.08840208e-08 4.62704232e-07 3.82602774e-09 4.62804232e-07 1.9345039e-08 4.62904232e-07 5.23100646e-09 4.63004232e-07 1.80626872e-08 4.63104232e-07 6.40116754e-09 4.63204232e-07 1.69951488e-08
+ 4.63304232e-07 7.37485326e-09 4.63404232e-07 1.61072775e-08 4.63504232e-07 8.1842742e-09 4.63604232e-07 1.53695615e-08 4.63704232e-07 8.85646259e-09 4.63804232e-07 1.47572435e-08 4.63904232e-07 9.41408912e-09 4.64004232e-07 1.42496092e-08
+ 4.64104232e-07 9.87609011e-09 4.64204232e-07 1.38293653e-08 4.64304232e-07 1.02579408e-08 4.64404232e-07 1.34824605e-08 4.64504232e-07 1.05733335e-08 4.64604232e-07 1.31955881e-08 4.64704232e-07 1.0834203e-08 4.64804232e-07 1.2958563e-08
+ 4.64904232e-07 1.10493929e-08 4.65004232e-07 1.27633176e-08 4.65104232e-07 1.12264358e-08 4.65204232e-07 1.26028727e-08 4.65304232e-07 1.13717579e-08 4.65404232e-07 1.247132e-08 4.65504232e-07 1.14908049e-08 4.65604232e-07 1.2363581e-08
+ 4.65704232e-07 1.15882853e-08 4.65804232e-07 1.22755164e-08 4.65904232e-07 1.16677001e-08 4.66004232e-07 1.22039679e-08 4.66104232e-07 1.17321323e-08 4.66204232e-07 1.21459761e-08 4.66304232e-07 1.17842884e-08 4.66404232e-07 1.20991123e-08
+ 4.66504232e-07 1.18263538e-08 4.66604232e-07 1.20613942e-08 4.66704232e-07 1.18601356e-08 4.66804232e-07 1.20310978e-08 4.66904232e-07 1.18872595e-08 4.67004232e-07 1.20070315e-08 4.67104232e-07 1.1908574e-08 4.67204232e-07 1.19880783e-08
+ 4.67304232e-07 1.19254169e-08 4.67404232e-07 1.19731435e-08 4.67504232e-07 1.19386231e-08 4.67604232e-07 1.19615011e-08 4.67704232e-07 1.19488513e-08 4.67804232e-07 1.1952549e-08 4.67904232e-07 1.19566547e-08 4.68004232e-07 1.19457784e-08
+ 4.68104232e-07 1.19624985e-08 4.68204232e-07 1.19407655e-08 4.68304232e-07 1.19667685e-08 4.68404232e-07 1.19371595e-08 4.68504232e-07 1.19697978e-08 4.68604232e-07 1.19346251e-08 4.68704232e-07 1.19718619e-08 4.68804232e-07 1.1933019e-08
+ 4.68904232e-07 1.19730706e-08 4.69004232e-07 1.19321402e-08 4.69104232e-07 1.19736656e-08 4.69204232e-07 1.19317915e-08 4.69304232e-07 1.19738031e-08 4.69404232e-07 1.19318359e-08 4.69504232e-07 1.19735953e-08 4.69604232e-07 1.19321916e-08
+ 4.69704232e-07 1.19731111e-08 4.69804232e-07 1.19327847e-08 4.69904232e-07 1.19724275e-08 4.70004232e-07 1.19335431e-08 4.70104232e-07 1.19716068e-08 4.70204232e-07 1.1934414e-08 4.70304232e-07 1.19706962e-08 4.70404232e-07 1.19353556e-08
+ 4.70504232e-07 1.19697314e-08 4.70604232e-07 1.19363368e-08 4.70704232e-07 1.19687406e-08 4.70804232e-07 1.19373321e-08 4.70904232e-07 1.19677454e-08 4.71004232e-07 1.19383235e-08 4.71104232e-07 1.19667619e-08 4.71204232e-07 1.1939296e-08
+ 4.71304232e-07 1.19658028e-08 4.71404232e-07 1.19402393e-08 4.71504232e-07 1.19648766e-08 4.71604232e-07 1.19411469e-08 4.71704232e-07 1.19639893e-08 4.71804232e-07 1.1942013e-08 4.71904232e-07 1.19631447e-08 4.72004232e-07 1.19428352e-08
+ 4.72104232e-07 1.19623458e-08 4.72204232e-07 1.19436107e-08 4.72304232e-07 1.19615935e-08 4.72404232e-07 1.19443397e-08 4.72504232e-07 1.19608878e-08 4.72604232e-07 1.1945022e-08 4.72704232e-07 1.19602288e-08 4.72804232e-07 1.19456584e-08
+ 4.72904232e-07 1.19596146e-08 4.73004232e-07 1.19462507e-08 4.73104232e-07 1.19590438e-08 4.73204232e-07 1.19468002e-08 4.73304232e-07 1.1958515e-08 4.73404232e-07 1.19473089e-08 4.73504232e-07 1.19580261e-08 4.73604232e-07 1.19477786e-08
+ 4.73704232e-07 1.1957575e-08 4.73804232e-07 1.19482113e-08 4.73904232e-07 1.19571606e-08 4.74004232e-07 1.19486087e-08 4.74104232e-07 1.19567797e-08 4.74204232e-07 1.19489733e-08 4.74304232e-07 1.19564303e-08 4.74404232e-07 1.19493079e-08
+ 4.74504232e-07 1.19561109e-08 4.74604232e-07 1.19496138e-08 4.74704232e-07 1.1955818e-08 4.74804232e-07 1.19498936e-08 4.74904232e-07 1.19555505e-08 4.75004232e-07 1.19501491e-08 4.75104232e-07 1.1955306e-08 4.75204232e-07 1.19503829e-08
+ 4.75304232e-07 1.19550829e-08 4.75404232e-07 1.19505964e-08 4.75504232e-07 1.19548786e-08 4.75604232e-07 1.19507919e-08 4.75704232e-07 1.19546916e-08 4.75804232e-07 1.19509708e-08 4.75904232e-07 1.19545206e-08 4.76004232e-07 1.19511338e-08
+ 4.76104232e-07 1.19543651e-08 4.76204232e-07 1.19512819e-08 4.76304232e-07 1.19542241e-08 4.76404232e-07 1.19514164e-08 4.76504232e-07 1.19540959e-08 4.76604232e-07 1.19515391e-08 4.76704232e-07 1.19539788e-08 4.76804232e-07 1.19516502e-08
+ 4.76904232e-07 1.1953873e-08 4.77004232e-07 1.19517514e-08 4.77104232e-07 1.19537765e-08 4.77204232e-07 1.19518435e-08 4.77304232e-07 1.19536886e-08 4.77404232e-07 1.19519276e-08 4.77504232e-07 1.19536083e-08 4.77604232e-07 1.19520039e-08
+ 4.77704232e-07 1.19535355e-08 4.77804232e-07 1.19520734e-08 4.77904232e-07 1.19534692e-08 4.78004232e-07 1.19521368e-08 4.78104232e-07 1.19534085e-08 4.78204232e-07 1.19521944e-08 4.78304232e-07 1.19533536e-08 4.78404232e-07 1.19522471e-08
+ 4.78504232e-07 1.19533033e-08 4.78604232e-07 1.1952295e-08 4.78704232e-07 1.19532578e-08 4.78804232e-07 1.19523388e-08 4.78904232e-07 1.19532159e-08 4.79004232e-07 1.19523786e-08 4.79104232e-07 1.19531779e-08 4.79204232e-07 1.19524149e-08
+ 4.79304232e-07 1.19531433e-08 4.79404232e-07 1.19524481e-08 4.79504232e-07 1.19531115e-08 4.79604232e-07 1.19524783e-08 4.79704232e-07 1.19530826e-08 4.79804232e-07 1.19525062e-08 4.79904232e-07 1.19530563e-08 4.80004232e-07 1.19525311e-08
+ 4.80104232e-07 1.19530322e-08 4.80204232e-07 1.19525541e-08 4.80304232e-07 1.19530107e-08 4.80404232e-07 1.19525747e-08 4.80504232e-07 1.19529904e-08 4.80604232e-07 1.19525938e-08 4.80704232e-07 1.19529726e-08 4.80804232e-07 1.1952611e-08
+ 4.80904232e-07 1.19529558e-08 4.81004232e-07 1.19526269e-08 4.81104232e-07 1.19529408e-08 4.81204232e-07 1.19526414e-08 4.81304232e-07 1.19529271e-08 4.81404232e-07 1.19526548e-08 4.81504232e-07 1.19529142e-08 4.81604232e-07 1.19526669e-08
+ 4.81704232e-07 1.19529029e-08 4.81804232e-07 1.19526778e-08 4.81904232e-07 1.19528926e-08 4.82004232e-07 1.19526874e-08 4.82104232e-07 1.1952883e-08 4.82204232e-07 1.19526968e-08 4.82304232e-07 1.19528741e-08 4.82404232e-07 1.19527052e-08
+ 4.82504232e-07 1.19528661e-08 4.82604232e-07 1.19527126e-08 4.82704232e-07 1.19528589e-08 4.82804232e-07 1.19527198e-08 4.82904232e-07 1.19528524e-08 4.83004232e-07 1.19527259e-08 4.83104232e-07 1.19528467e-08 4.83204232e-07 1.19527314e-08
+ 4.83304232e-07 1.19528411e-08 4.83404232e-07 1.19527365e-08 4.83504232e-07 1.19528362e-08 4.83604232e-07 1.19527412e-08 4.83704232e-07 1.19528319e-08 4.83804232e-07 1.19527455e-08 4.83904232e-07 1.19528278e-08 4.84004232e-07 1.19527493e-08
+ 4.84104232e-07 1.19528241e-08 4.84204232e-07 1.19527531e-08 4.84304232e-07 1.19528209e-08 4.84404232e-07 1.1952756e-08 4.84504232e-07 1.19528177e-08 4.84604232e-07 1.19527588e-08 4.84704232e-07 1.1952815e-08 4.84804232e-07 1.19527614e-08
+ 4.84904232e-07 1.19528125e-08 4.85004232e-07 1.19527641e-08 4.85104232e-07 1.19528104e-08 4.85204232e-07 1.19527661e-08 4.85304232e-07 1.19528082e-08 4.85404232e-07 1.19527681e-08 4.85504232e-07 1.19528062e-08 4.85604232e-07 1.19527703e-08
+ 4.85704232e-07 1.19528042e-08 4.85804232e-07 1.19527718e-08 4.85904232e-07 1.19528027e-08 4.86004232e-07 1.19527733e-08 4.86104232e-07 1.19528012e-08 4.86204232e-07 1.19527747e-08 4.86304232e-07 1.19528002e-08 4.86404232e-07 1.19527759e-08
+ 4.86504232e-07 1.19527987e-08 4.86604232e-07 1.19527772e-08 4.86704232e-07 1.19527978e-08 4.86804232e-07 1.19527779e-08 4.86904232e-07 1.19527966e-08 4.87004232e-07 1.19527791e-08 4.87104232e-07 1.19527961e-08 4.87204232e-07 1.19527798e-08
+ 4.87304232e-07 1.19527952e-08 4.87404232e-07 1.19527809e-08 4.87504232e-07 1.19527944e-08 4.87604232e-07 1.19527814e-08 4.87704232e-07 1.19527939e-08 4.87804232e-07 1.1952782e-08 4.87904232e-07 1.19527931e-08 4.88004232e-07 1.19527825e-08
+ 4.88104232e-07 1.19527927e-08 4.88204232e-07 1.19527831e-08 4.88304232e-07 1.19527922e-08 4.88404232e-07 1.19527835e-08 4.88504232e-07 1.19527918e-08 4.88604232e-07 1.19527839e-08 4.88704232e-07 1.19527913e-08 4.88804232e-07 1.19527843e-08
+ 4.88904232e-07 1.19527912e-08 4.89004232e-07 1.19527847e-08 4.89104232e-07 1.19527906e-08 4.89204232e-07 1.19527848e-08 4.89304232e-07 1.19527906e-08 4.89404232e-07 1.19527853e-08 4.89504232e-07 1.195279e-08 4.89604232e-07 1.19527856e-08
+ 4.89704232e-07 1.19527897e-08 4.89804232e-07 1.19527858e-08 4.89904232e-07 1.19527896e-08 4.90004232e-07 1.1952786e-08 4.90104232e-07 1.19527896e-08 4.90204232e-07 1.19527863e-08 4.90304232e-07 1.19527894e-08 4.90404232e-07 1.19527863e-08
+ 4.90504232e-07 1.19527892e-08 4.90604232e-07 1.19527864e-08 4.90704232e-07 1.19527892e-08 4.90804232e-07 1.19527866e-08 4.90904232e-07 1.19527891e-08 4.91004232e-07 1.19527869e-08 4.91104232e-07 1.19527889e-08 4.91204232e-07 1.19527866e-08
+ 4.91304232e-07 1.19527888e-08 4.91404232e-07 1.19527869e-08 4.91504232e-07 1.19527884e-08 4.91604232e-07 1.19527872e-08 4.91704232e-07 1.19527885e-08 4.91804232e-07 1.19527873e-08 4.91904232e-07 1.19527886e-08 4.92004232e-07 1.19527874e-08
+ 4.92104232e-07 1.19527884e-08 4.92204232e-07 1.19527875e-08 4.92304232e-07 1.19527884e-08 4.92404232e-07 1.19527874e-08 4.92504232e-07 1.19527883e-08 4.92604232e-07 1.19527876e-08 4.92704232e-07 1.19527882e-08 4.92804232e-07 1.19527876e-08
+ 4.92904232e-07 1.1952788e-08 4.93004232e-07 1.19527878e-08 4.93104232e-07 1.1952788e-08 4.93204232e-07 1.19527877e-08 4.93304232e-07 1.19527881e-08 4.93404232e-07 1.19527878e-08 4.93504232e-07 1.19527881e-08 4.93604232e-07 1.19527875e-08
+ 4.93704232e-07 1.19527878e-08 4.93804232e-07 1.19527879e-08 4.93904232e-07 1.1952788e-08 4.94004232e-07 1.19527878e-08 4.94104232e-07 1.19527881e-08 4.94204232e-07 1.19527877e-08 4.94304232e-07 1.1952788e-08 4.94404232e-07 1.1952788e-08
+ 4.94504232e-07 1.19527876e-08 4.94604232e-07 1.19527878e-08 4.94704232e-07 1.19527879e-08 4.94804232e-07 1.19527876e-08 4.94904232e-07 1.19527879e-08 4.95004232e-07 1.1952788e-08 4.95104232e-07 1.19527879e-08 4.95204232e-07 1.19527882e-08
+ 4.95304232e-07 1.19527878e-08 4.95404232e-07 1.19527878e-08 4.95504232e-07 1.19527879e-08 4.95604232e-07 1.19527877e-08 4.95704232e-07 1.19527878e-08 4.95804232e-07 1.1952788e-08 4.95904232e-07 1.19527877e-08 4.96004232e-07 1.19527879e-08
+ 4.96104232e-07 1.1952788e-08 4.96204232e-07 1.19527876e-08 4.96304232e-07 1.19527877e-08 4.96404232e-07 1.1952788e-08 4.96504232e-07 1.1952788e-08 4.96604232e-07 1.19527878e-08 4.96704232e-07 1.19527879e-08 4.96804232e-07 1.1952788e-08
+ 4.96904232e-07 1.1952788e-08 4.97004232e-07 1.1952788e-08 4.97104232e-07 1.19527879e-08 4.97204232e-07 1.19527879e-08 4.97304232e-07 1.1952788e-08 4.97404232e-07 1.19527881e-08 4.97504232e-07 1.19527879e-08 4.97604232e-07 1.1952788e-08
+ 4.97704232e-07 1.19527878e-08 4.97804232e-07 1.19527878e-08 4.97904232e-07 1.19527876e-08 4.98004232e-07 1.19527879e-08 4.98104232e-07 1.19527878e-08 4.98204232e-07 1.19527879e-08 4.98304232e-07 1.19527878e-08 4.98404232e-07 1.1952788e-08
+ 4.98504232e-07 1.19527878e-08 4.98604232e-07 1.1952788e-08 4.98704232e-07 1.19527878e-08 4.98804232e-07 1.1952788e-08 4.98904232e-07 1.19527879e-08 4.99004232e-07 1.19527881e-08 4.99104232e-07 1.19527879e-08 4.99204232e-07 1.19527881e-08
+ 4.99304232e-07 1.19527879e-08 4.99404232e-07 1.1952788e-08 4.99504232e-07 1.1952788e-08 4.99604232e-07 1.1952788e-08 4.99704232e-07 1.1952788e-08 4.99804232e-07 1.1952788e-08 4.99904232e-07 1.1952788e-08 5e-07 1.19527881e-08
+ 5.0001e-07 1.19897009e-08 5.0003e-07 1.17744011e-08 5.0007e-07 1.22290809e-08 5.0015e-07 1.16424026e-08 5.0025e-07 1.22714108e-08 5.0035e-07 1.16453998e-08 5.0045e-07 1.22303623e-08 5.0055e-07 1.17276505e-08
+ 5.0065e-07 1.1820677e-08 5.0075e-07 2.88720796e-08 5.0085e-07 -5.4410992e-07 5.00932051e-07 7.37313015e-06 5.01e-07 -4.67316346e-05 5.01008488e-07 -5.13612331e-05 5.01025463e-07 -3.72346547e-05 5.01059414e-07 -3.10057984e-05
+ 5.0109062e-07 0.000250461008 5.0114347e-07 0.00049480124 5.01199151e-07 0.00157091292 5.01299151e-07 -0.0175241145 5.01399151e-07 0.171158646 5.01499151e-07 4.36372901 5.01599151e-07 5.20242883 5.01699151e-07 4.8824605
+ 5.01799151e-07 5.06724446 5.01893327e-07 4.9583704 5.01993327e-07 5.0269427 5.02093327e-07 4.98189925 5.02193327e-07 5.0121594 5.02293327e-07 4.99168783 5.02393327e-07 5.00564959 5.02493327e-07 4.99611607
+ 5.02593327e-07 5.00265018 5.02693327e-07 4.99817445 5.02793327e-07 5.0012475 5.02893327e-07 4.99913996 5.02993327e-07 5.00058806 5.03093327e-07 4.99959445 5.03193327e-07 5.0002773 5.03293327e-07 4.99980878
+ 5.03393327e-07 5.00013066 5.03493327e-07 4.99990996 5.03593327e-07 5.00006141 5.03693327e-07 4.99995775 5.03793327e-07 5.0000287 5.03893327e-07 4.99998031 5.03993327e-07 5.00001327 5.04093327e-07 4.99999095
+ 5.04193327e-07 5.00000601 5.04293327e-07 4.99999594 5.04393327e-07 5.00000262 5.04493327e-07 4.99999825 5.04593327e-07 5.00000105 5.04693327e-07 4.99999931 5.04793327e-07 5.00000035 5.04893327e-07 4.99999978
+ 5.04993327e-07 5.00000005 5.05093327e-07 4.99999997 5.05193327e-07 4.99999993 5.05293327e-07 5.00000003 5.05393327e-07 4.9999999 5.05493327e-07 5.00000005 5.05593327e-07 4.9999999 5.05693327e-07 5.00000004
+ 5.05793327e-07 4.99999991 5.05893327e-07 5.00000002 5.05993327e-07 4.99999993 5.06093327e-07 5.00000001 5.06193327e-07 4.99999994 5.06293327e-07 5.0 5.06393327e-07 4.99999995 5.06493327e-07 4.99999998
+ 5.06593327e-07 4.99999996 5.06693327e-07 4.99999998 5.06793327e-07 4.99999997 5.06893327e-07 4.99999997 5.06993327e-07 4.99999997 5.07093327e-07 4.99999997 5.07193327e-07 4.99999998 5.07293327e-07 4.99999996
+ 5.07393327e-07 4.99999998 5.07493327e-07 4.99999996 5.07593327e-07 4.99999998 5.07693327e-07 4.99999996 5.07793327e-07 4.99999998 5.07893327e-07 4.99999996 5.07993327e-07 4.99999998 5.08093327e-07 4.99999996
+ 5.08193327e-07 4.99999998 5.08293327e-07 4.99999996 5.08393327e-07 4.99999998 5.08493327e-07 4.99999996 5.08593327e-07 4.99999998 5.08693327e-07 4.99999996 5.08793327e-07 4.99999998 5.08893327e-07 4.99999996
+ 5.08993327e-07 4.99999998 5.09093327e-07 4.99999996 5.09193327e-07 4.99999998 5.09293327e-07 4.99999997 5.09393327e-07 4.99999998 5.09493327e-07 4.99999997 5.09593327e-07 4.99999998 5.09693327e-07 4.99999997
+ 5.09793327e-07 4.99999998 5.09893327e-07 4.99999997 5.09993327e-07 4.99999998 5.10093327e-07 4.99999997 5.10193327e-07 4.99999998 5.10293327e-07 4.99999997 5.10393327e-07 4.99999998 5.10493327e-07 4.99999997
+ 5.10593327e-07 4.99999998 5.10693327e-07 4.99999997 5.10793327e-07 4.99999998 5.10893327e-07 4.99999997 5.10993327e-07 4.99999997 5.11093327e-07 4.99999997 5.11193327e-07 4.99999997 5.11293327e-07 4.99999997
+ 5.11393327e-07 4.99999997 5.11493327e-07 4.99999997 5.11593327e-07 4.99999997 5.11693327e-07 4.99999997 5.11793327e-07 4.99999997 5.11893327e-07 4.99999997 5.11993327e-07 4.99999997 5.12093327e-07 4.99999997
+ 5.12193327e-07 4.99999997 5.12293327e-07 4.99999997 5.12393327e-07 4.99999997 5.12493327e-07 4.99999997 5.12593327e-07 4.99999997 5.12693327e-07 4.99999997 5.12793327e-07 4.99999997 5.12893327e-07 4.99999997
+ 5.12993327e-07 4.99999997 5.13093327e-07 4.99999997 5.13193327e-07 4.99999997 5.13293327e-07 4.99999997 5.13393327e-07 4.99999997 5.13493327e-07 4.99999997 5.13593327e-07 4.99999997 5.13693327e-07 4.99999997
+ 5.13793327e-07 4.99999997 5.13893327e-07 4.99999997 5.13993327e-07 4.99999997 5.14093327e-07 4.99999997 5.14193327e-07 4.99999997 5.14293327e-07 4.99999997 5.14393327e-07 4.99999997 5.14493327e-07 4.99999997
+ 5.14593327e-07 4.99999997 5.14693327e-07 4.99999997 5.14793327e-07 4.99999997 5.14893327e-07 4.99999997 5.14993327e-07 4.99999997 5.15093327e-07 4.99999997 5.15193327e-07 4.99999997 5.15293327e-07 4.99999997
+ 5.15393327e-07 4.99999997 5.15493327e-07 4.99999997 5.15593327e-07 4.99999997 5.15693327e-07 4.99999997 5.15793327e-07 4.99999997 5.15893327e-07 4.99999997 5.15993327e-07 4.99999997 5.16093327e-07 4.99999997
+ 5.16193327e-07 4.99999997 5.16293327e-07 4.99999997 5.16393327e-07 4.99999997 5.16493327e-07 4.99999997 5.16593327e-07 4.99999997 5.16693327e-07 4.99999997 5.16793327e-07 4.99999997 5.16893327e-07 4.99999997
+ 5.16993327e-07 4.99999997 5.17093327e-07 4.99999997 5.17193327e-07 4.99999997 5.17293327e-07 4.99999997 5.17393327e-07 4.99999997 5.17493327e-07 4.99999997 5.17593327e-07 4.99999997 5.17693327e-07 4.99999997
+ 5.17793327e-07 4.99999997 5.17893327e-07 4.99999997 5.17993327e-07 4.99999997 5.18093327e-07 4.99999997 5.18193327e-07 4.99999997 5.18293327e-07 4.99999997 5.18393327e-07 4.99999997 5.18493327e-07 4.99999997
+ 5.18593327e-07 4.99999997 5.18693327e-07 4.99999997 5.18793327e-07 4.99999997 5.18893327e-07 4.99999997 5.18993327e-07 4.99999997 5.19093327e-07 4.99999997 5.19193327e-07 4.99999997 5.19293327e-07 4.99999997
+ 5.19393327e-07 4.99999997 5.19493327e-07 4.99999997 5.19593327e-07 4.99999997 5.19693327e-07 4.99999997 5.19793327e-07 4.99999997 5.19893327e-07 4.99999997 5.19993327e-07 4.99999997 5.20093327e-07 4.99999997
+ 5.20193327e-07 4.99999997 5.20293327e-07 4.99999997 5.20393327e-07 4.99999997 5.20493327e-07 4.99999997 5.20593327e-07 4.99999997 5.20693327e-07 4.99999997 5.20793327e-07 4.99999997 5.20893327e-07 4.99999997
+ 5.20993327e-07 4.99999997 5.21093327e-07 4.99999997 5.21193327e-07 4.99999997 5.21293327e-07 4.99999997 5.21393327e-07 4.99999997 5.21493327e-07 4.99999997 5.21593327e-07 4.99999997 5.21693327e-07 4.99999997
+ 5.21793327e-07 4.99999997 5.21893327e-07 4.99999997 5.21993327e-07 4.99999997 5.22093327e-07 4.99999997 5.22193327e-07 4.99999997 5.22293327e-07 4.99999997 5.22393327e-07 4.99999997 5.22493327e-07 4.99999997
+ 5.22593327e-07 4.99999997 5.22693327e-07 4.99999997 5.22793327e-07 4.99999997 5.22893327e-07 4.99999997 5.22993327e-07 4.99999997 5.23093327e-07 4.99999997 5.23193327e-07 4.99999997 5.23293327e-07 4.99999997
+ 5.23393327e-07 4.99999997 5.23493327e-07 4.99999997 5.23593327e-07 4.99999997 5.23693327e-07 4.99999997 5.23793327e-07 4.99999997 5.23893327e-07 4.99999997 5.23993327e-07 4.99999997 5.24093327e-07 4.99999997
+ 5.24193327e-07 4.99999997 5.24293327e-07 4.99999997 5.24393327e-07 4.99999997 5.24493327e-07 4.99999997 5.24593327e-07 4.99999997 5.24693327e-07 4.99999997 5.24793327e-07 4.99999997 5.24893327e-07 4.99999997
+ 5.24993327e-07 4.99999997 5.25093327e-07 4.99999997 5.25193327e-07 4.99999997 5.25293327e-07 4.99999997 5.25393327e-07 4.99999997 5.25493327e-07 4.99999997 5.25593327e-07 4.99999997 5.25693327e-07 4.99999997
+ 5.25793327e-07 4.99999997 5.25893327e-07 4.99999997 5.25993327e-07 4.99999997 5.26093327e-07 4.99999997 5.26193327e-07 4.99999997 5.26293327e-07 4.99999997 5.26393327e-07 4.99999997 5.26493327e-07 4.99999997
+ 5.26593327e-07 4.99999997 5.26693327e-07 4.99999997 5.26793327e-07 4.99999997 5.26893327e-07 4.99999997 5.26993327e-07 4.99999997 5.27093327e-07 4.99999997 5.27193327e-07 4.99999997 5.27293327e-07 4.99999997
+ 5.27393327e-07 4.99999997 5.27493327e-07 4.99999997 5.27593327e-07 4.99999997 5.27693327e-07 4.99999997 5.27793327e-07 4.99999997 5.27893327e-07 4.99999997 5.27993327e-07 4.99999997 5.28093327e-07 4.99999997
+ 5.28193327e-07 4.99999997 5.28293327e-07 4.99999997 5.28393327e-07 4.99999997 5.28493327e-07 4.99999997 5.28593327e-07 4.99999997 5.28693327e-07 4.99999997 5.28793327e-07 4.99999997 5.28893327e-07 4.99999997
+ 5.28993327e-07 4.99999997 5.29093327e-07 4.99999997 5.29193327e-07 4.99999997 5.29293327e-07 4.99999997 5.29393327e-07 4.99999997 5.29493327e-07 4.99999997 5.29593327e-07 4.99999997 5.29693327e-07 4.99999997
+ 5.29793327e-07 4.99999997 5.29893327e-07 4.99999997 5.29993327e-07 4.99999997 5.30093327e-07 4.99999997 5.30193327e-07 4.99999997 5.30293327e-07 4.99999997 5.30393327e-07 4.99999997 5.30493327e-07 4.99999997
+ 5.30593327e-07 4.99999997 5.30693327e-07 4.99999997 5.30793327e-07 4.99999997 5.30893327e-07 4.99999997 5.30993327e-07 4.99999997 5.31093327e-07 4.99999997 5.31193327e-07 4.99999997 5.31293327e-07 4.99999997
+ 5.31393327e-07 4.99999997 5.31493327e-07 4.99999997 5.31593327e-07 4.99999997 5.31693327e-07 4.99999997 5.31793327e-07 4.99999997 5.31893327e-07 4.99999997 5.31993327e-07 4.99999997 5.32093327e-07 4.99999997
+ 5.32193327e-07 4.99999997 5.32293327e-07 4.99999997 5.32393327e-07 4.99999997 5.32493327e-07 4.99999997 5.32593327e-07 4.99999997 5.32693327e-07 4.99999997 5.32793327e-07 4.99999997 5.32893327e-07 4.99999997
+ 5.32993327e-07 4.99999997 5.33093327e-07 4.99999997 5.33193327e-07 4.99999997 5.33293327e-07 4.99999997 5.33393327e-07 4.99999997 5.33493327e-07 4.99999997 5.33593327e-07 4.99999997 5.33693327e-07 4.99999997
+ 5.33793327e-07 4.99999997 5.33893327e-07 4.99999997 5.33993327e-07 4.99999997 5.34093327e-07 4.99999997 5.34193327e-07 4.99999997 5.34293327e-07 4.99999997 5.34393327e-07 4.99999997 5.34493327e-07 4.99999997
+ 5.34593327e-07 4.99999997 5.34693327e-07 4.99999997 5.34793327e-07 4.99999997 5.34893327e-07 4.99999997 5.34993327e-07 4.99999997 5.35093327e-07 4.99999997 5.35193327e-07 4.99999997 5.35293327e-07 4.99999997
+ 5.35393327e-07 4.99999997 5.35493327e-07 4.99999997 5.35593327e-07 4.99999997 5.35693327e-07 4.99999997 5.35793327e-07 4.99999997 5.35893327e-07 4.99999997 5.35993327e-07 4.99999997 5.36093327e-07 4.99999997
+ 5.36193327e-07 4.99999997 5.36293327e-07 4.99999997 5.36393327e-07 4.99999997 5.36493327e-07 4.99999997 5.36593327e-07 4.99999997 5.36693327e-07 4.99999997 5.36793327e-07 4.99999997 5.36893327e-07 4.99999997
+ 5.36993327e-07 4.99999997 5.37093327e-07 4.99999997 5.37193327e-07 4.99999997 5.37293327e-07 4.99999997 5.37393327e-07 4.99999997 5.37493327e-07 4.99999997 5.37593327e-07 4.99999997 5.37693327e-07 4.99999997
+ 5.37793327e-07 4.99999997 5.37893327e-07 4.99999997 5.37993327e-07 4.99999997 5.38093327e-07 4.99999997 5.38193327e-07 4.99999997 5.38293327e-07 4.99999997 5.38393327e-07 4.99999997 5.38493327e-07 4.99999997
+ 5.38593327e-07 4.99999997 5.38693327e-07 4.99999997 5.38793327e-07 4.99999997 5.38893327e-07 4.99999997 5.38993327e-07 4.99999997 5.39093327e-07 4.99999997 5.39193327e-07 4.99999997 5.39293327e-07 4.99999997
+ 5.39393327e-07 4.99999997 5.39493327e-07 4.99999997 5.39593327e-07 4.99999997 5.39693327e-07 4.99999997 5.39793327e-07 4.99999997 5.39893327e-07 4.99999997 5.39993327e-07 4.99999997 5.40093327e-07 4.99999997
+ 5.40193327e-07 4.99999997 5.40293327e-07 4.99999997 5.40393327e-07 4.99999997 5.40493327e-07 4.99999997 5.40593327e-07 4.99999997 5.40693327e-07 4.99999997 5.40793327e-07 4.99999997 5.40893327e-07 4.99999997
+ 5.40993327e-07 4.99999997 5.41093327e-07 4.99999997 5.41193327e-07 4.99999997 5.41293327e-07 4.99999997 5.41393327e-07 4.99999997 5.41493327e-07 4.99999997 5.41593327e-07 4.99999997 5.41693327e-07 4.99999997
+ 5.41793327e-07 4.99999997 5.41893327e-07 4.99999997 5.41993327e-07 4.99999997 5.42093327e-07 4.99999997 5.42193327e-07 4.99999997 5.42293327e-07 4.99999997 5.42393327e-07 4.99999997 5.42493327e-07 4.99999997
+ 5.42593327e-07 4.99999997 5.42693327e-07 4.99999997 5.42793327e-07 4.99999997 5.42893327e-07 4.99999997 5.42993327e-07 4.99999997 5.43093327e-07 4.99999997 5.43193327e-07 4.99999997 5.43293327e-07 4.99999997
+ 5.43393327e-07 4.99999997 5.43493327e-07 4.99999997 5.43593327e-07 4.99999997 5.43693327e-07 4.99999997 5.43793327e-07 4.99999997 5.43893327e-07 4.99999997 5.43993327e-07 4.99999997 5.44093327e-07 4.99999997
+ 5.44193327e-07 4.99999997 5.44293327e-07 4.99999997 5.44393327e-07 4.99999997 5.44493327e-07 4.99999997 5.44593327e-07 4.99999997 5.44693327e-07 4.99999997 5.44793327e-07 4.99999997 5.44893327e-07 4.99999997
+ 5.44993327e-07 4.99999997 5.45093327e-07 4.99999997 5.45193327e-07 4.99999997 5.45293327e-07 4.99999997 5.45393327e-07 4.99999997 5.45493327e-07 4.99999997 5.45593327e-07 4.99999997 5.45693327e-07 4.99999997
+ 5.45793327e-07 4.99999997 5.45893327e-07 4.99999997 5.45993327e-07 4.99999997 5.46093327e-07 4.99999997 5.46193327e-07 4.99999997 5.46293327e-07 4.99999997 5.46393327e-07 4.99999997 5.46493327e-07 4.99999997
+ 5.46593327e-07 4.99999997 5.46693327e-07 4.99999997 5.46793327e-07 4.99999997 5.46893327e-07 4.99999997 5.46993327e-07 4.99999997 5.47093327e-07 4.99999997 5.47193327e-07 4.99999997 5.47293327e-07 4.99999997
+ 5.47393327e-07 4.99999997 5.47493327e-07 4.99999997 5.47593327e-07 4.99999997 5.47693327e-07 4.99999997 5.47793327e-07 4.99999997 5.47893327e-07 4.99999997 5.47993327e-07 4.99999997 5.48093327e-07 4.99999997
+ 5.48193327e-07 4.99999997 5.48293327e-07 4.99999997 5.48393327e-07 4.99999997 5.48493327e-07 4.99999997 5.48593327e-07 4.99999997 5.48693327e-07 4.99999997 5.48793327e-07 4.99999997 5.48893327e-07 4.99999997
+ 5.48993327e-07 4.99999997 5.49093327e-07 4.99999997 5.49193327e-07 4.99999997 5.49293327e-07 4.99999997 5.49393327e-07 4.99999997 5.49493327e-07 4.99999997 5.49593327e-07 4.99999997 5.49693327e-07 4.99999997
+ 5.49793327e-07 4.99999997 5.49893327e-07 4.99999997 5.49993327e-07 4.99999997 5.50093327e-07 4.99999997 5.50193327e-07 4.99999997 5.50293327e-07 4.99999997 5.50393327e-07 4.99999997 5.50493327e-07 4.99999997
+ 5.50593327e-07 4.99999997 5.50693327e-07 4.99999997 5.50793327e-07 4.99999997 5.50893327e-07 4.99999997 5.50993327e-07 4.99999997 5.51e-07 4.99999997 5.5101e-07 4.99999997 5.5103e-07 4.99999997
+ 5.5107e-07 4.99999997 5.5115e-07 4.99999997 5.5125e-07 4.99999997 5.5135e-07 4.99999997 5.5145e-07 4.99999997 5.5155e-07 4.99999997 5.5165e-07 4.99999997 5.5175e-07 4.99999997
+ 5.5185e-07 4.99999997 5.51930828e-07 5.00000065 5.52e-07 5.00000149 5.52008608e-07 4.99999288 5.52025825e-07 4.99997549 5.52060258e-07 4.99999257 5.52106188e-07 5.00004375 5.52150118e-07 5.00000856
+ 5.5219811e-07 4.99994581 5.52255501e-07 5.00002983 5.52312176e-07 4.99999321 5.52404431e-07 5.00000355 5.52490774e-07 5.00000011 5.52590774e-07 4.99999756 5.52690774e-07 5.00000329 5.52790774e-07 4.99999639
+ 5.52890774e-07 5.0000034 5.52990774e-07 4.99999687 5.53090774e-07 5.00000266 5.53190774e-07 4.9999977 5.53290774e-07 5.00000186 5.53390774e-07 4.99999842 5.53490774e-07 5.00000123 5.53590774e-07 4.99999895
+ 5.53690774e-07 5.00000079 5.53790774e-07 4.99999931 5.53890774e-07 5.00000051 5.53990774e-07 4.99999954 5.54090774e-07 5.00000033 5.54190774e-07 4.99999968 5.54290774e-07 5.00000021 5.54390774e-07 4.99999977
+ 5.54490774e-07 5.00000014 5.54590774e-07 4.99999983 5.54690774e-07 5.00000009 5.54790774e-07 4.99999987 5.54890774e-07 5.00000007 5.54990774e-07 4.99999989 5.55090774e-07 5.00000005 5.55190774e-07 4.99999991
+ 5.55290774e-07 5.00000003 5.55390774e-07 4.99999992 5.55490774e-07 5.00000002 5.55590774e-07 4.99999993 5.55690774e-07 5.00000001 5.55790774e-07 4.99999993 5.55890774e-07 5.00000001 5.55990774e-07 4.99999994
+ 5.56090774e-07 5.0 5.56190774e-07 4.99999994 5.56290774e-07 5.0 5.56390774e-07 4.99999995 5.56490774e-07 5.0 5.56590774e-07 4.99999995 5.56690774e-07 4.99999999 5.56790774e-07 4.99999995
+ 5.56890774e-07 4.99999999 5.56990774e-07 4.99999996 5.57090774e-07 4.99999999 5.57190774e-07 4.99999996 5.57290774e-07 4.99999999 5.57390774e-07 4.99999996 5.57490774e-07 4.99999998 5.57590774e-07 4.99999996
+ 5.57690774e-07 4.99999998 5.57790774e-07 4.99999996 5.57890774e-07 4.99999998 5.57990774e-07 4.99999996 5.58090774e-07 4.99999998 5.58190774e-07 4.99999997 5.58290774e-07 4.99999998 5.58390774e-07 4.99999997
+ 5.58490774e-07 4.99999998 5.58590774e-07 4.99999997 5.58690774e-07 4.99999998 5.58790774e-07 4.99999997 5.58890774e-07 4.99999998 5.58990774e-07 4.99999997 5.59090774e-07 4.99999998 5.59190774e-07 4.99999997
+ 5.59290774e-07 4.99999997 5.59390774e-07 4.99999997 5.59490774e-07 4.99999997 5.59590774e-07 4.99999997 5.59690774e-07 4.99999997 5.59790774e-07 4.99999997 5.59890774e-07 4.99999997 5.59990774e-07 4.99999997
+ 5.60090774e-07 4.99999997 5.60190774e-07 4.99999997 5.60290774e-07 4.99999997 5.60390774e-07 4.99999997 5.60490774e-07 4.99999997 5.60590774e-07 4.99999997 5.60690774e-07 4.99999997 5.60790774e-07 4.99999997
+ 5.60890774e-07 4.99999997 5.60990774e-07 4.99999997 5.61090774e-07 4.99999997 5.61190774e-07 4.99999997 5.61290774e-07 4.99999997 5.61390774e-07 4.99999997 5.61490774e-07 4.99999997 5.61590774e-07 4.99999997
+ 5.61690774e-07 4.99999997 5.61790774e-07 4.99999997 5.61890774e-07 4.99999997 5.61990774e-07 4.99999997 5.62090774e-07 4.99999997 5.62190774e-07 4.99999997 5.62290774e-07 4.99999997 5.62390774e-07 4.99999997
+ 5.62490774e-07 4.99999997 5.62590774e-07 4.99999997 5.62690774e-07 4.99999997 5.62790774e-07 4.99999997 5.62890774e-07 4.99999997 5.62990774e-07 4.99999997 5.63090774e-07 4.99999997 5.63190774e-07 4.99999997
+ 5.63290774e-07 4.99999997 5.63390774e-07 4.99999997 5.63490774e-07 4.99999997 5.63590774e-07 4.99999997 5.63690774e-07 4.99999997 5.63790774e-07 4.99999997 5.63890774e-07 4.99999997 5.63990774e-07 4.99999997
+ 5.64090774e-07 4.99999997 5.64190774e-07 4.99999997 5.64290774e-07 4.99999997 5.64390774e-07 4.99999997 5.64490774e-07 4.99999997 5.64590774e-07 4.99999997 5.64690774e-07 4.99999997 5.64790774e-07 4.99999997
+ 5.64890774e-07 4.99999997 5.64990774e-07 4.99999997 5.65090774e-07 4.99999997 5.65190774e-07 4.99999997 5.65290774e-07 4.99999997 5.65390774e-07 4.99999997 5.65490774e-07 4.99999997 5.65590774e-07 4.99999997
+ 5.65690774e-07 4.99999997 5.65790774e-07 4.99999997 5.65890774e-07 4.99999997 5.65990774e-07 4.99999997 5.66090774e-07 4.99999997 5.66190774e-07 4.99999997 5.66290774e-07 4.99999997 5.66390774e-07 4.99999997
+ 5.66490774e-07 4.99999997 5.66590774e-07 4.99999997 5.66690774e-07 4.99999997 5.66790774e-07 4.99999997 5.66890774e-07 4.99999997 5.66990774e-07 4.99999997 5.67090774e-07 4.99999997 5.67190774e-07 4.99999997
+ 5.67290774e-07 4.99999997 5.67390774e-07 4.99999997 5.67490774e-07 4.99999997 5.67590774e-07 4.99999997 5.67690774e-07 4.99999997 5.67790774e-07 4.99999997 5.67890774e-07 4.99999997 5.67990774e-07 4.99999997
+ 5.68090774e-07 4.99999997 5.68190774e-07 4.99999997 5.68290774e-07 4.99999997 5.68390774e-07 4.99999997 5.68490774e-07 4.99999997 5.68590774e-07 4.99999997 5.68690774e-07 4.99999997 5.68790774e-07 4.99999997
+ 5.68890774e-07 4.99999997 5.68990774e-07 4.99999997 5.69090774e-07 4.99999997 5.69190774e-07 4.99999997 5.69290774e-07 4.99999997 5.69390774e-07 4.99999997 5.69490774e-07 4.99999997 5.69590774e-07 4.99999997
+ 5.69690774e-07 4.99999997 5.69790774e-07 4.99999997 5.69890774e-07 4.99999997 5.69990774e-07 4.99999997 5.70090774e-07 4.99999997 5.70190774e-07 4.99999997 5.70290774e-07 4.99999997 5.70390774e-07 4.99999997
+ 5.70490774e-07 4.99999997 5.70590774e-07 4.99999997 5.70690774e-07 4.99999997 5.70790774e-07 4.99999997 5.70890774e-07 4.99999997 5.70990774e-07 4.99999997 5.71090774e-07 4.99999997 5.71190774e-07 4.99999997
+ 5.71290774e-07 4.99999997 5.71390774e-07 4.99999997 5.71490774e-07 4.99999997 5.71590774e-07 4.99999997 5.71690774e-07 4.99999997 5.71790774e-07 4.99999997 5.71890774e-07 4.99999997 5.71990774e-07 4.99999997
+ 5.72090774e-07 4.99999997 5.72190774e-07 4.99999997 5.72290774e-07 4.99999997 5.72390774e-07 4.99999997 5.72490774e-07 4.99999997 5.72590774e-07 4.99999997 5.72690774e-07 4.99999997 5.72790774e-07 4.99999997
+ 5.72890774e-07 4.99999997 5.72990774e-07 4.99999997 5.73090774e-07 4.99999997 5.73190774e-07 4.99999997 5.73290774e-07 4.99999997 5.73390774e-07 4.99999997 5.73490774e-07 4.99999997 5.73590774e-07 4.99999997
+ 5.73690774e-07 4.99999997 5.73790774e-07 4.99999997 5.73890774e-07 4.99999997 5.73990774e-07 4.99999997 5.74090774e-07 4.99999997 5.74190774e-07 4.99999997 5.74290774e-07 4.99999997 5.74390774e-07 4.99999997
+ 5.74490774e-07 4.99999997 5.74590774e-07 4.99999997 5.74690774e-07 4.99999997 5.74790774e-07 4.99999997 5.74890774e-07 4.99999997 5.74990774e-07 4.99999997 5.75090774e-07 4.99999997 5.75190774e-07 4.99999997
+ 5.75290774e-07 4.99999997 5.75390774e-07 4.99999997 5.75490774e-07 4.99999997 5.75590774e-07 4.99999997 5.75690774e-07 4.99999997 5.75790774e-07 4.99999997 5.75890774e-07 4.99999997 5.75990774e-07 4.99999997
+ 5.76090774e-07 4.99999997 5.76190774e-07 4.99999997 5.76290774e-07 4.99999997 5.76390774e-07 4.99999997 5.76490774e-07 4.99999997 5.76590774e-07 4.99999997 5.76690774e-07 4.99999997 5.76790774e-07 4.99999997
+ 5.76890774e-07 4.99999997 5.76990774e-07 4.99999997 5.77090774e-07 4.99999997 5.77190774e-07 4.99999997 5.77290774e-07 4.99999997 5.77390774e-07 4.99999997 5.77490774e-07 4.99999997 5.77590774e-07 4.99999997
+ 5.77690774e-07 4.99999997 5.77790774e-07 4.99999997 5.77890774e-07 4.99999997 5.77990774e-07 4.99999997 5.78090774e-07 4.99999997 5.78190774e-07 4.99999997 5.78290774e-07 4.99999997 5.78390774e-07 4.99999997
+ 5.78490774e-07 4.99999997 5.78590774e-07 4.99999997 5.78690774e-07 4.99999997 5.78790774e-07 4.99999997 5.78890774e-07 4.99999997 5.78990774e-07 4.99999997 5.79090774e-07 4.99999997 5.79190774e-07 4.99999997
+ 5.79290774e-07 4.99999997 5.79390774e-07 4.99999997 5.79490774e-07 4.99999997 5.79590774e-07 4.99999997 5.79690774e-07 4.99999997 5.79790774e-07 4.99999997 5.79890774e-07 4.99999997 5.79990774e-07 4.99999997
+ 5.80090774e-07 4.99999997 5.80190774e-07 4.99999997 5.80290774e-07 4.99999997 5.80390774e-07 4.99999997 5.80490774e-07 4.99999997 5.80590774e-07 4.99999997 5.80690774e-07 4.99999997 5.80790774e-07 4.99999997
+ 5.80890774e-07 4.99999997 5.80990774e-07 4.99999997 5.81090774e-07 4.99999997 5.81190774e-07 4.99999997 5.81290774e-07 4.99999997 5.81390774e-07 4.99999997 5.81490774e-07 4.99999997 5.81590774e-07 4.99999997
+ 5.81690774e-07 4.99999997 5.81790774e-07 4.99999997 5.81890774e-07 4.99999997 5.81990774e-07 4.99999997 5.82090774e-07 4.99999997 5.82190774e-07 4.99999997 5.82290774e-07 4.99999997 5.82390774e-07 4.99999997
+ 5.82490774e-07 4.99999997 5.82590774e-07 4.99999997 5.82690774e-07 4.99999997 5.82790774e-07 4.99999997 5.82890774e-07 4.99999997 5.82990774e-07 4.99999997 5.83090774e-07 4.99999997 5.83190774e-07 4.99999997
+ 5.83290774e-07 4.99999997 5.83390774e-07 4.99999997 5.83490774e-07 4.99999997 5.83590774e-07 4.99999997 5.83690774e-07 4.99999997 5.83790774e-07 4.99999997 5.83890774e-07 4.99999997 5.83990774e-07 4.99999997
+ 5.84090774e-07 4.99999997 5.84190774e-07 4.99999997 5.84290774e-07 4.99999997 5.84390774e-07 4.99999997 5.84490774e-07 4.99999997 5.84590774e-07 4.99999997 5.84690774e-07 4.99999997 5.84790774e-07 4.99999997
+ 5.84890774e-07 4.99999997 5.84990774e-07 4.99999997 5.85090774e-07 4.99999997 5.85190774e-07 4.99999997 5.85290774e-07 4.99999997 5.85390774e-07 4.99999997 5.85490774e-07 4.99999997 5.85590774e-07 4.99999997
+ 5.85690774e-07 4.99999997 5.85790774e-07 4.99999997 5.85890774e-07 4.99999997 5.85990774e-07 4.99999997 5.86090774e-07 4.99999997 5.86190774e-07 4.99999997 5.86290774e-07 4.99999997 5.86390774e-07 4.99999997
+ 5.86490774e-07 4.99999997 5.86590774e-07 4.99999997 5.86690774e-07 4.99999997 5.86790774e-07 4.99999997 5.86890774e-07 4.99999997 5.86990774e-07 4.99999997 5.87090774e-07 4.99999997 5.87190774e-07 4.99999997
+ 5.87290774e-07 4.99999997 5.87390774e-07 4.99999997 5.87490774e-07 4.99999997 5.87590774e-07 4.99999997 5.87690774e-07 4.99999997 5.87790774e-07 4.99999997 5.87890774e-07 4.99999997 5.87990774e-07 4.99999997
+ 5.88090774e-07 4.99999997 5.88190774e-07 4.99999997 5.88290774e-07 4.99999997 5.88390774e-07 4.99999997 5.88490774e-07 4.99999997 5.88590774e-07 4.99999997 5.88690774e-07 4.99999997 5.88790774e-07 4.99999997
+ 5.88890774e-07 4.99999997 5.88990774e-07 4.99999997 5.89090774e-07 4.99999997 5.89190774e-07 4.99999997 5.89290774e-07 4.99999997 5.89390774e-07 4.99999997 5.89490774e-07 4.99999997 5.89590774e-07 4.99999997
+ 5.89690774e-07 4.99999997 5.89790774e-07 4.99999997 5.89890774e-07 4.99999997 5.89990774e-07 4.99999997 5.90090774e-07 4.99999997 5.90190774e-07 4.99999997 5.90290774e-07 4.99999997 5.90390774e-07 4.99999997
+ 5.90490774e-07 4.99999997 5.90590774e-07 4.99999997 5.90690774e-07 4.99999997 5.90790774e-07 4.99999997 5.90890774e-07 4.99999997 5.90990774e-07 4.99999997 5.91090774e-07 4.99999997 5.91190774e-07 4.99999997
+ 5.91290774e-07 4.99999997 5.91390774e-07 4.99999997 5.91490774e-07 4.99999997 5.91590774e-07 4.99999997 5.91690774e-07 4.99999997 5.91790774e-07 4.99999997 5.91890774e-07 4.99999997 5.91990774e-07 4.99999997
+ 5.92090774e-07 4.99999997 5.92190774e-07 4.99999997 5.92290774e-07 4.99999997 5.92390774e-07 4.99999997 5.92490774e-07 4.99999997 5.92590774e-07 4.99999997 5.92690774e-07 4.99999997 5.92790774e-07 4.99999997
+ 5.92890774e-07 4.99999997 5.92990774e-07 4.99999997 5.93090774e-07 4.99999997 5.93190774e-07 4.99999997 5.93290774e-07 4.99999997 5.93390774e-07 4.99999997 5.93490774e-07 4.99999997 5.93590774e-07 4.99999997
+ 5.93690774e-07 4.99999997 5.93790774e-07 4.99999997 5.93890774e-07 4.99999997 5.93990774e-07 4.99999997 5.94090774e-07 4.99999997 5.94190774e-07 4.99999997 5.94290774e-07 4.99999997 5.94390774e-07 4.99999997
+ 5.94490774e-07 4.99999997 5.94590774e-07 4.99999997 5.94690774e-07 4.99999997 5.94790774e-07 4.99999997 5.94890774e-07 4.99999997 5.94990774e-07 4.99999997 5.95090774e-07 4.99999997 5.95190774e-07 4.99999997
+ 5.95290774e-07 4.99999997 5.95390774e-07 4.99999997 5.95490774e-07 4.99999997 5.95590774e-07 4.99999997 5.95690774e-07 4.99999997 5.95790774e-07 4.99999997 5.95890774e-07 4.99999997 5.95990774e-07 4.99999997
+ 5.96090774e-07 4.99999997 5.96190774e-07 4.99999997 5.96290774e-07 4.99999997 5.96390774e-07 4.99999997 5.96490774e-07 4.99999997 5.96590774e-07 4.99999997 5.96690774e-07 4.99999997 5.96790774e-07 4.99999997
+ 5.96890774e-07 4.99999997 5.96990774e-07 4.99999997 5.97090774e-07 4.99999997 5.97190774e-07 4.99999997 5.97290774e-07 4.99999997 5.97390774e-07 4.99999997 5.97490774e-07 4.99999997 5.97590774e-07 4.99999997
+ 5.97690774e-07 4.99999997 5.97790774e-07 4.99999997 5.97890774e-07 4.99999997 5.97990774e-07 4.99999997 5.98090774e-07 4.99999997 5.98190774e-07 4.99999997 5.98290774e-07 4.99999997 5.98390774e-07 4.99999997
+ 5.98490774e-07 4.99999997 5.98590774e-07 4.99999997 5.98690774e-07 4.99999997 5.98790774e-07 4.99999997 5.98890774e-07 4.99999997 5.98990774e-07 4.99999997 5.99090774e-07 4.99999997 5.99190774e-07 4.99999997
+ 5.99290774e-07 4.99999997 5.99390774e-07 4.99999997 5.99490774e-07 4.99999997 5.99590774e-07 4.99999997 5.99690774e-07 4.99999997 5.99790774e-07 4.99999997 5.99890774e-07 4.99999997 5.99990774e-07 4.99999997
+ 6e-07 4.99999997 6.0001e-07 4.99999997 6.0003e-07 4.99999997 6.0007e-07 4.99999997 6.0015e-07 4.99999997 6.0025e-07 4.99999997 6.0035e-07 4.99999997 6.0045e-07 4.99999997
+ 6.0055e-07 4.99999997 6.0065e-07 4.99999997 6.0075e-07 5.00000001 6.0085e-07 4.99999718 6.00932239e-07 5.00000338 6.01e-07 5.00008492 6.01008502e-07 5.000115 6.01025505e-07 5.00022464
+ 6.01059511e-07 4.99960722 6.01090728e-07 4.99799758 6.01143656e-07 4.99699984 6.01199398e-07 5.02510852 6.01276452e-07 4.95223975 6.01342062e-07 2.70342682 6.01411951e-07 0.0431011932 6.01487979e-07 0.0413288898
+ 6.01566956e-07 -0.0198570509 6.01643585e-07 0.0200526747 6.01743585e-07 -0.0178801195 6.01843585e-07 0.0163673972 6.01943585e-07 -0.0148974057 6.02043585e-07 0.0136306143 6.02143585e-07 -0.0124132097 6.02243585e-07 0.0113552946
+ 6.02343585e-07 -0.0103461822 6.02443585e-07 0.0094630689 6.02543585e-07 -0.00862578629 6.02643585e-07 0.00788868402 6.02743585e-07 -0.00719330222 6.02843585e-07 0.00657807192 6.02943585e-07 -0.006000042 6.03043585e-07 0.00548651241
+ 6.03143585e-07 -0.00500567123 6.03243585e-07 0.00457700773 6.03343585e-07 -0.00417676053 6.03443585e-07 0.00381891884 6.03543585e-07 -0.0034855792 6.03643585e-07 0.00318684373 6.03743585e-07 -0.00290910243 6.03843585e-07 0.00265969964
+ 6.03943585e-07 -0.00242819624 6.04043585e-07 0.00221997183 6.04143585e-07 -0.00202694784 6.04243585e-07 0.00185309768 6.04343585e-07 -0.00169211461 6.04443585e-07 0.00154696059 6.04543585e-07 -0.00141266991 6.04643585e-07 0.00129147307
+ 6.04743585e-07 -0.00117942793 6.04843585e-07 0.00107823278 6.04943585e-07 -0.000984733296 6.05043585e-07 0.000900238043 6.05143585e-07 -0.000822203994 6.05243585e-07 0.000751652326 6.05343585e-07 -0.000684967497 6.05443585e-07 0.000628009411
+ 6.05543585e-07 -0.000573313512 6.05643585e-07 0.000524119197 6.05743585e-07 -0.000478719923 6.05843585e-07 0.000437643874 6.05943585e-07 -0.000399739745 6.06043585e-07 0.000365442996 6.06143585e-07 -0.000333794097 6.06243585e-07 0.00030515815
+ 6.06343585e-07 -0.000278730355 6.06443585e-07 0.000254821376 6.06543585e-07 -0.00023159652 6.06643585e-07 0.000212980054 6.06743585e-07 -0.000193420857 6.06843585e-07 0.000177921478 6.06943585e-07 -0.000161548089 6.07043585e-07 0.000149658205
+ 6.07143585e-07 -0.000134776618 6.07243585e-07 0.000124935858 6.07343585e-07 -0.000112502013 6.07443585e-07 0.00010430023 6.07543585e-07 -9.39128182e-05 6.07643585e-07 8.7076031e-05 6.07743585e-07 -7.83977713e-05 6.07843585e-07 7.26984165e-05
+ 6.07943585e-07 -6.54475826e-05 6.08043585e-07 6.06963617e-05 6.08143585e-07 -5.46376243e-05 6.08243585e-07 5.06769633e-05 6.08343585e-07 -4.56137591e-05 6.08443585e-07 4.23124246e-05 6.08543585e-07 -3.80805791e-05 6.08643585e-07 3.53292281e-05
+ 6.08743585e-07 -3.1791625e-05 6.08843585e-07 2.9499122e-05 6.08943585e-07 -2.65412486e-05 6.09043585e-07 2.46316109e-05 6.09143585e-07 -2.21578353e-05 6.09243585e-07 2.05676984e-05 6.09343585e-07 -1.84981586e-05 6.09443585e-07 1.71746699e-05
+ 6.09543585e-07 -1.5442675e-05 6.09643585e-07 1.43417422e-05 6.09743585e-07 -1.28916015e-05 6.09843585e-07 1.19764355e-05 6.09943585e-07 -1.07616446e-05 6.10043585e-07 1.00015461e-05 6.10143585e-07 -8.98327234e-06 6.10243585e-07 8.35262224e-06
+ 6.10343585e-07 -7.49844226e-06 6.10443585e-07 6.97585964e-06 6.10543585e-07 -6.25869755e-06 6.10643585e-07 5.82633423e-06 6.10743585e-07 -5.22358013e-06 6.10843585e-07 4.86653702e-06 6.10943585e-07 -4.35931147e-06 6.11043585e-07 4.06515128e-06
+ 6.11143585e-07 -3.63768999e-06 6.11243585e-07 3.39603008e-06 6.11343585e-07 -3.03517004e-06 6.11443585e-07 2.8373427e-06 6.11543585e-07 -2.53209303e-06 6.11643585e-07 2.37085708e-06 6.11743585e-07 -2.11203389e-06 6.11843585e-07 1.98135588e-06
+ 6.11943585e-07 -1.76130989e-06 6.12043585e-07 1.65614584e-06 6.12143585e-07 -1.46847298e-06 6.12243585e-07 1.38460953e-06 6.12343585e-07 -1.22396639e-06 6.12443585e-07 1.15788736e-06 6.12543585e-07 -1.01981312e-06 6.12643585e-07 9.68583023e-07
+ 6.12743585e-07 -8.49353044e-07 6.12843585e-07 8.10520995e-07 6.12943585e-07 -7.07025355e-07 6.13043585e-07 6.78545058e-07 6.13143585e-07 -5.88187152e-07 6.13243585e-07 5.68350126e-07 6.13343585e-07 -4.88961596e-07 6.13443585e-07 4.76341167e-07
+ 6.13543585e-07 -4.06111844e-07 6.13643585e-07 3.9951709e-07 6.13743585e-07 -3.3693541e-07 6.13843585e-07 3.35371832e-07 6.13943585e-07 -2.79175661e-07 6.14043585e-07 2.81812899e-07 6.14143585e-07 -2.30948406e-07 6.14243585e-07 2.37093157e-07
+ 6.14343585e-07 -1.90680431e-07 6.14443585e-07 1.99753817e-07 6.14543585e-07 -1.57058162e-07 6.14643585e-07 1.68576846e-07 6.14743585e-07 -1.28984815e-07 6.14843585e-07 1.4254523e-07 6.14943585e-07 -1.05544617e-07 6.15043585e-07 1.20809799e-07
+ 6.15143585e-07 -8.59729299e-08 6.15243585e-07 1.0266153e-07 6.15343585e-07 -6.96340728e-08 6.15443585e-07 8.75136771e-08 6.15543585e-07 -5.59972485e-08 6.15643585e-07 7.48717104e-08 6.15743585e-07 -4.46163239e-08 6.15843585e-07 6.43210656e-08
+ 6.15943585e-07 -3.51181102e-08 6.16043585e-07 5.55157795e-08 6.16143585e-07 -2.71911567e-08 6.16243585e-07 4.81671263e-08 6.16343585e-07 -2.05755379e-08 6.16443585e-07 4.2034142e-08 6.16543585e-07 -1.50403401e-08 6.16643585e-07 3.69030002e-08
+ 6.16743585e-07 -1.04355916e-08 6.16843585e-07 3.26339482e-08 6.16943585e-07 -6.59228286e-09 6.17043585e-07 2.90710201e-08 6.17143585e-07 -3.38468512e-09 6.17243585e-07 2.60974314e-08 6.17343585e-07 -7.07655962e-10 6.17443585e-07 2.36157065e-08
+ 6.17543585e-07 1.52656238e-09 6.17643585e-07 2.15643591e-08 6.17743585e-07 3.37429326e-09 6.17843585e-07 1.9875483e-08 6.17943585e-07 4.89591384e-09 6.18043585e-07 1.84846782e-08 6.18143585e-07 6.14898488e-09 6.18243585e-07 1.73393336e-08
+ 6.18343585e-07 7.1809042e-09 6.18443585e-07 1.63961285e-08 6.18543585e-07 8.03070202e-09 6.18643585e-07 1.56193889e-08 6.18743585e-07 8.730519e-09 6.18843585e-07 1.48828709e-08 6.18943585e-07 9.29306102e-09 6.19043585e-07 1.43671892e-08
+ 6.19143585e-07 9.76114514e-09 6.19243585e-07 1.39422636e-08 6.19343585e-07 1.01468814e-08 6.19443585e-07 1.35921051e-08 6.19543585e-07 1.04647404e-08 6.19643585e-07 1.33035664e-08 6.19743585e-07 1.07266619e-08 6.19843585e-07 1.30658055e-08
+ 6.19943585e-07 1.09424891e-08 6.20043585e-07 1.2869888e-08 6.20143585e-07 1.11203324e-08 6.20243585e-07 1.27084505e-08 6.20343585e-07 1.12668762e-08 6.20443585e-07 1.25754253e-08 6.20543585e-07 1.13876285e-08 6.20643585e-07 1.24658125e-08
+ 6.20743585e-07 1.14871282e-08 6.20843585e-07 1.23754922e-08 6.20943585e-07 1.15691149e-08 6.21043585e-07 1.23010691e-08 6.21143585e-07 1.16366712e-08 6.21243585e-07 1.22397455e-08 6.21343585e-07 1.16923362e-08 6.21443585e-07 1.2189216e-08
+ 6.21543585e-07 1.17382027e-08 6.21643585e-07 1.2147581e-08 6.21743585e-07 1.17759953e-08 6.21843585e-07 1.21132755e-08 6.21943585e-07 1.18071351e-08 6.22043585e-07 1.20850087e-08 6.22143585e-07 1.18327929e-08 6.22243585e-07 1.20617188e-08
+ 6.22343585e-07 1.18539331e-08 6.22443585e-07 1.20425292e-08 6.22543585e-07 1.18713516e-08 6.22643585e-07 1.20267179e-08 6.22743585e-07 1.18857028e-08 6.22843585e-07 1.20136909e-08 6.22943585e-07 1.18975271e-08 6.23043585e-07 1.20029576e-08
+ 6.23143585e-07 1.19072691e-08 6.23243585e-07 1.19941146e-08 6.23343585e-07 1.19152952e-08 6.23443585e-07 1.19868294e-08 6.23543585e-07 1.19219075e-08 6.23643585e-07 1.1980827e-08 6.23743585e-07 1.19273553e-08 6.23843585e-07 1.1975882e-08
+ 6.23943585e-07 1.19318434e-08 6.24043585e-07 1.19718084e-08 6.24143585e-07 1.19355402e-08 6.24243585e-07 1.19684525e-08 6.24343585e-07 1.1938586e-08 6.24443585e-07 1.19656882e-08 6.24543585e-07 1.19410948e-08 6.24643585e-07 1.19634108e-08
+ 6.24743585e-07 1.19431612e-08 6.24843585e-07 1.19615351e-08 6.24943585e-07 1.19448633e-08 6.25043585e-07 1.19599901e-08 6.25143585e-07 1.19462654e-08 6.25243585e-07 1.19587172e-08 6.25343585e-07 1.19474203e-08 6.25443585e-07 1.19576688e-08
+ 6.25543585e-07 1.1948371e-08 6.25643585e-07 1.19568059e-08 6.25743585e-07 1.19491541e-08 6.25843585e-07 1.19560951e-08 6.25943585e-07 1.19497992e-08 6.26043585e-07 1.19555095e-08 6.26143585e-07 1.19503302e-08 6.26243585e-07 1.19550275e-08
+ 6.26343585e-07 1.19507671e-08 6.26443585e-07 1.1954631e-08 6.26543585e-07 1.1951127e-08 6.26643585e-07 1.19543042e-08 6.26743585e-07 1.19514233e-08 6.26843585e-07 1.19540354e-08 6.26943585e-07 1.19516671e-08 6.27043585e-07 1.19538139e-08
+ 6.27143585e-07 1.19518674e-08 6.27243585e-07 1.19536314e-08 6.27343585e-07 1.19520328e-08 6.27443585e-07 1.19534817e-08 6.27543585e-07 1.19521685e-08 6.27643585e-07 1.19533584e-08 6.27743585e-07 1.19522803e-08 6.27843585e-07 1.19532566e-08
+ 6.27943585e-07 1.19523721e-08 6.28043585e-07 1.19531736e-08 6.28143585e-07 1.19524477e-08 6.28243585e-07 1.19531047e-08 6.28343585e-07 1.19525098e-08 6.28443585e-07 1.19530486e-08 6.28543585e-07 1.19525605e-08 6.28643585e-07 1.19530018e-08
+ 6.28743585e-07 1.19526027e-08 6.28843585e-07 1.19529638e-08 6.28943585e-07 1.19526368e-08 6.29043585e-07 1.19529326e-08 6.29143585e-07 1.19526652e-08 6.29243585e-07 1.19529066e-08 6.29343585e-07 1.19526883e-08 6.29443585e-07 1.19528853e-08
+ 6.29543585e-07 1.19527075e-08 6.29643585e-07 1.19528683e-08 6.29743585e-07 1.19527231e-08 6.29843585e-07 1.19528538e-08 6.29943585e-07 1.19527358e-08 6.30043585e-07 1.19528424e-08 6.30143585e-07 1.19527458e-08 6.30243585e-07 1.19528328e-08
+ 6.30343585e-07 1.19527545e-08 6.30443585e-07 1.19528251e-08 6.30543585e-07 1.19527617e-08 6.30643585e-07 1.19528185e-08 6.30743585e-07 1.19527671e-08 6.30843585e-07 1.19528134e-08 6.30943585e-07 1.19527717e-08 6.31043585e-07 1.1952809e-08
+ 6.31143585e-07 1.19527757e-08 6.31243585e-07 1.19528053e-08 6.31343585e-07 1.19527789e-08 6.31443585e-07 1.19528027e-08 6.31543585e-07 1.19527812e-08 6.31643585e-07 1.19528004e-08 6.31743585e-07 1.19527832e-08 6.31843585e-07 1.19527984e-08
+ 6.31943585e-07 1.1952785e-08 6.32043585e-07 1.19527969e-08 6.32143585e-07 1.19527859e-08 6.32243585e-07 1.19527958e-08 6.32343585e-07 1.19527871e-08 6.32443585e-07 1.19527946e-08 6.32543585e-07 1.19527879e-08 6.32643585e-07 1.1952794e-08
+ 6.32743585e-07 1.19527884e-08 6.32843585e-07 1.1952793e-08 6.32943585e-07 1.19527891e-08 6.33043585e-07 1.19527925e-08 6.33143585e-07 1.19527895e-08 6.33243585e-07 1.19527919e-08 6.33343585e-07 1.19527899e-08 6.33443585e-07 1.19527917e-08
+ 6.33543585e-07 1.19527901e-08 6.33643585e-07 1.19527914e-08 6.33743585e-07 1.19527905e-08 6.33843585e-07 1.19527909e-08 6.33943585e-07 1.19527905e-08 6.34043585e-07 1.19527909e-08 6.34143585e-07 1.19527906e-08 6.34243585e-07 1.19527909e-08
+ 6.34343585e-07 1.19527906e-08 6.34443585e-07 1.19527908e-08 6.34543585e-07 1.19527906e-08 6.34643585e-07 1.19527906e-08 6.34743585e-07 1.19527907e-08 6.34843585e-07 1.19527905e-08 6.34943585e-07 1.19527906e-08 6.35043585e-07 1.19527905e-08
+ 6.35143585e-07 1.19527906e-08 6.35243585e-07 1.19527903e-08 6.35343585e-07 1.19527907e-08 6.35443585e-07 1.195279e-08 6.35543585e-07 1.19527907e-08 6.35643585e-07 1.19527902e-08 6.35743585e-07 1.19527905e-08 6.35843585e-07 1.195279e-08
+ 6.35943585e-07 1.19527905e-08 6.36043585e-07 1.19527903e-08 6.36143585e-07 1.19527903e-08 6.36243585e-07 1.19527904e-08 6.36343585e-07 1.19527902e-08 6.36443585e-07 1.19527901e-08 6.36543585e-07 1.19527905e-08 6.36643585e-07 1.19527901e-08
+ 6.36743585e-07 1.19527898e-08 6.36843585e-07 1.19527903e-08 6.36943585e-07 1.195279e-08 6.37043585e-07 1.195279e-08 6.37143585e-07 1.19527901e-08 6.37243585e-07 1.19527901e-08 6.37343585e-07 1.19527902e-08 6.37443585e-07 1.19527899e-08
+ 6.37543585e-07 1.19527901e-08 6.37643585e-07 1.19527899e-08 6.37743585e-07 1.19527904e-08 6.37843585e-07 1.19527895e-08 6.37943585e-07 1.19527903e-08 6.38043585e-07 1.19527898e-08 6.38143585e-07 1.19527903e-08 6.38243585e-07 1.19527899e-08
+ 6.38343585e-07 1.19527901e-08 6.38443585e-07 1.19527899e-08 6.38543585e-07 1.195279e-08 6.38643585e-07 1.19527898e-08 6.38743585e-07 1.19527902e-08 6.38843585e-07 1.19527895e-08 6.38943585e-07 1.19527901e-08 6.39043585e-07 1.19527896e-08
+ 6.39143585e-07 1.19527901e-08 6.39243585e-07 1.19527898e-08 6.39343585e-07 1.195279e-08 6.39443585e-07 1.19527898e-08 6.39543585e-07 1.19527901e-08 6.39643585e-07 1.19527897e-08 6.39743585e-07 1.195279e-08 6.39843585e-07 1.19527897e-08
+ 6.39943585e-07 1.19527898e-08 6.40043585e-07 1.19527895e-08 6.40143585e-07 1.19527901e-08 6.40243585e-07 1.19527892e-08 6.40343585e-07 1.19527899e-08 6.40443585e-07 1.19527897e-08 6.40543585e-07 1.195279e-08 6.40643585e-07 1.19527896e-08
+ 6.40743585e-07 1.19527899e-08 6.40843585e-07 1.19527898e-08 6.40943585e-07 1.19527896e-08 6.41043585e-07 1.19527895e-08 6.41143585e-07 1.19527898e-08 6.41243585e-07 1.19527896e-08 6.41343585e-07 1.19527898e-08 6.41443585e-07 1.19527896e-08
+ 6.41543585e-07 1.19527898e-08 6.41643585e-07 1.19527894e-08 6.41743585e-07 1.19527896e-08 6.41843585e-07 1.19527892e-08 6.41943585e-07 1.19527895e-08 6.42043585e-07 1.19527895e-08 6.42143585e-07 1.19527898e-08 6.42243585e-07 1.19527892e-08
+ 6.42343585e-07 1.19527897e-08 6.42443585e-07 1.19527895e-08 6.42543585e-07 1.19527896e-08 6.42643585e-07 1.19527894e-08 6.42743585e-07 1.19527894e-08 6.42843585e-07 1.19527895e-08 6.42943585e-07 1.19527894e-08 6.43043585e-07 1.19527896e-08
+ 6.43143585e-07 1.19527894e-08 6.43243585e-07 1.19527894e-08 6.43343585e-07 1.19527896e-08 6.43443585e-07 1.19527895e-08 6.43543585e-07 1.19527896e-08 6.43643585e-07 1.19527893e-08 6.43743585e-07 1.19527893e-08 6.43843585e-07 1.19527893e-08
+ 6.43943585e-07 1.19527894e-08 6.44043585e-07 1.19527893e-08 6.44143585e-07 1.19527895e-08 6.44243585e-07 1.19527895e-08 6.44343585e-07 1.19527895e-08 6.44443585e-07 1.19527894e-08 6.44543585e-07 1.19527895e-08 6.44643585e-07 1.19527896e-08
+ 6.44743585e-07 1.19527894e-08 6.44843585e-07 1.19527893e-08 6.44943585e-07 1.19527892e-08 6.45043585e-07 1.19527894e-08 6.45143585e-07 1.19527893e-08 6.45243585e-07 1.19527891e-08 6.45343585e-07 1.19527895e-08 6.45443585e-07 1.19527893e-08
+ 6.45543585e-07 1.19527891e-08 6.45643585e-07 1.19527892e-08 6.45743585e-07 1.19527894e-08 6.45843585e-07 1.19527895e-08 6.45943585e-07 1.19527892e-08 6.46043585e-07 1.19527891e-08 6.46143585e-07 1.19527893e-08 6.46243585e-07 1.19527893e-08
+ 6.46343585e-07 1.19527892e-08 6.46443585e-07 1.19527893e-08 6.46543585e-07 1.19527892e-08 6.46643585e-07 1.19527894e-08 6.46743585e-07 1.19527892e-08 6.46843585e-07 1.19527893e-08 6.46943585e-07 1.19527891e-08 6.47043585e-07 1.19527893e-08
+ 6.47143585e-07 1.1952789e-08 6.47243585e-07 1.19527891e-08 6.47343585e-07 1.19527891e-08 6.47443585e-07 1.19527895e-08 6.47543585e-07 1.19527889e-08 6.47643585e-07 1.19527893e-08 6.47743585e-07 1.19527891e-08 6.47843585e-07 1.19527892e-08
+ 6.47943585e-07 1.1952789e-08 6.48043585e-07 1.19527893e-08 6.48143585e-07 1.1952789e-08 6.48243585e-07 1.19527893e-08 6.48343585e-07 1.19527888e-08 6.48443585e-07 1.19527895e-08 6.48543585e-07 1.19527888e-08 6.48643585e-07 1.19527892e-08
+ 6.48743585e-07 1.19527889e-08 6.48843585e-07 1.19527892e-08 6.48943585e-07 1.19527891e-08 6.49043585e-07 1.19527893e-08 6.49143585e-07 1.1952789e-08 6.49243585e-07 1.19527893e-08 6.49343585e-07 1.19527887e-08 6.49443585e-07 1.19527891e-08
+ 6.49543585e-07 1.19527888e-08 6.49643585e-07 1.19527893e-08 6.49743585e-07 1.1952789e-08 6.49843585e-07 1.19527894e-08 6.49943585e-07 1.19527888e-08 6.50043585e-07 1.19527892e-08 6.50143585e-07 1.19527889e-08 6.50243585e-07 1.19527893e-08
+ 6.50343585e-07 1.19527889e-08 6.50443585e-07 1.19527895e-08 6.50543585e-07 1.19527889e-08 6.50643585e-07 1.19527894e-08 6.50743585e-07 1.19527887e-08 6.50843585e-07 1.19527894e-08 6.50943585e-07 1.19527887e-08 6.51e-07 1.19527896e-08
+ 6.5101e-07 1.19387339e-08 6.5103e-07 1.20209579e-08 6.5107e-07 1.18456563e-08 6.5115e-07 1.20751985e-08 6.5125e-07 1.18257281e-08 6.5135e-07 1.20743629e-08 6.5145e-07 1.18466579e-08 6.5155e-07 1.2036145e-08
+ 6.5165e-07 1.18950759e-08 6.5175e-07 1.19816166e-08 6.5185e-07 1.19573518e-08 6.51930828e-07 1.29898242e-07 6.52e-07 1.68693818e-06 6.52008608e-07 -4.63455704e-06 6.52025825e-07 -7.9808205e-06 6.52060258e-07 1.5061975e-06
+ 6.52106181e-07 1.0973022e-05 6.52150081e-07 -1.19545368e-05 6.52198026e-07 8.69407648e-06 6.5225538e-07 -7.92726691e-06 6.52312019e-07 6.0886179e-06 6.52404231e-07 -4.35191802e-06 6.52504231e-07 2.87067141e-06 6.52604231e-07 -1.60647351e-06
+ 6.52704231e-07 7.0938315e-07 6.52804231e-07 6.21050554e-08 6.52904231e-07 -6.67617034e-07 6.53004231e-07 1.2280794e-06 6.53104231e-07 -1.66857258e-06 6.53204231e-07 2.08522619e-06 6.53304231e-07 -2.39320129e-06 6.53404231e-07 2.68781493e-06
+ 6.53504231e-07 -2.88197065e-06 6.53604231e-07 3.07280994e-06 6.53704231e-07 -3.17200642e-06 6.53804231e-07 3.2781936e-06 6.53904231e-07 -3.30170758e-06 6.54004231e-07 3.34196797e-06 6.54104231e-07 -3.30788027e-06 6.54204231e-07 3.2991216e-06
+ 6.54304231e-07 -3.2232367e-06 6.54404231e-07 3.17983294e-06 6.54504231e-07 -3.07526771e-06 6.54604231e-07 3.00890095e-06 6.54704231e-07 -2.88611918e-06 6.54804231e-07 2.80595288e-06 6.54904231e-07 -2.67303462e-06 6.55004231e-07 2.58603942e-06
+ 6.55104231e-07 -2.44904115e-06 6.55204231e-07 2.36036454e-06 6.55304231e-07 -2.22368841e-06 6.55404231e-07 2.13700757e-06 6.55504231e-07 -2.00373963e-06 6.55604231e-07 1.92157875e-06 6.55704231e-07 -1.79378453e-06 6.55804231e-07 1.71778029e-06
+ 6.55904231e-07 -1.59674487e-06 6.56004231e-07 1.52786046e-06 6.56104231e-07 -1.41428355e-06 6.56204231e-07 1.3529841e-06 6.56304231e-07 -1.24713754e-06 6.56404231e-07 1.19352802e-06 6.56504231e-07 -1.09537836e-06 6.56604231e-07 1.04931085e-06
+ 6.56704231e-07 -9.58614228e-07 6.56804231e-07 9.19769769e-07 6.56904231e-07 -8.36142431e-07 6.57004231e-07 8.04091186e-07 6.57104231e-07 -7.27063187e-07 6.57204231e-07 7.01312281e-07 6.57304231e-07 -6.30369486e-07 6.57404231e-07 6.10398102e-07
+ 6.57504231e-07 -5.45011509e-07 6.57604231e-07 5.30294844e-07 6.57704231e-07 -4.69940202e-07 6.57804231e-07 4.59965237e-07 6.57904231e-07 -4.04136037e-07 6.58004231e-07 3.98412181e-07 6.58104231e-07 -3.46628439e-07 6.58204231e-07 3.44694536e-07
+ 6.58304231e-07 -2.96508308e-07 6.58404231e-07 2.97936752e-07 6.58504231e-07 -2.52935085e-07 6.58604231e-07 2.57333733e-07 6.58704231e-07 -2.1513933e-07 6.58804231e-07 2.22150053e-07 6.58904231e-07 -1.82418412e-07 6.59004231e-07 1.9171647e-07
+ 6.59104231e-07 -1.54139153e-07 6.59204231e-07 1.65436835e-07 6.59304231e-07 -1.29741724e-07 6.59404231e-07 1.42784958e-07 6.59504231e-07 -1.08731077e-07 6.59604231e-07 1.23294537e-07 6.59704231e-07 -9.06683015e-08 6.59804231e-07 1.06552593e-07
+ 6.59904231e-07 -7.5165328e-08 6.60004231e-07 9.2194631e-08 6.60104231e-07 -6.1880455e-08 6.60204231e-07 7.99012531e-08 6.60304231e-07 -5.0515895e-08 6.60404231e-07 6.93947395e-08 6.60504231e-07 -4.0813082e-08 6.60604231e-07 6.04320326e-08
+ 6.60704231e-07 -3.25414544e-08 6.60804231e-07 5.27962643e-08 6.60904231e-07 -2.54989315e-08 6.61004231e-07 4.62991432e-08 6.61104231e-07 -1.95102628e-08 6.61204231e-07 4.07775697e-08 6.61304231e-07 -1.44238236e-08 6.61404231e-07 3.60905903e-08
+ 6.61504231e-07 -1.01087194e-08 6.61604231e-07 3.21166457e-08 6.61704231e-07 -6.45216383e-09 6.61804231e-07 2.87510622e-08 6.61904231e-07 -3.35709155e-09 6.62004231e-07 2.59038328e-08 6.62104231e-07 -7.40147582e-10 6.62204231e-07 2.34977897e-08
+ 6.62304231e-07 1.46047882e-09 6.62404231e-07 2.14846645e-08 6.62504231e-07 3.2971606e-09 6.62604231e-07 1.98091944e-08 6.62704231e-07 4.82515061e-09 6.62804231e-07 1.84160882e-08 6.62904231e-07 6.0949224e-09 6.63004231e-07 1.72590653e-08
+ 6.63104231e-07 7.14889656e-09 6.63204231e-07 1.62992532e-08 6.63304231e-07 8.02268554e-09 6.63404231e-07 1.55040344e-08 6.63504231e-07 8.74615705e-09 6.63604231e-07 1.4846065e-08 6.63704231e-07 9.34433925e-09 6.63804231e-07 1.43024406e-08
+ 6.63904231e-07 9.83818962e-09 6.64004231e-07 1.38540378e-08 6.64104231e-07 1.0245185e-08 6.64204231e-07 1.34848201e-08 6.64304231e-07 1.0579713e-08 6.64404231e-07 1.31818535e-08 6.64504231e-07 1.08542379e-08 6.64604231e-07 1.293309e-08
+ 6.64704231e-07 1.10795435e-08 6.64804231e-07 1.27292155e-08 6.64904231e-07 1.12638395e-08 6.65004231e-07 1.25627463e-08 6.65104231e-07 1.14141357e-08 6.65204231e-07 1.24270858e-08 6.65304231e-07 1.15365053e-08 6.65404231e-07 1.23168959e-08
+ 6.65504231e-07 1.16355321e-08 6.65604231e-07 1.22280072e-08 6.65704231e-07 1.17152599e-08 6.65804231e-07 1.21565573e-08 6.65904231e-07 1.17792245e-08 6.66004231e-07 1.20993641e-08 6.66104231e-07 1.18302937e-08 6.66204231e-07 1.20538322e-08
+ 6.66304231e-07 1.18708183e-08 6.66404231e-07 1.20178358e-08 6.66504231e-07 1.19027244e-08 6.66604231e-07 1.1989619e-08 6.66704231e-07 1.19276164e-08 6.66804231e-07 1.19676439e-08 6.66904231e-07 1.1946949e-08 6.67004231e-07 1.19508727e-08
+ 6.67104231e-07 1.19614316e-08 6.67204231e-07 1.19383222e-08 6.67304231e-07 1.19722685e-08 6.67404231e-07 1.19290236e-08 6.67504231e-07 1.19801835e-08 6.67604231e-07 1.19223501e-08 6.67704231e-07 1.19857468e-08 6.67804231e-07 1.19177778e-08
+ 6.67904231e-07 1.19894366e-08 6.68004231e-07 1.19148714e-08 6.68104231e-07 1.19916496e-08 6.68204231e-07 1.19132703e-08 6.68304231e-07 1.19927119e-08 6.68404231e-07 1.19126811e-08 6.68504231e-07 1.19929032e-08 6.68604231e-07 1.19128184e-08
+ 6.68704231e-07 1.19924515e-08 6.68804231e-07 1.19135801e-08 6.68904231e-07 1.19914317e-08 6.69004231e-07 1.19147993e-08 6.69104231e-07 1.19900508e-08 6.69204231e-07 1.19163127e-08 6.69304231e-07 1.19884329e-08 6.69404231e-07 1.19180127e-08
+ 6.69504231e-07 1.19866634e-08 6.69604231e-07 1.19198411e-08 6.69704231e-07 1.19847903e-08 6.69804231e-07 1.19217443e-08 6.69904231e-07 1.19828696e-08 6.70004231e-07 1.19236705e-08 6.70104231e-07 1.19809474e-08 6.70204231e-07 1.19255819e-08
+ 6.70304231e-07 1.19790537e-08 6.70404231e-07 1.19274518e-08 6.70504231e-07 1.19772121e-08 6.70604231e-07 1.19292611e-08 6.70704231e-07 1.19754386e-08 6.70804231e-07 1.19309964e-08 6.70904231e-07 1.19737437e-08 6.71004231e-07 1.19326492e-08
+ 6.71104231e-07 1.19721343e-08 6.71204231e-07 1.19342136e-08 6.71304231e-07 1.19706149e-08 6.71404231e-07 1.19356878e-08 6.71504231e-07 1.19691864e-08 6.71604231e-07 1.19370708e-08 6.71704231e-07 1.1967849e-08 6.71804231e-07 1.1938363e-08
+ 6.71904231e-07 1.19666018e-08 6.72004231e-07 1.19395658e-08 6.72104231e-07 1.19654424e-08 6.72204231e-07 1.19406827e-08 6.72304231e-07 1.19643672e-08 6.72404231e-07 1.19417168e-08 6.72504231e-07 1.19633727e-08 6.72604231e-07 1.19426723e-08
+ 6.72704231e-07 1.19624554e-08 6.72804231e-07 1.19435533e-08 6.72904231e-07 1.19616097e-08 6.73004231e-07 1.1944364e-08 6.73104231e-07 1.19608331e-08 6.73204231e-07 1.19451072e-08 6.73304231e-07 1.19601215e-08 6.73404231e-07 1.19457902e-08
+ 6.73504231e-07 1.19594654e-08 6.73604231e-07 1.19464193e-08 6.73704231e-07 1.19588636e-08 6.73804231e-07 1.19469944e-08 6.73904231e-07 1.19583144e-08 6.74004231e-07 1.19475189e-08 6.74104231e-07 1.19578135e-08 6.74204231e-07 1.1947997e-08
+ 6.74304231e-07 1.19573573e-08 6.74404231e-07 1.19484327e-08 6.74504231e-07 1.19569411e-08 6.74604231e-07 1.19488295e-08 6.74704231e-07 1.19565626e-08 6.74804231e-07 1.19491909e-08 6.74904231e-07 1.19562178e-08 6.75004231e-07 1.19495197e-08
+ 6.75104231e-07 1.19559043e-08 6.75204231e-07 1.19498187e-08 6.75304231e-07 1.19556191e-08 6.75404231e-07 1.19500906e-08 6.75504231e-07 1.19553597e-08 6.75604231e-07 1.19503383e-08 6.75704231e-07 1.19551232e-08 6.75804231e-07 1.19505643e-08
+ 6.75904231e-07 1.19549075e-08 6.76004231e-07 1.19507697e-08 6.76104231e-07 1.19547121e-08 6.76204231e-07 1.19509559e-08 6.76304231e-07 1.19545346e-08 6.76404231e-07 1.19511245e-08 6.76504231e-07 1.19543743e-08 6.76604231e-07 1.19512774e-08
+ 6.76704231e-07 1.19542286e-08 6.76804231e-07 1.19514159e-08 6.76904231e-07 1.19540967e-08 6.77004231e-07 1.1951542e-08 6.77104231e-07 1.19539768e-08 6.77204231e-07 1.19516558e-08 6.77304231e-07 1.1953868e-08 6.77404231e-07 1.19517598e-08
+ 6.77504231e-07 1.1953769e-08 6.77604231e-07 1.19518539e-08 6.77704231e-07 1.19536795e-08 6.77804231e-07 1.19519395e-08 6.77904231e-07 1.19535977e-08 6.78004231e-07 1.19520173e-08 6.78104231e-07 1.19535235e-08 6.78204231e-07 1.19520877e-08
+ 6.78304231e-07 1.19534563e-08 6.78404231e-07 1.19521518e-08 6.78504231e-07 1.19533954e-08 6.78604231e-07 1.195221e-08 6.78704231e-07 1.19533397e-08 6.78804231e-07 1.19522632e-08 6.78904231e-07 1.19532891e-08 6.79004231e-07 1.19523112e-08
+ 6.79104231e-07 1.19532433e-08 6.79204231e-07 1.1952355e-08 6.79304231e-07 1.19532014e-08 6.79404231e-07 1.19523948e-08 6.79504231e-07 1.19531634e-08 6.79604231e-07 1.1952431e-08 6.79704231e-07 1.19531292e-08 6.79804231e-07 1.19524639e-08
+ 6.79904231e-07 1.19530979e-08 6.80004231e-07 1.19524936e-08 6.80104231e-07 1.19530694e-08 6.80204231e-07 1.19525209e-08 6.80304231e-07 1.19530436e-08 6.80404231e-07 1.19525454e-08 6.80504231e-07 1.19530202e-08 6.80604231e-07 1.19525678e-08
+ 6.80704231e-07 1.19529989e-08 6.80804231e-07 1.19525882e-08 6.80904231e-07 1.19529795e-08 6.81004231e-07 1.19526065e-08 6.81104231e-07 1.1952962e-08 6.81204231e-07 1.19526236e-08 6.81304231e-07 1.19529458e-08 6.81404231e-07 1.19526388e-08
+ 6.81504231e-07 1.19529312e-08 6.81604231e-07 1.19526528e-08 6.81704231e-07 1.19529178e-08 6.81804231e-07 1.19526654e-08 6.81904231e-07 1.19529058e-08 6.82004231e-07 1.19526766e-08 6.82104231e-07 1.19528951e-08 6.82204231e-07 1.19526871e-08
+ 6.82304231e-07 1.19528849e-08 6.82404231e-07 1.19526965e-08 6.82504231e-07 1.1952876e-08 6.82604231e-07 1.19527051e-08 6.82704231e-07 1.1952868e-08 6.82804231e-07 1.19527125e-08 6.82904231e-07 1.19528603e-08 6.83004231e-07 1.19527197e-08
+ 6.83104231e-07 1.19528536e-08 6.83204231e-07 1.19527265e-08 6.83304231e-07 1.19528476e-08 6.83404231e-07 1.19527322e-08 6.83504231e-07 1.1952842e-08 6.83604231e-07 1.19527372e-08 6.83704231e-07 1.19528371e-08 6.83804231e-07 1.1952742e-08
+ 6.83904231e-07 1.19528326e-08 6.84004231e-07 1.19527464e-08 6.84104231e-07 1.19528284e-08 6.84204231e-07 1.19527503e-08 6.84304231e-07 1.19528246e-08 6.84404231e-07 1.19527539e-08 6.84504231e-07 1.19528215e-08 6.84604231e-07 1.19527572e-08
+ 6.84704231e-07 1.19528182e-08 6.84804231e-07 1.195276e-08 6.84904231e-07 1.19528154e-08 6.85004231e-07 1.19527629e-08 6.85104231e-07 1.19528129e-08 6.85204231e-07 1.19527651e-08 6.85304231e-07 1.19528105e-08 6.85404231e-07 1.19527676e-08
+ 6.85504231e-07 1.19528084e-08 6.85604231e-07 1.19527695e-08 6.85704231e-07 1.19528063e-08 6.85804231e-07 1.19527714e-08 6.85904231e-07 1.19528047e-08 6.86004231e-07 1.1952773e-08 6.86104231e-07 1.19528031e-08 6.86204231e-07 1.19527745e-08
+ 6.86304231e-07 1.19528017e-08 6.86404231e-07 1.19527759e-08 6.86504231e-07 1.19528006e-08 6.86604231e-07 1.19527768e-08 6.86704231e-07 1.19527992e-08 6.86804231e-07 1.19527781e-08 6.86904231e-07 1.19527984e-08 6.87004231e-07 1.1952779e-08
+ 6.87104231e-07 1.19527973e-08 6.87204231e-07 1.19527801e-08 6.87304231e-07 1.19527965e-08 6.87404231e-07 1.19527808e-08 6.87504231e-07 1.19527956e-08 6.87604231e-07 1.19527814e-08 6.87704231e-07 1.19527948e-08 6.87804231e-07 1.19527823e-08
+ 6.87904231e-07 1.19527944e-08 6.88004231e-07 1.19527827e-08 6.88104231e-07 1.19527936e-08 6.88204231e-07 1.19527833e-08 6.88304231e-07 1.19527931e-08 6.88404231e-07 1.19527838e-08 6.88504231e-07 1.19527926e-08 6.88604231e-07 1.19527842e-08
+ 6.88704231e-07 1.19527925e-08 6.88804231e-07 1.19527845e-08 6.88904231e-07 1.1952792e-08 6.89004231e-07 1.19527847e-08 6.89104231e-07 1.19527917e-08 6.89204231e-07 1.19527851e-08 6.89304231e-07 1.19527916e-08 6.89404231e-07 1.19527854e-08
+ 6.89504231e-07 1.19527913e-08 6.89604231e-07 1.19527858e-08 6.89704231e-07 1.19527906e-08 6.89804231e-07 1.19527862e-08 6.89904231e-07 1.19527904e-08 6.90004231e-07 1.19527864e-08 6.90104231e-07 1.19527904e-08 6.90204231e-07 1.19527867e-08
+ 6.90304231e-07 1.19527899e-08 6.90404231e-07 1.19527869e-08 6.90504231e-07 1.195279e-08 6.90604231e-07 1.1952787e-08 6.90704231e-07 1.19527896e-08 6.90804231e-07 1.19527872e-08 6.90904231e-07 1.19527898e-08 6.91004231e-07 1.19527873e-08
+ 6.91104231e-07 1.19527898e-08 6.91204231e-07 1.19527872e-08 6.91304231e-07 1.19527897e-08 6.91404231e-07 1.19527874e-08 6.91504231e-07 1.19527895e-08 6.91604231e-07 1.19527873e-08 6.91704231e-07 1.19527895e-08 6.91804231e-07 1.19527873e-08
+ 6.91904231e-07 1.19527892e-08 6.92004231e-07 1.19527874e-08 6.92104231e-07 1.19527893e-08 6.92204231e-07 1.19527875e-08 6.92304231e-07 1.19527893e-08 6.92404231e-07 1.19527878e-08 6.92504231e-07 1.19527893e-08 6.92604231e-07 1.19527876e-08
+ 6.92704231e-07 1.19527891e-08 6.92804231e-07 1.19527878e-08 6.92904231e-07 1.19527892e-08 6.93004231e-07 1.19527876e-08 6.93104231e-07 1.19527891e-08 6.93204231e-07 1.1952788e-08 6.93304231e-07 1.1952789e-08 6.93404231e-07 1.19527879e-08
+ 6.93504231e-07 1.1952789e-08 6.93604231e-07 1.19527881e-08 6.93704231e-07 1.19527887e-08 6.93804231e-07 1.1952788e-08 6.93904231e-07 1.19527889e-08 6.94004231e-07 1.19527881e-08 6.94104231e-07 1.19527889e-08 6.94204231e-07 1.19527881e-08
+ 6.94304231e-07 1.19527887e-08 6.94404231e-07 1.19527883e-08 6.94504231e-07 1.19527883e-08 6.94604231e-07 1.19527883e-08 6.94704231e-07 1.19527883e-08 6.94804231e-07 1.19527884e-08 6.94904231e-07 1.19527885e-08 6.95004231e-07 1.19527882e-08
+ 6.95104231e-07 1.19527884e-08 6.95204231e-07 1.19527886e-08 6.95304231e-07 1.19527885e-08 6.95404231e-07 1.19527887e-08 6.95504231e-07 1.19527883e-08 6.95604231e-07 1.19527886e-08 6.95704231e-07 1.19527885e-08 6.95804231e-07 1.19527885e-08
+ 6.95904231e-07 1.19527884e-08 6.96004231e-07 1.19527886e-08 6.96104231e-07 1.19527885e-08 6.96204231e-07 1.19527883e-08 6.96304231e-07 1.19527883e-08 6.96404231e-07 1.19527885e-08 6.96504231e-07 1.19527884e-08 6.96604231e-07 1.19527886e-08
+ 6.96704231e-07 1.19527883e-08 6.96804231e-07 1.19527881e-08 6.96904231e-07 1.19527885e-08 6.97004231e-07 1.19527885e-08 6.97104231e-07 1.19527885e-08 6.97204231e-07 1.19527882e-08 6.97304231e-07 1.19527886e-08 6.97404231e-07 1.19527884e-08
+ 6.97504231e-07 1.19527884e-08 6.97604231e-07 1.19527884e-08 6.97704231e-07 1.19527883e-08 6.97804231e-07 1.19527883e-08 6.97904231e-07 1.19527885e-08 6.98004231e-07 1.19527884e-08 6.98104231e-07 1.19527885e-08 6.98204231e-07 1.19527884e-08
+ 6.98304231e-07 1.19527884e-08 6.98404231e-07 1.19527885e-08 6.98504231e-07 1.19527884e-08 6.98604231e-07 1.19527884e-08 6.98704231e-07 1.19527884e-08 6.98804231e-07 1.19527883e-08 6.98904231e-07 1.19527883e-08 6.99004231e-07 1.19527886e-08
+ 6.99104231e-07 1.19527882e-08 6.99204231e-07 1.19527885e-08 6.99304231e-07 1.19527884e-08 6.99404231e-07 1.19527882e-08 6.99504231e-07 1.19527883e-08 6.99604231e-07 1.19527885e-08 6.99704231e-07 1.19527883e-08 6.99804231e-07 1.19527885e-08
+ 6.99904231e-07 1.19527884e-08 7e-07 1.19527882e-08 7.0001e-07 1.19885671e-08 7.0003e-07 1.17808827e-08 7.0007e-07 1.22180336e-08 7.0015e-07 1.1655688e-08 7.0025e-07 1.22568031e-08 7.0035e-07 1.16606774e-08
+ 7.0045e-07 1.22151902e-08 7.0055e-07 1.17418277e-08 7.0065e-07 1.18107333e-08 7.0075e-07 2.87697415e-08 7.0085e-07 -5.432075e-07 7.00931988e-07 7.32055252e-06 7.01e-07 -4.5908469e-05 7.01008484e-07 -5.04559152e-05
+ 7.01025451e-07 -3.69618015e-05 7.01059385e-07 -3.09903885e-05 7.01090588e-07 0.000242070373 7.01143428e-07 0.000483109234 7.011991e-07 0.00152689372 7.012991e-07 -0.0155867066 7.013991e-07 0.117270425 7.014991e-07 4.30152836
+ 7.01578678e-07 5.13555996 7.01663998e-07 4.92548528 7.01763998e-07 5.04581425 7.01858547e-07 4.97061047 7.01958547e-07 5.01945309 7.02058547e-07 4.98680161 7.02158547e-07 5.00891418 7.02258547e-07 4.99390118
+ 7.02358547e-07 5.00413809 7.02458547e-07 4.99716775 7.02558547e-07 5.00191851 7.02658547e-07 4.99869244 7.02758547e-07 5.00087968 7.02858547e-07 4.99940653 7.02958547e-07 5.00039318 7.03058547e-07 4.99974055
+ 7.03158547e-07 5.0001661 7.03258547e-07 4.9998959 7.03358547e-07 5.00006105 7.03458547e-07 4.99996722 7.03558547e-07 5.00001337 7.03658547e-07 4.99999907 7.03758547e-07 4.99999272 7.03858547e-07 5.00001245
+ 7.03958547e-07 4.99998442 7.04058547e-07 5.00001725 7.04158547e-07 4.99998194 7.04258547e-07 5.00001816 7.04358547e-07 4.99998204 7.04458547e-07 5.00001738 7.04558547e-07 4.99998323 7.04658547e-07 5.00001594
+ 7.04758547e-07 4.9999848 7.04858547e-07 5.00001432 7.04958547e-07 4.99998643 7.05058547e-07 5.00001272 7.05158547e-07 4.99998798 7.05258547e-07 5.00001123 7.05358547e-07 4.9999894 7.05458547e-07 5.00000988
+ 7.05558547e-07 4.99999068 7.05658547e-07 5.00000868 7.05758547e-07 4.99999181 7.05858547e-07 5.00000762 7.05958547e-07 4.99999281 7.06058547e-07 5.00000668 7.06158547e-07 4.99999369 7.06258547e-07 5.00000585
+ 7.06358547e-07 4.99999446 7.06458547e-07 5.00000513 7.06558547e-07 4.99999514 7.06658547e-07 5.00000449 7.06758547e-07 4.99999573 7.06858547e-07 5.00000394 7.06958547e-07 4.99999626 7.07058547e-07 5.00000345
+ 7.07158547e-07 4.99999671 7.07258547e-07 5.00000302 7.07358547e-07 4.99999712 7.07458547e-07 5.00000264 7.07558547e-07 4.99999747 7.07658547e-07 5.00000231 7.07758547e-07 4.99999778 7.07858547e-07 5.00000203
+ 7.07958547e-07 4.99999805 7.08058547e-07 5.00000177 7.08158547e-07 4.99999828 7.08258547e-07 5.00000155 7.08358547e-07 4.99999849 7.08458547e-07 5.00000136 7.08558547e-07 4.99999868 7.08658547e-07 5.00000119
+ 7.08758547e-07 4.99999884 7.08858547e-07 5.00000104 7.08958547e-07 4.99999898 7.09058547e-07 5.0000009 7.09158547e-07 4.9999991 7.09258547e-07 5.00000079 7.09358547e-07 4.99999921 7.09458547e-07 5.00000069
+ 7.09558547e-07 4.9999993 7.09658547e-07 5.0000006 7.09758547e-07 4.99999938 7.09858547e-07 5.00000052 7.09958547e-07 4.99999946 7.10058547e-07 5.00000045 7.10158547e-07 4.99999952 7.10258547e-07 5.0000004
+ 7.10358547e-07 4.99999958 7.10458547e-07 5.00000034 7.10558547e-07 4.99999962 7.10658547e-07 5.0000003 7.10758547e-07 4.99999967 7.10858547e-07 5.00000026 7.10958547e-07 4.99999971 7.11058547e-07 5.00000022
+ 7.11158547e-07 4.99999973 7.11258547e-07 5.00000019 7.11358547e-07 4.99999976 7.11458547e-07 5.00000016 7.11558547e-07 4.99999979 7.11658547e-07 5.00000014 7.11758547e-07 4.99999981 7.11858547e-07 5.00000012
+ 7.11958547e-07 4.99999983 7.12058547e-07 5.0000001 7.12158547e-07 4.99999985 7.12258547e-07 5.00000008 7.12358547e-07 4.99999986 7.12458547e-07 5.00000007 7.12558547e-07 4.99999988 7.12658547e-07 5.00000006
+ 7.12758547e-07 4.99999989 7.12858547e-07 5.00000005 7.12958547e-07 4.9999999 7.13058547e-07 5.00000004 7.13158547e-07 4.99999991 7.13258547e-07 5.00000003 7.13358547e-07 4.99999992 7.13458547e-07 5.00000002
+ 7.13558547e-07 4.99999992 7.13658547e-07 5.00000002 7.13758547e-07 4.99999993 7.13858547e-07 5.00000001 7.13958547e-07 4.99999994 7.14058547e-07 5.0 7.14158547e-07 4.99999994 7.14258547e-07 5.0
+ 7.14358547e-07 4.99999994 7.14458547e-07 5.0 7.14558547e-07 4.99999995 7.14658547e-07 4.99999999 7.14758547e-07 4.99999995 7.14858547e-07 4.99999999 7.14958547e-07 4.99999995 7.15058547e-07 4.99999999
+ 7.15158547e-07 4.99999996 7.15258547e-07 4.99999999 7.15358547e-07 4.99999996 7.15458547e-07 4.99999998 7.15558547e-07 4.99999996 7.15658547e-07 4.99999998 7.15758547e-07 4.99999996 7.15858547e-07 4.99999998
+ 7.15958547e-07 4.99999996 7.16058547e-07 4.99999998 7.16158547e-07 4.99999996 7.16258547e-07 4.99999998 7.16358547e-07 4.99999997 7.16458547e-07 4.99999998 7.16558547e-07 4.99999997 7.16658547e-07 4.99999998
+ 7.16758547e-07 4.99999997 7.16858547e-07 4.99999998 7.16958547e-07 4.99999997 7.17058547e-07 4.99999998 7.17158547e-07 4.99999997 7.17258547e-07 4.99999998 7.17358547e-07 4.99999997 7.17458547e-07 4.99999998
+ 7.17558547e-07 4.99999997 7.17658547e-07 4.99999998 7.17758547e-07 4.99999997 7.17858547e-07 4.99999997 7.17958547e-07 4.99999997 7.18058547e-07 4.99999997 7.18158547e-07 4.99999997 7.18258547e-07 4.99999997
+ 7.18358547e-07 4.99999997 7.18458547e-07 4.99999997 7.18558547e-07 4.99999997 7.18658547e-07 4.99999997 7.18758547e-07 4.99999997 7.18858547e-07 4.99999997 7.18958547e-07 4.99999997 7.19058547e-07 4.99999997
+ 7.19158547e-07 4.99999997 7.19258547e-07 4.99999997 7.19358547e-07 4.99999997 7.19458547e-07 4.99999997 7.19558547e-07 4.99999997 7.19658547e-07 4.99999997 7.19758547e-07 4.99999997 7.19858547e-07 4.99999997
+ 7.19958547e-07 4.99999997 7.20058547e-07 4.99999997 7.20158547e-07 4.99999997 7.20258547e-07 4.99999997 7.20358547e-07 4.99999997 7.20458547e-07 4.99999997 7.20558547e-07 4.99999997 7.20658547e-07 4.99999997
+ 7.20758547e-07 4.99999997 7.20858547e-07 4.99999997 7.20958547e-07 4.99999997 7.21058547e-07 4.99999997 7.21158547e-07 4.99999997 7.21258547e-07 4.99999997 7.21358547e-07 4.99999997 7.21458547e-07 4.99999997
+ 7.21558547e-07 4.99999997 7.21658547e-07 4.99999997 7.21758547e-07 4.99999997 7.21858547e-07 4.99999997 7.21958547e-07 4.99999997 7.22058547e-07 4.99999997 7.22158547e-07 4.99999997 7.22258547e-07 4.99999997
+ 7.22358547e-07 4.99999997 7.22458547e-07 4.99999997 7.22558547e-07 4.99999997 7.22658547e-07 4.99999997 7.22758547e-07 4.99999997 7.22858547e-07 4.99999997 7.22958547e-07 4.99999997 7.23058547e-07 4.99999997
+ 7.23158547e-07 4.99999997 7.23258547e-07 4.99999997 7.23358547e-07 4.99999997 7.23458547e-07 4.99999997 7.23558547e-07 4.99999997 7.23658547e-07 4.99999997 7.23758547e-07 4.99999997 7.23858547e-07 4.99999997
+ 7.23958547e-07 4.99999997 7.24058547e-07 4.99999997 7.24158547e-07 4.99999997 7.24258547e-07 4.99999997 7.24358547e-07 4.99999997 7.24458547e-07 4.99999997 7.24558547e-07 4.99999997 7.24658547e-07 4.99999997
+ 7.24758547e-07 4.99999997 7.24858547e-07 4.99999997 7.24958547e-07 4.99999997 7.25058547e-07 4.99999997 7.25158547e-07 4.99999997 7.25258547e-07 4.99999997 7.25358547e-07 4.99999997 7.25458547e-07 4.99999997
+ 7.25558547e-07 4.99999997 7.25658547e-07 4.99999997 7.25758547e-07 4.99999997 7.25858547e-07 4.99999997 7.25958547e-07 4.99999997 7.26058547e-07 4.99999997 7.26158547e-07 4.99999997 7.26258547e-07 4.99999997
+ 7.26358547e-07 4.99999997 7.26458547e-07 4.99999997 7.26558547e-07 4.99999997 7.26658547e-07 4.99999997 7.26758547e-07 4.99999997 7.26858547e-07 4.99999997 7.26958547e-07 4.99999997 7.27058547e-07 4.99999997
+ 7.27158547e-07 4.99999997 7.27258547e-07 4.99999997 7.27358547e-07 4.99999997 7.27458547e-07 4.99999997 7.27558547e-07 4.99999997 7.27658547e-07 4.99999997 7.27758547e-07 4.99999997 7.27858547e-07 4.99999997
+ 7.27958547e-07 4.99999997 7.28058547e-07 4.99999997 7.28158547e-07 4.99999997 7.28258547e-07 4.99999997 7.28358547e-07 4.99999997 7.28458547e-07 4.99999997 7.28558547e-07 4.99999997 7.28658547e-07 4.99999997
+ 7.28758547e-07 4.99999997 7.28858547e-07 4.99999997 7.28958547e-07 4.99999997 7.29058547e-07 4.99999997 7.29158547e-07 4.99999997 7.29258547e-07 4.99999997 7.29358547e-07 4.99999997 7.29458547e-07 4.99999997
+ 7.29558547e-07 4.99999997 7.29658547e-07 4.99999997 7.29758547e-07 4.99999997 7.29858547e-07 4.99999997 7.29958547e-07 4.99999997 7.30058547e-07 4.99999997 7.30158547e-07 4.99999997 7.30258547e-07 4.99999997
+ 7.30358547e-07 4.99999997 7.30458547e-07 4.99999997 7.30558547e-07 4.99999997 7.30658547e-07 4.99999997 7.30758547e-07 4.99999997 7.30858547e-07 4.99999997 7.30958547e-07 4.99999997 7.31058547e-07 4.99999997
+ 7.31158547e-07 4.99999997 7.31258547e-07 4.99999997 7.31358547e-07 4.99999997 7.31458547e-07 4.99999997 7.31558547e-07 4.99999997 7.31658547e-07 4.99999997 7.31758547e-07 4.99999997 7.31858547e-07 4.99999997
+ 7.31958547e-07 4.99999997 7.32058547e-07 4.99999997 7.32158547e-07 4.99999997 7.32258547e-07 4.99999997 7.32358547e-07 4.99999997 7.32458547e-07 4.99999997 7.32558547e-07 4.99999997 7.32658547e-07 4.99999997
+ 7.32758547e-07 4.99999997 7.32858547e-07 4.99999997 7.32958547e-07 4.99999997 7.33058547e-07 4.99999997 7.33158547e-07 4.99999997 7.33258547e-07 4.99999997 7.33358547e-07 4.99999997 7.33458547e-07 4.99999997
+ 7.33558547e-07 4.99999997 7.33658547e-07 4.99999997 7.33758547e-07 4.99999997 7.33858547e-07 4.99999997 7.33958547e-07 4.99999997 7.34058547e-07 4.99999997 7.34158547e-07 4.99999997 7.34258547e-07 4.99999997
+ 7.34358547e-07 4.99999997 7.34458547e-07 4.99999997 7.34558547e-07 4.99999997 7.34658547e-07 4.99999997 7.34758547e-07 4.99999997 7.34858547e-07 4.99999997 7.34958547e-07 4.99999997 7.35058547e-07 4.99999997
+ 7.35158547e-07 4.99999997 7.35258547e-07 4.99999997 7.35358547e-07 4.99999997 7.35458547e-07 4.99999997 7.35558547e-07 4.99999997 7.35658547e-07 4.99999997 7.35758547e-07 4.99999997 7.35858547e-07 4.99999997
+ 7.35958547e-07 4.99999997 7.36058547e-07 4.99999997 7.36158547e-07 4.99999997 7.36258547e-07 4.99999997 7.36358547e-07 4.99999997 7.36458547e-07 4.99999997 7.36558547e-07 4.99999997 7.36658547e-07 4.99999997
+ 7.36758547e-07 4.99999997 7.36858547e-07 4.99999997 7.36958547e-07 4.99999997 7.37058547e-07 4.99999997 7.37158547e-07 4.99999997 7.37258547e-07 4.99999997 7.37358547e-07 4.99999997 7.37458547e-07 4.99999997
+ 7.37558547e-07 4.99999997 7.37658547e-07 4.99999997 7.37758547e-07 4.99999997 7.37858547e-07 4.99999997 7.37958547e-07 4.99999997 7.38058547e-07 4.99999997 7.38158547e-07 4.99999997 7.38258547e-07 4.99999997
+ 7.38358547e-07 4.99999997 7.38458547e-07 4.99999997 7.38558547e-07 4.99999997 7.38658547e-07 4.99999997 7.38758547e-07 4.99999997 7.38858547e-07 4.99999997 7.38958547e-07 4.99999997 7.39058547e-07 4.99999997
+ 7.39158547e-07 4.99999997 7.39258547e-07 4.99999997 7.39358547e-07 4.99999997 7.39458547e-07 4.99999997 7.39558547e-07 4.99999997 7.39658547e-07 4.99999997 7.39758547e-07 4.99999997 7.39858547e-07 4.99999997
+ 7.39958547e-07 4.99999997 7.40058547e-07 4.99999997 7.40158547e-07 4.99999997 7.40258547e-07 4.99999997 7.40358547e-07 4.99999997 7.40458547e-07 4.99999997 7.40558547e-07 4.99999997 7.40658547e-07 4.99999997
+ 7.40758547e-07 4.99999997 7.40858547e-07 4.99999997 7.40958547e-07 4.99999997 7.41058547e-07 4.99999997 7.41158547e-07 4.99999997 7.41258547e-07 4.99999997 7.41358547e-07 4.99999997 7.41458547e-07 4.99999997
+ 7.41558547e-07 4.99999997 7.41658547e-07 4.99999997 7.41758547e-07 4.99999997 7.41858547e-07 4.99999997 7.41958547e-07 4.99999997 7.42058547e-07 4.99999997 7.42158547e-07 4.99999997 7.42258547e-07 4.99999997
+ 7.42358547e-07 4.99999997 7.42458547e-07 4.99999997 7.42558547e-07 4.99999997 7.42658547e-07 4.99999997 7.42758547e-07 4.99999997 7.42858547e-07 4.99999997 7.42958547e-07 4.99999997 7.43058547e-07 4.99999997
+ 7.43158547e-07 4.99999997 7.43258547e-07 4.99999997 7.43358547e-07 4.99999997 7.43458547e-07 4.99999997 7.43558547e-07 4.99999997 7.43658547e-07 4.99999997 7.43758547e-07 4.99999997 7.43858547e-07 4.99999997
+ 7.43958547e-07 4.99999997 7.44058547e-07 4.99999997 7.44158547e-07 4.99999997 7.44258547e-07 4.99999997 7.44358547e-07 4.99999997 7.44458547e-07 4.99999997 7.44558547e-07 4.99999997 7.44658547e-07 4.99999997
+ 7.44758547e-07 4.99999997 7.44858547e-07 4.99999997 7.44958547e-07 4.99999997 7.45058547e-07 4.99999997 7.45158547e-07 4.99999997 7.45258547e-07 4.99999997 7.45358547e-07 4.99999997 7.45458547e-07 4.99999997
+ 7.45558547e-07 4.99999997 7.45658547e-07 4.99999997 7.45758547e-07 4.99999997 7.45858547e-07 4.99999997 7.45958547e-07 4.99999997 7.46058547e-07 4.99999997 7.46158547e-07 4.99999997 7.46258547e-07 4.99999997
+ 7.46358547e-07 4.99999997 7.46458547e-07 4.99999997 7.46558547e-07 4.99999997 7.46658547e-07 4.99999997 7.46758547e-07 4.99999997 7.46858547e-07 4.99999997 7.46958547e-07 4.99999997 7.47058547e-07 4.99999997
+ 7.47158547e-07 4.99999997 7.47258547e-07 4.99999997 7.47358547e-07 4.99999997 7.47458547e-07 4.99999997 7.47558547e-07 4.99999997 7.47658547e-07 4.99999997 7.47758547e-07 4.99999997 7.47858547e-07 4.99999997
+ 7.47958547e-07 4.99999997 7.48058547e-07 4.99999997 7.48158547e-07 4.99999997 7.48258547e-07 4.99999997 7.48358547e-07 4.99999997 7.48458547e-07 4.99999997 7.48558547e-07 4.99999997 7.48658547e-07 4.99999997
+ 7.48758547e-07 4.99999997 7.48858547e-07 4.99999997 7.48958547e-07 4.99999997 7.49058547e-07 4.99999997 7.49158547e-07 4.99999997 7.49258547e-07 4.99999997 7.49358547e-07 4.99999997 7.49458547e-07 4.99999997
+ 7.49558547e-07 4.99999997 7.49658547e-07 4.99999997 7.49758547e-07 4.99999997 7.49858547e-07 4.99999997 7.49958547e-07 4.99999997 7.50058547e-07 4.99999997 7.50158547e-07 4.99999997 7.50258547e-07 4.99999997
+ 7.50358547e-07 4.99999997 7.50458547e-07 4.99999997 7.50558547e-07 4.99999997 7.50658547e-07 4.99999997 7.50758547e-07 4.99999997 7.50858547e-07 4.99999997 7.50958547e-07 4.99999997 7.51e-07 4.99999997
+ 7.5101e-07 4.99999997 7.5103e-07 4.99999997 7.5107e-07 4.99999997 7.5115e-07 4.99999997 7.5125e-07 4.99999997 7.5135e-07 4.99999997 7.5145e-07 4.99999997 7.5155e-07 4.99999997
+ 7.5165e-07 4.99999997 7.5175e-07 4.99999997 7.5185e-07 4.99999997 7.51930828e-07 5.00000066 7.52e-07 5.00000151 7.52008608e-07 4.9999927 7.52025825e-07 4.99997482 7.52060258e-07 4.99999285
+ 7.52106188e-07 5.00004461 7.52150118e-07 5.00000795 7.5219811e-07 4.99994547 7.522555e-07 5.00002987 7.52312176e-07 4.9999935 7.52404431e-07 5.0000036 7.52490759e-07 4.99999971 7.52590759e-07 4.99999801
+ 7.52690759e-07 5.00000291 7.52790759e-07 4.99999668 7.52890759e-07 5.00000318 7.52990759e-07 4.99999704 7.53090759e-07 5.00000252 7.53190759e-07 4.99999781 7.53290759e-07 5.00000177 7.53390759e-07 4.9999985
+ 7.53490759e-07 5.00000116 7.53590759e-07 4.99999902 7.53690759e-07 5.00000073 7.53790759e-07 4.99999937 7.53890759e-07 5.00000045 7.53990759e-07 4.99999959 7.54090759e-07 5.00000027 7.54190759e-07 4.99999973
+ 7.54290759e-07 5.00000017 7.54390759e-07 4.99999981 7.54490759e-07 5.0000001 7.54590759e-07 4.99999986 7.54690759e-07 5.00000006 7.54790759e-07 4.99999989 7.54890759e-07 5.00000004 7.54990759e-07 4.99999991
+ 7.55090759e-07 5.00000002 7.55190759e-07 4.99999992 7.55290759e-07 5.00000002 7.55390759e-07 4.99999993 7.55490759e-07 5.00000001 7.55590759e-07 4.99999994 7.55690759e-07 5.0 7.55790759e-07 4.99999994
+ 7.55890759e-07 5.0 7.55990759e-07 4.99999994 7.56090759e-07 5.0 7.56190759e-07 4.99999995 7.56290759e-07 5.0 7.56390759e-07 4.99999995 7.56490759e-07 4.99999999 7.56590759e-07 4.99999995
+ 7.56690759e-07 4.99999999 7.56790759e-07 4.99999995 7.56890759e-07 4.99999999 7.56990759e-07 4.99999995 7.57090759e-07 4.99999999 7.57190759e-07 4.99999996 7.57290759e-07 4.99999999 7.57390759e-07 4.99999996
+ 7.57490759e-07 4.99999999 7.57590759e-07 4.99999996 7.57690759e-07 4.99999998 7.57790759e-07 4.99999996 7.57890759e-07 4.99999998 7.57990759e-07 4.99999996 7.58090759e-07 4.99999998 7.58190759e-07 4.99999996
+ 7.58290759e-07 4.99999998 7.58390759e-07 4.99999996 7.58490759e-07 4.99999998 7.58590759e-07 4.99999997 7.58690759e-07 4.99999998 7.58790759e-07 4.99999997 7.58890759e-07 4.99999998 7.58990759e-07 4.99999997
+ 7.59090759e-07 4.99999998 7.59190759e-07 4.99999997 7.59290759e-07 4.99999998 7.59390759e-07 4.99999997 7.59490759e-07 4.99999998 7.59590759e-07 4.99999997 7.59690759e-07 4.99999998 7.59790759e-07 4.99999997
+ 7.59890759e-07 4.99999998 7.59990759e-07 4.99999997 7.60090759e-07 4.99999997 7.60190759e-07 4.99999997 7.60290759e-07 4.99999997 7.60390759e-07 4.99999997 7.60490759e-07 4.99999997 7.60590759e-07 4.99999997
+ 7.60690759e-07 4.99999997 7.60790759e-07 4.99999997 7.60890759e-07 4.99999997 7.60990759e-07 4.99999997 7.61090759e-07 4.99999997 7.61190759e-07 4.99999997 7.61290759e-07 4.99999997 7.61390759e-07 4.99999997
+ 7.61490759e-07 4.99999997 7.61590759e-07 4.99999997 7.61690759e-07 4.99999997 7.61790759e-07 4.99999997 7.61890759e-07 4.99999997 7.61990759e-07 4.99999997 7.62090759e-07 4.99999997 7.62190759e-07 4.99999997
+ 7.62290759e-07 4.99999997 7.62390759e-07 4.99999997 7.62490759e-07 4.99999997 7.62590759e-07 4.99999997 7.62690759e-07 4.99999997 7.62790759e-07 4.99999997 7.62890759e-07 4.99999997 7.62990759e-07 4.99999997
+ 7.63090759e-07 4.99999997 7.63190759e-07 4.99999997 7.63290759e-07 4.99999997 7.63390759e-07 4.99999997 7.63490759e-07 4.99999997 7.63590759e-07 4.99999997 7.63690759e-07 4.99999997 7.63790759e-07 4.99999997
+ 7.63890759e-07 4.99999997 7.63990759e-07 4.99999997 7.64090759e-07 4.99999997 7.64190759e-07 4.99999997 7.64290759e-07 4.99999997 7.64390759e-07 4.99999997 7.64490759e-07 4.99999997 7.64590759e-07 4.99999997
+ 7.64690759e-07 4.99999997 7.64790759e-07 4.99999997 7.64890759e-07 4.99999997 7.64990759e-07 4.99999997 7.65090759e-07 4.99999997 7.65190759e-07 4.99999997 7.65290759e-07 4.99999997 7.65390759e-07 4.99999997
+ 7.65490759e-07 4.99999997 7.65590759e-07 4.99999997 7.65690759e-07 4.99999997 7.65790759e-07 4.99999997 7.65890759e-07 4.99999997 7.65990759e-07 4.99999997 7.66090759e-07 4.99999997 7.66190759e-07 4.99999997
+ 7.66290759e-07 4.99999997 7.66390759e-07 4.99999997 7.66490759e-07 4.99999997 7.66590759e-07 4.99999997 7.66690759e-07 4.99999997 7.66790759e-07 4.99999997 7.66890759e-07 4.99999997 7.66990759e-07 4.99999997
+ 7.67090759e-07 4.99999997 7.67190759e-07 4.99999997 7.67290759e-07 4.99999997 7.67390759e-07 4.99999997 7.67490759e-07 4.99999997 7.67590759e-07 4.99999997 7.67690759e-07 4.99999997 7.67790759e-07 4.99999997
+ 7.67890759e-07 4.99999997 7.67990759e-07 4.99999997 7.68090759e-07 4.99999997 7.68190759e-07 4.99999997 7.68290759e-07 4.99999997 7.68390759e-07 4.99999997 7.68490759e-07 4.99999997 7.68590759e-07 4.99999997
+ 7.68690759e-07 4.99999997 7.68790759e-07 4.99999997 7.68890759e-07 4.99999997 7.68990759e-07 4.99999997 7.69090759e-07 4.99999997 7.69190759e-07 4.99999997 7.69290759e-07 4.99999997 7.69390759e-07 4.99999997
+ 7.69490759e-07 4.99999997 7.69590759e-07 4.99999997 7.69690759e-07 4.99999997 7.69790759e-07 4.99999997 7.69890759e-07 4.99999997 7.69990759e-07 4.99999997 7.70090759e-07 4.99999997 7.70190759e-07 4.99999997
+ 7.70290759e-07 4.99999997 7.70390759e-07 4.99999997 7.70490759e-07 4.99999997 7.70590759e-07 4.99999997 7.70690759e-07 4.99999997 7.70790759e-07 4.99999997 7.70890759e-07 4.99999997 7.70990759e-07 4.99999997
+ 7.71090759e-07 4.99999997 7.71190759e-07 4.99999997 7.71290759e-07 4.99999997 7.71390759e-07 4.99999997 7.71490759e-07 4.99999997 7.71590759e-07 4.99999997 7.71690759e-07 4.99999997 7.71790759e-07 4.99999997
+ 7.71890759e-07 4.99999997 7.71990759e-07 4.99999997 7.72090759e-07 4.99999997 7.72190759e-07 4.99999997 7.72290759e-07 4.99999997 7.72390759e-07 4.99999997 7.72490759e-07 4.99999997 7.72590759e-07 4.99999997
+ 7.72690759e-07 4.99999997 7.72790759e-07 4.99999997 7.72890759e-07 4.99999997 7.72990759e-07 4.99999997 7.73090759e-07 4.99999997 7.73190759e-07 4.99999997 7.73290759e-07 4.99999997 7.73390759e-07 4.99999997
+ 7.73490759e-07 4.99999997 7.73590759e-07 4.99999997 7.73690759e-07 4.99999997 7.73790759e-07 4.99999997 7.73890759e-07 4.99999997 7.73990759e-07 4.99999997 7.74090759e-07 4.99999997 7.74190759e-07 4.99999997
+ 7.74290759e-07 4.99999997 7.74390759e-07 4.99999997 7.74490759e-07 4.99999997 7.74590759e-07 4.99999997 7.74690759e-07 4.99999997 7.74790759e-07 4.99999997 7.74890759e-07 4.99999997 7.74990759e-07 4.99999997
+ 7.75090759e-07 4.99999997 7.75190759e-07 4.99999997 7.75290759e-07 4.99999997 7.75390759e-07 4.99999997 7.75490759e-07 4.99999997 7.75590759e-07 4.99999997 7.75690759e-07 4.99999997 7.75790759e-07 4.99999997
+ 7.75890759e-07 4.99999997 7.75990759e-07 4.99999997 7.76090759e-07 4.99999997 7.76190759e-07 4.99999997 7.76290759e-07 4.99999997 7.76390759e-07 4.99999997 7.76490759e-07 4.99999997 7.76590759e-07 4.99999997
+ 7.76690759e-07 4.99999997 7.76790759e-07 4.99999997 7.76890759e-07 4.99999997 7.76990759e-07 4.99999997 7.77090759e-07 4.99999997 7.77190759e-07 4.99999997 7.77290759e-07 4.99999997 7.77390759e-07 4.99999997
+ 7.77490759e-07 4.99999997 7.77590759e-07 4.99999997 7.77690759e-07 4.99999997 7.77790759e-07 4.99999997 7.77890759e-07 4.99999997 7.77990759e-07 4.99999997 7.78090759e-07 4.99999997 7.78190759e-07 4.99999997
+ 7.78290759e-07 4.99999997 7.78390759e-07 4.99999997 7.78490759e-07 4.99999997 7.78590759e-07 4.99999997 7.78690759e-07 4.99999997 7.78790759e-07 4.99999997 7.78890759e-07 4.99999997 7.78990759e-07 4.99999997
+ 7.79090759e-07 4.99999997 7.79190759e-07 4.99999997 7.79290759e-07 4.99999997 7.79390759e-07 4.99999997 7.79490759e-07 4.99999997 7.79590759e-07 4.99999997 7.79690759e-07 4.99999997 7.79790759e-07 4.99999997
+ 7.79890759e-07 4.99999997 7.79990759e-07 4.99999997 7.80090759e-07 4.99999997 7.80190759e-07 4.99999997 7.80290759e-07 4.99999997 7.80390759e-07 4.99999997 7.80490759e-07 4.99999997 7.80590759e-07 4.99999997
+ 7.80690759e-07 4.99999997 7.80790759e-07 4.99999997 7.80890759e-07 4.99999997 7.80990759e-07 4.99999997 7.81090759e-07 4.99999997 7.81190759e-07 4.99999997 7.81290759e-07 4.99999997 7.81390759e-07 4.99999997
+ 7.81490759e-07 4.99999997 7.81590759e-07 4.99999997 7.81690759e-07 4.99999997 7.81790759e-07 4.99999997 7.81890759e-07 4.99999997 7.81990759e-07 4.99999997 7.82090759e-07 4.99999997 7.82190759e-07 4.99999997
+ 7.82290759e-07 4.99999997 7.82390759e-07 4.99999997 7.82490759e-07 4.99999997 7.82590759e-07 4.99999997 7.82690759e-07 4.99999997 7.82790759e-07 4.99999997 7.82890759e-07 4.99999997 7.82990759e-07 4.99999997
+ 7.83090759e-07 4.99999997 7.83190759e-07 4.99999997 7.83290759e-07 4.99999997 7.83390759e-07 4.99999997 7.83490759e-07 4.99999997 7.83590759e-07 4.99999997 7.83690759e-07 4.99999997 7.83790759e-07 4.99999997
+ 7.83890759e-07 4.99999997 7.83990759e-07 4.99999997 7.84090759e-07 4.99999997 7.84190759e-07 4.99999997 7.84290759e-07 4.99999997 7.84390759e-07 4.99999997 7.84490759e-07 4.99999997 7.84590759e-07 4.99999997
+ 7.84690759e-07 4.99999997 7.84790759e-07 4.99999997 7.84890759e-07 4.99999997 7.84990759e-07 4.99999997 7.85090759e-07 4.99999997 7.85190759e-07 4.99999997 7.85290759e-07 4.99999997 7.85390759e-07 4.99999997
+ 7.85490759e-07 4.99999997 7.85590759e-07 4.99999997 7.85690759e-07 4.99999997 7.85790759e-07 4.99999997 7.85890759e-07 4.99999997 7.85990759e-07 4.99999997 7.86090759e-07 4.99999997 7.86190759e-07 4.99999997
+ 7.86290759e-07 4.99999997 7.86390759e-07 4.99999997 7.86490759e-07 4.99999997 7.86590759e-07 4.99999997 7.86690759e-07 4.99999997 7.86790759e-07 4.99999997 7.86890759e-07 4.99999997 7.86990759e-07 4.99999997
+ 7.87090759e-07 4.99999997 7.87190759e-07 4.99999997 7.87290759e-07 4.99999997 7.87390759e-07 4.99999997 7.87490759e-07 4.99999997 7.87590759e-07 4.99999997 7.87690759e-07 4.99999997 7.87790759e-07 4.99999997
+ 7.87890759e-07 4.99999997 7.87990759e-07 4.99999997 7.88090759e-07 4.99999997 7.88190759e-07 4.99999997 7.88290759e-07 4.99999997 7.88390759e-07 4.99999997 7.88490759e-07 4.99999997 7.88590759e-07 4.99999997
+ 7.88690759e-07 4.99999997 7.88790759e-07 4.99999997 7.88890759e-07 4.99999997 7.88990759e-07 4.99999997 7.89090759e-07 4.99999997 7.89190759e-07 4.99999997 7.89290759e-07 4.99999997 7.89390759e-07 4.99999997
+ 7.89490759e-07 4.99999997 7.89590759e-07 4.99999997 7.89690759e-07 4.99999997 7.89790759e-07 4.99999997 7.89890759e-07 4.99999997 7.89990759e-07 4.99999997 7.90090759e-07 4.99999997 7.90190759e-07 4.99999997
+ 7.90290759e-07 4.99999997 7.90390759e-07 4.99999997 7.90490759e-07 4.99999997 7.90590759e-07 4.99999997 7.90690759e-07 4.99999997 7.90790759e-07 4.99999997 7.90890759e-07 4.99999997 7.90990759e-07 4.99999997
+ 7.91090759e-07 4.99999997 7.91190759e-07 4.99999997 7.91290759e-07 4.99999997 7.91390759e-07 4.99999997 7.91490759e-07 4.99999997 7.91590759e-07 4.99999997 7.91690759e-07 4.99999997 7.91790759e-07 4.99999997
+ 7.91890759e-07 4.99999997 7.91990759e-07 4.99999997 7.92090759e-07 4.99999997 7.92190759e-07 4.99999997 7.92290759e-07 4.99999997 7.92390759e-07 4.99999997 7.92490759e-07 4.99999997 7.92590759e-07 4.99999997
+ 7.92690759e-07 4.99999997 7.92790759e-07 4.99999997 7.92890759e-07 4.99999997 7.92990759e-07 4.99999997 7.93090759e-07 4.99999997 7.93190759e-07 4.99999997 7.93290759e-07 4.99999997 7.93390759e-07 4.99999997
+ 7.93490759e-07 4.99999997 7.93590759e-07 4.99999997 7.93690759e-07 4.99999997 7.93790759e-07 4.99999997 7.93890759e-07 4.99999997 7.93990759e-07 4.99999997 7.94090759e-07 4.99999997 7.94190759e-07 4.99999997
+ 7.94290759e-07 4.99999997 7.94390759e-07 4.99999997 7.94490759e-07 4.99999997 7.94590759e-07 4.99999997 7.94690759e-07 4.99999997 7.94790759e-07 4.99999997 7.94890759e-07 4.99999997 7.94990759e-07 4.99999997
+ 7.95090759e-07 4.99999997 7.95190759e-07 4.99999997 7.95290759e-07 4.99999997 7.95390759e-07 4.99999997 7.95490759e-07 4.99999997 7.95590759e-07 4.99999997 7.95690759e-07 4.99999997 7.95790759e-07 4.99999997
+ 7.95890759e-07 4.99999997 7.95990759e-07 4.99999997 7.96090759e-07 4.99999997 7.96190759e-07 4.99999997 7.96290759e-07 4.99999997 7.96390759e-07 4.99999997 7.96490759e-07 4.99999997 7.96590759e-07 4.99999997
+ 7.96690759e-07 4.99999997 7.96790759e-07 4.99999997 7.96890759e-07 4.99999997 7.96990759e-07 4.99999997 7.97090759e-07 4.99999997 7.97190759e-07 4.99999997 7.97290759e-07 4.99999997 7.97390759e-07 4.99999997
+ 7.97490759e-07 4.99999997 7.97590759e-07 4.99999997 7.97690759e-07 4.99999997 7.97790759e-07 4.99999997 7.97890759e-07 4.99999997 7.97990759e-07 4.99999997 7.98090759e-07 4.99999997 7.98190759e-07 4.99999997
+ 7.98290759e-07 4.99999997 7.98390759e-07 4.99999997 7.98490759e-07 4.99999997 7.98590759e-07 4.99999997 7.98690759e-07 4.99999997 7.98790759e-07 4.99999997 7.98890759e-07 4.99999997 7.98990759e-07 4.99999997
+ 7.99090759e-07 4.99999997 7.99190759e-07 4.99999997 7.99290759e-07 4.99999997 7.99390759e-07 4.99999997 7.99490759e-07 4.99999997 7.99590759e-07 4.99999997 7.99690759e-07 4.99999997 7.99790759e-07 4.99999997
+ 7.99890759e-07 4.99999997 7.99990759e-07 4.99999997 8e-07 4.99999997 8.0001e-07 4.99999997 8.0003e-07 4.99999997 8.0007e-07 4.99999997 8.0015e-07 4.99999997 8.0025e-07 4.99999997
+ 8.0035e-07 4.99999997 8.0045e-07 4.99999997 8.0055e-07 4.99999997 8.0065e-07 4.99999997 8.0075e-07 5.00000001 8.0085e-07 4.99999717 8.00931913e-07 5.00000328 8.01e-07 5.00008601
+ 8.01008477e-07 5.00011635 8.01025432e-07 5.00022698 8.01059342e-07 4.99960029 8.01090545e-07 4.99796703 8.01143412e-07 4.99703072 8.01199108e-07 5.02828621 8.01266691e-07 4.9918975 8.01329415e-07 3.49023986
+ 8.01394829e-07 0.154819829 8.01464618e-07 -0.00376126514 8.01533535e-07 0.0257937047 8.01610366e-07 -0.0174819665 8.01709241e-07 0.0166256226 8.01809241e-07 -0.0151036136 8.01909241e-07 0.0138168911 8.02009241e-07 -0.0125784687
+ 8.02109241e-07 0.011505171 8.02209241e-07 -0.010481817 8.02309241e-07 0.00958739706 8.02409241e-07 -0.00873958877 8.02509241e-07 0.00799375037 8.02609241e-07 -0.00729006223 8.02709241e-07 0.00666768862 8.02809241e-07 -0.00608276976
+ 8.02909241e-07 0.00556317247 8.03009241e-07 -0.00507645127 8.03109241e-07 0.00464253506 8.03209241e-07 -0.00423720493 8.03309241e-07 0.00387478758 8.03409241e-07 -0.00353704076 8.03509241e-07 0.00323432261 8.03609241e-07 -0.00295276769
+ 8.03709241e-07 0.00269991248 8.03809241e-07 -0.00246512287 8.03909241e-07 0.00225392144 8.04009241e-07 -0.00205807943 8.04109241e-07 0.00188167602 8.04209241e-07 -0.00171828798 8.04309241e-07 0.00157095524 8.04409241e-07 -0.00143462118
+ 8.04509241e-07 0.00131157363 8.04609241e-07 -0.00119779915 8.04709241e-07 0.00109503818 8.04809241e-07 -0.00100008016 8.04909241e-07 0.000914264687 8.05009241e-07 -0.000835004145 8.05109241e-07 0.000763342619 8.05209241e-07 -0.00069717962
+ 8.05309241e-07 0.000637339801 8.05409241e-07 -0.000582106412 8.05509241e-07 0.000532139928 8.05609241e-07 -0.000486027981 8.05709241e-07 0.000444307246 8.05809241e-07 -0.000405808347 8.05909241e-07 0.000370973849 8.06009241e-07 -0.000338829481
+ 8.06109241e-07 0.000309745686 8.06209241e-07 -0.000282905677 8.06309241e-07 0.000258624171 8.06409241e-07 -0.000236212099 8.06509241e-07 0.000215940793 8.06609241e-07 -0.000197225188 8.06709241e-07 0.000180302581 8.06809241e-07 -0.000164672908
+ 8.06909241e-07 0.000151581252 8.07009241e-07 -0.000137330071 8.07109241e-07 0.000125617353 8.07209241e-07 -0.000114721651 8.07309241e-07 0.000104886816 8.07409241e-07 -9.57863029e-05 8.07509241e-07 8.75782273e-05 8.07609241e-07 -7.99758898e-05
+ 8.07709241e-07 7.31262283e-05 8.07809241e-07 -6.67747637e-05 8.07909241e-07 6.14617377e-05 8.08009241e-07 -5.56877955e-05 8.08109241e-07 5.12854283e-05 8.08209241e-07 -4.64651204e-05 8.08309241e-07 4.27945085e-05 8.08409241e-07 -3.85326677e-05
+ 8.08509241e-07 3.57459199e-05 8.08609241e-07 -3.21645777e-05 8.08709241e-07 2.98427245e-05 8.08809241e-07 -2.68487335e-05 8.08909241e-07 2.49148683e-05 8.09009241e-07 -2.24112808e-05 8.09109241e-07 2.08011545e-05 8.09209241e-07 -1.87070504e-05
+ 8.09309241e-07 1.73671183e-05 8.09409241e-07 -1.56148482e-05 8.09509241e-07 1.45003217e-05 8.09609241e-07 -1.30334472e-05 8.09709241e-07 1.2107067e-05 8.09809241e-07 -1.08784781e-05 8.09909241e-07 1.01091346e-05 8.10009241e-07 -9.07948871e-06
+ 8.10109241e-07 8.44121874e-06 8.10209241e-07 -7.57766587e-06 8.10309241e-07 7.04880191e-06 8.10409241e-07 -6.3239152e-06 8.10509241e-07 5.8863742e-06 8.10609241e-07 -5.27725522e-06 8.10709241e-07 4.91594507e-06 8.10809241e-07 -4.40347637e-06
+ 8.10909241e-07 4.10580046e-06 8.11009241e-07 -3.67402123e-06 8.11109241e-07 3.42946531e-06 8.11209241e-07 -3.06505021e-06 8.11309241e-07 2.8648379e-06 8.11409241e-07 -2.55666197e-06 8.11509241e-07 2.39346732e-06 8.11609241e-07 -2.13224273e-06
+ 8.11709241e-07 1.99995037e-06 8.11809241e-07 -1.77792302e-06 8.11909241e-07 1.67142791e-06 8.12009241e-07 -1.48212383e-06 8.12109241e-07 1.39716414e-06 8.12209241e-07 -1.23517925e-06 8.12309241e-07 1.16819841e-06 8.12409241e-07 -1.0290213e-06
+ 8.12509241e-07 9.77049652e-07 8.12609241e-07 -8.56913387e-07 8.12709241e-07 8.17471684e-07 8.12809241e-07 -7.13231541e-07 8.12909241e-07 6.84250153e-07 8.13009241e-07 -5.93280523e-07 8.13109241e-07 5.73031515e-07 8.13209241e-07 -4.93140772e-07
+ 8.13309241e-07 4.80181928e-07 8.13409241e-07 -4.09540301e-07 8.13509241e-07 4.02667501e-07 8.13609241e-07 -3.39747397e-07 8.13709241e-07 3.37955414e-07 8.13809241e-07 -2.81481545e-07 8.13909241e-07 2.83931202e-07 8.14009241e-07 -2.32838909e-07
+ 8.14109241e-07 2.38829636e-07 8.14209241e-07 -1.92230101e-07 8.14309241e-07 2.01177043e-07 8.14409241e-07 -1.58328245e-07 8.14509241e-07 1.69743148e-07 8.14609241e-07 -1.30025615e-07 8.14709241e-07 1.43500865e-07 8.14809241e-07 -1.06397437e-07
+ 8.14909241e-07 1.21592743e-07 8.15009241e-07 -8.66716736e-08 8.15109241e-07 1.03302951e-07 8.15209241e-07 -7.02059618e-08 8.15309241e-07 8.80380011e-08 8.15409241e-07 -5.64647247e-08 8.15509241e-07 7.53001782e-08 8.15609241e-07 -4.49983217e-08
+ 8.15709241e-07 6.46710726e-08 8.15809241e-07 -3.54301521e-08 8.15909241e-07 5.5801589e-08 8.16009241e-07 -2.74459685e-08 8.16109241e-07 4.84004266e-08 8.16209241e-07 -2.07835451e-08 8.16309241e-07 4.22245088e-08 8.16409241e-07 -1.52102918e-08
+ 8.16509241e-07 3.70584681e-08 8.16609241e-07 -1.05742361e-08 8.16709241e-07 3.27607126e-08 8.16809241e-07 -6.70534886e-09 8.16909241e-07 2.91743369e-08 8.17009241e-07 -3.47686099e-09 8.17109241e-07 2.61816047e-08 8.17209241e-07 -7.82778814e-10
+ 8.17309241e-07 2.36842577e-08 8.17409241e-07 1.46535367e-09 8.17509241e-07 2.16193711e-08 8.17609241e-07 3.32511205e-09 8.17709241e-07 1.99196331e-08 8.17809241e-07 4.85641755e-09 8.17909241e-07 1.85200861e-08 8.18009241e-07 6.11728254e-09
+ 8.18109241e-07 1.73677094e-08 8.18209241e-07 7.15547221e-09 8.18309241e-07 1.64188494e-08 8.18409241e-07 8.01030936e-09 8.18509241e-07 1.56375695e-08 8.18609241e-07 8.7141723e-09 8.18709241e-07 1.48973149e-08 8.18809241e-07 9.27994537e-09
+ 8.18909241e-07 1.43787412e-08 8.19009241e-07 9.75062581e-09 8.19109241e-07 1.39514974e-08 8.19209241e-07 1.01384438e-08 8.19309241e-07 1.35994825e-08 8.19409241e-07 1.04579696e-08 8.19509241e-07 1.33094584e-08 8.19609241e-07 1.07212254e-08
+ 8.19709241e-07 1.30705116e-08 8.19809241e-07 1.09381179e-08 8.19909241e-07 1.28736473e-08 8.20009241e-07 1.11168121e-08 8.20109241e-07 1.27114549e-08 8.20209241e-07 1.12640354e-08 8.20309241e-07 1.25778278e-08 8.20409241e-07 1.13853303e-08
+ 8.20509241e-07 1.24677355e-08 8.20609241e-07 1.14852626e-08 8.20709241e-07 1.23770332e-08 8.20809241e-07 1.15675949e-08 8.20909241e-07 1.23023062e-08 8.21009241e-07 1.16354266e-08 8.21109241e-07 1.22407405e-08 8.21209241e-07 1.16913121e-08
+ 8.21309241e-07 1.21900182e-08 8.21409241e-07 1.17373551e-08 8.21509241e-07 1.21482295e-08 8.21609241e-07 1.17752891e-08 8.21709241e-07 1.2113801e-08 8.21809241e-07 1.18065423e-08 8.21909241e-07 1.20854362e-08 8.22009241e-07 1.18322916e-08
+ 8.22109241e-07 1.20620668e-08 8.22209241e-07 1.18535064e-08 8.22309241e-07 1.20428138e-08 8.22409241e-07 1.18709849e-08 8.22509241e-07 1.20269515e-08 8.22609241e-07 1.18853851e-08 8.22709241e-07 1.20138834e-08 8.22809241e-07 1.18972497e-08
+ 8.22909241e-07 1.20031166e-08 8.23009241e-07 1.19070248e-08 8.23109241e-07 1.19942465e-08 8.23209241e-07 1.19150786e-08 8.23309241e-07 1.19869385e-08 8.23409241e-07 1.19217138e-08 8.23509241e-07 1.19809181e-08 8.23609241e-07 1.1927181e-08
+ 8.23709241e-07 1.19759581e-08 8.23809241e-07 1.19316854e-08 8.23909241e-07 1.19718719e-08 8.24009241e-07 1.19353963e-08 8.24109241e-07 1.19685051e-08 8.24209241e-07 1.19384543e-08 8.24309241e-07 1.19657318e-08 8.24409241e-07 1.19409732e-08
+ 8.24509241e-07 1.1963447e-08 8.24609241e-07 1.19430492e-08 8.24709241e-07 1.19615647e-08 8.24809241e-07 1.19447596e-08 8.24909241e-07 1.19600138e-08 8.25009241e-07 1.19461686e-08 8.25109241e-07 1.19587365e-08 8.25209241e-07 1.19473297e-08
+ 8.25309241e-07 1.19576843e-08 8.25409241e-07 1.19482865e-08 8.25509241e-07 1.19568178e-08 8.25609241e-07 1.19490745e-08 8.25709241e-07 1.19561035e-08 8.25809241e-07 1.19497241e-08 8.25909241e-07 1.19555155e-08 8.26009241e-07 1.19502596e-08
+ 8.26109241e-07 1.19550309e-08 8.26209241e-07 1.19507006e-08 8.26309241e-07 1.19546319e-08 8.26409241e-07 1.1951064e-08 8.26509241e-07 1.19543034e-08 8.26609241e-07 1.19513638e-08 8.26709241e-07 1.19540326e-08 8.26809241e-07 1.19516104e-08
+ 8.26909241e-07 1.19538095e-08 8.27009241e-07 1.19518142e-08 8.27109241e-07 1.19536262e-08 8.27209241e-07 1.19519823e-08 8.27309241e-07 1.19534746e-08 8.27409241e-07 1.19521203e-08 8.27509241e-07 1.19533501e-08 8.27609241e-07 1.19522346e-08
+ 8.27709241e-07 1.19532476e-08 8.27809241e-07 1.19523288e-08 8.27909241e-07 1.19531633e-08 8.28009241e-07 1.19524061e-08 8.28109241e-07 1.19530941e-08 8.28209241e-07 1.19524703e-08 8.28309241e-07 1.19530367e-08 8.28409241e-07 1.1952523e-08
+ 8.28509241e-07 1.19529898e-08 8.28609241e-07 1.19525667e-08 8.28709241e-07 1.19529514e-08 8.28809241e-07 1.19526025e-08 8.28909241e-07 1.19529196e-08 8.29009241e-07 1.19526322e-08 8.29109241e-07 1.19528936e-08 8.29209241e-07 1.1952657e-08
+ 8.29309241e-07 1.1952872e-08 8.29409241e-07 1.19526772e-08 8.29509241e-07 1.19528542e-08 8.29609241e-07 1.1952694e-08 8.29709241e-07 1.19528397e-08 8.29809241e-07 1.19527078e-08 8.29909241e-07 1.19528279e-08 8.30009241e-07 1.19527193e-08
+ 8.30109241e-07 1.19528183e-08 8.30209241e-07 1.19527286e-08 8.30309241e-07 1.19528107e-08 8.30409241e-07 1.19527364e-08 8.30509241e-07 1.19528039e-08 8.30609241e-07 1.19527432e-08 8.30709241e-07 1.19527988e-08 8.30809241e-07 1.19527485e-08
+ 8.30909241e-07 1.19527944e-08 8.31009241e-07 1.19527531e-08 8.31109241e-07 1.19527911e-08 8.31209241e-07 1.19527569e-08 8.31309241e-07 1.19527882e-08 8.31409241e-07 1.19527599e-08 8.31509241e-07 1.19527857e-08 8.31609241e-07 1.1952763e-08
+ 8.31709241e-07 1.1952784e-08 8.31809241e-07 1.19527652e-08 8.31909241e-07 1.19527823e-08 8.32009241e-07 1.19527672e-08 8.32109241e-07 1.19527811e-08 8.32209241e-07 1.19527687e-08 8.32309241e-07 1.19527801e-08 8.32409241e-07 1.19527702e-08
+ 8.32509241e-07 1.19527795e-08 8.32609241e-07 1.1952771e-08 8.32709241e-07 1.19527792e-08 8.32809241e-07 1.19527722e-08 8.32909241e-07 1.19527787e-08 8.33009241e-07 1.19527729e-08 8.33109241e-07 1.19527784e-08 8.33209241e-07 1.19527736e-08
+ 8.33309241e-07 1.19527783e-08 8.33409241e-07 1.19527742e-08 8.33509241e-07 1.19527784e-08 8.33609241e-07 1.19527749e-08 8.33709241e-07 1.19527782e-08 8.33809241e-07 1.19527753e-08 8.33909241e-07 1.1952778e-08 8.34009241e-07 1.19527759e-08
+ 8.34109241e-07 1.19527779e-08 8.34209241e-07 1.19527763e-08 8.34309241e-07 1.1952778e-08 8.34409241e-07 1.19527768e-08 8.34509241e-07 1.19527783e-08 8.34609241e-07 1.1952777e-08 8.34709241e-07 1.19527783e-08 8.34809241e-07 1.19527775e-08
+ 8.34909241e-07 1.19527785e-08 8.35009241e-07 1.19527773e-08 8.35109241e-07 1.19527785e-08 8.35209241e-07 1.19527778e-08 8.35309241e-07 1.19527787e-08 8.35409241e-07 1.1952778e-08 8.35509241e-07 1.1952779e-08 8.35609241e-07 1.19527782e-08
+ 8.35709241e-07 1.19527792e-08 8.35809241e-07 1.19527784e-08 8.35909241e-07 1.19527791e-08 8.36009241e-07 1.19527785e-08 8.36109241e-07 1.19527793e-08 8.36209241e-07 1.19527785e-08 8.36309241e-07 1.19527795e-08 8.36409241e-07 1.19527789e-08
+ 8.36509241e-07 1.19527797e-08 8.36609241e-07 1.1952779e-08 8.36709241e-07 1.19527799e-08 8.36809241e-07 1.19527794e-08 8.36909241e-07 1.19527799e-08 8.37009241e-07 1.19527796e-08 8.37109241e-07 1.195278e-08 8.37209241e-07 1.19527798e-08
+ 8.37309241e-07 1.19527802e-08 8.37409241e-07 1.195278e-08 8.37509241e-07 1.195278e-08 8.37609241e-07 1.195278e-08 8.37709241e-07 1.19527803e-08 8.37809241e-07 1.19527802e-08 8.37909241e-07 1.19527803e-08 8.38009241e-07 1.19527806e-08
+ 8.38109241e-07 1.19527808e-08 8.38209241e-07 1.19527805e-08 8.38309241e-07 1.19527807e-08 8.38409241e-07 1.19527807e-08 8.38509241e-07 1.19527809e-08 8.38609241e-07 1.19527809e-08 8.38709241e-07 1.19527811e-08 8.38809241e-07 1.19527807e-08
+ 8.38909241e-07 1.19527811e-08 8.39009241e-07 1.19527809e-08 8.39109241e-07 1.19527815e-08 8.39209241e-07 1.19527807e-08 8.39309241e-07 1.19527816e-08 8.39409241e-07 1.19527811e-08 8.39509241e-07 1.19527817e-08 8.39609241e-07 1.19527811e-08
+ 8.39709241e-07 1.19527816e-08 8.39809241e-07 1.19527817e-08 8.39909241e-07 1.19527818e-08 8.40009241e-07 1.19527817e-08 8.40109241e-07 1.19527821e-08 8.40209241e-07 1.19527815e-08 8.40309241e-07 1.19527822e-08 8.40409241e-07 1.19527814e-08
+ 8.40509241e-07 1.19527823e-08 8.40609241e-07 1.19527817e-08 8.40709241e-07 1.19527823e-08 8.40809241e-07 1.19527818e-08 8.40909241e-07 1.19527824e-08 8.41009241e-07 1.19527822e-08 8.41109241e-07 1.19527821e-08 8.41209241e-07 1.19527824e-08
+ 8.41309241e-07 1.19527824e-08 8.41409241e-07 1.19527823e-08 8.41509241e-07 1.19527822e-08 8.41609241e-07 1.19527826e-08 8.41709241e-07 1.19527826e-08 8.41809241e-07 1.19527827e-08 8.41909241e-07 1.19527827e-08 8.42009241e-07 1.19527824e-08
+ 8.42109241e-07 1.19527828e-08 8.42209241e-07 1.19527825e-08 8.42309241e-07 1.19527829e-08 8.42409241e-07 1.19527825e-08 8.42509241e-07 1.19527829e-08 8.42609241e-07 1.19527829e-08 8.42709241e-07 1.19527831e-08 8.42809241e-07 1.19527829e-08
+ 8.42909241e-07 1.19527829e-08 8.43009241e-07 1.1952783e-08 8.43109241e-07 1.19527832e-08 8.43209241e-07 1.1952783e-08 8.43309241e-07 1.1952783e-08 8.43409241e-07 1.1952783e-08 8.43509241e-07 1.19527832e-08 8.43609241e-07 1.19527833e-08
+ 8.43709241e-07 1.19527835e-08 8.43809241e-07 1.19527833e-08 8.43909241e-07 1.19527834e-08 8.44009241e-07 1.19527832e-08 8.44109241e-07 1.19527834e-08 8.44209241e-07 1.19527834e-08 8.44309241e-07 1.19527839e-08 8.44409241e-07 1.19527835e-08
+ 8.44509241e-07 1.19527835e-08 8.44609241e-07 1.19527837e-08 8.44709241e-07 1.19527838e-08 8.44809241e-07 1.19527836e-08 8.44909241e-07 1.19527836e-08 8.45009241e-07 1.19527838e-08 8.45109241e-07 1.19527839e-08 8.45209241e-07 1.19527837e-08
+ 8.45309241e-07 1.19527838e-08 8.45409241e-07 1.1952784e-08 8.45509241e-07 1.1952784e-08 8.45609241e-07 1.19527838e-08 8.45709241e-07 1.1952784e-08 8.45809241e-07 1.1952784e-08 8.45909241e-07 1.19527842e-08 8.46009241e-07 1.1952784e-08
+ 8.46109241e-07 1.19527839e-08 8.46209241e-07 1.19527842e-08 8.46309241e-07 1.19527844e-08 8.46409241e-07 1.19527841e-08 8.46509241e-07 1.19527843e-08 8.46609241e-07 1.19527846e-08 8.46709241e-07 1.19527842e-08 8.46809241e-07 1.19527845e-08
+ 8.46909241e-07 1.19527843e-08 8.47009241e-07 1.19527844e-08 8.47109241e-07 1.19527842e-08 8.47209241e-07 1.19527846e-08 8.47309241e-07 1.19527843e-08 8.47409241e-07 1.19527845e-08 8.47509241e-07 1.19527843e-08 8.47609241e-07 1.19527847e-08
+ 8.47709241e-07 1.19527846e-08 8.47809241e-07 1.19527844e-08 8.47909241e-07 1.19527846e-08 8.48009241e-07 1.19527844e-08 8.48109241e-07 1.19527849e-08 8.48209241e-07 1.19527847e-08 8.48309241e-07 1.19527848e-08 8.48409241e-07 1.19527847e-08
+ 8.48509241e-07 1.19527848e-08 8.48609241e-07 1.19527846e-08 8.48709241e-07 1.19527846e-08 8.48809241e-07 1.19527847e-08 8.48909241e-07 1.19527848e-08 8.49009241e-07 1.19527848e-08 8.49109241e-07 1.19527848e-08 8.49209241e-07 1.19527848e-08
+ 8.49309241e-07 1.19527846e-08 8.49409241e-07 1.19527851e-08 8.49509241e-07 1.19527847e-08 8.49609241e-07 1.19527853e-08 8.49709241e-07 1.19527847e-08 8.49809241e-07 1.19527852e-08 8.49909241e-07 1.19527852e-08 8.50009241e-07 1.19527853e-08
+ 8.50109241e-07 1.19527852e-08 8.50209241e-07 1.19527849e-08 8.50309241e-07 1.19527853e-08 8.50409241e-07 1.19527852e-08 8.50509241e-07 1.1952785e-08 8.50609241e-07 1.19527852e-08 8.50709241e-07 1.19527854e-08 8.50809241e-07 1.19527851e-08
+ 8.50909241e-07 1.19527856e-08 8.51e-07 1.19527852e-08 8.5101e-07 1.19386918e-08 8.5103e-07 1.20215821e-08 8.5107e-07 1.18440786e-08 8.5115e-07 1.2077572e-08 8.5125e-07 1.18225583e-08 8.5135e-07 1.2078315e-08
+ 8.5145e-07 1.18420536e-08 8.5155e-07 1.20411277e-08 8.5165e-07 1.18900523e-08 8.5175e-07 1.19863694e-08 8.5185e-07 1.19530395e-08 8.51930828e-07 1.24467922e-07 8.52e-07 1.72239017e-06 8.52008608e-07 -4.6155889e-06
+ 8.52025825e-07 -7.7865531e-06 8.52060258e-07 1.13509844e-06 8.52106181e-07 1.11144542e-05 8.52150081e-07 -1.1934542e-05 8.52198026e-07 9.08990105e-06 8.5225538e-07 -8.63563247e-06 8.52312019e-07 6.70440666e-06 8.52404232e-07 -4.84172578e-06
+ 8.52504232e-07 3.27464683e-06 8.52604232e-07 -1.93327282e-06 8.52704232e-07 9.69006195e-07 8.52804232e-07 -1.42030635e-07 8.52904232e-07 -5.08190821e-07 8.53004232e-07 1.1074106e-06 8.53104232e-07 -1.58170362e-06 8.53204232e-07 2.02780267e-06
+ 8.53304232e-07 -2.36191986e-06 8.53404232e-07 2.67940834e-06 8.53504232e-07 -2.89378902e-06 8.53604232e-07 3.10213512e-06 8.53704232e-07 -3.21656805e-06 8.53804232e-07 3.33567977e-06 8.53904232e-07 -3.37016818e-06 8.54004232e-07 3.41946247e-06
+ 8.54104232e-07 -3.39276677e-06 8.54204232e-07 3.38981241e-06 8.54304232e-07 -3.31838696e-06 8.54404232e-07 3.27818282e-06 8.54504232e-07 -3.175748e-06 8.54604232e-07 3.11054471e-06 8.54704232e-07 -2.98810251e-06 8.54804232e-07 2.90756109e-06
+ 8.54904232e-07 -2.77365299e-06 8.55004232e-07 2.68516151e-06 8.55104232e-07 -2.54622598e-06 8.55204232e-07 2.45527496e-06 8.55304232e-07 -2.31602352e-06 8.55404232e-07 2.22656391e-06 8.55504232e-07 -2.0903272e-06 8.55604232e-07 2.00509543e-06
+ 8.55704232e-07 -1.87412373e-06 8.55804232e-07 1.79491502e-06 8.55904232e-07 -1.67063204e-06 8.56004232e-07 1.59852859e-06 8.56104232e-07 -1.48173646e-06 8.56204232e-07 1.4172895e-06 8.56304232e-07 -1.30833291e-06 8.56404232e-07 1.25170759e-06
+ 8.56504232e-07 -1.15060305e-06 8.56604232e-07 1.10169152e-06 8.56704232e-07 -1.0082267e-06 8.56804232e-07 9.66733687e-07 8.56904232e-07 -8.80542186e-07 8.57004232e-07 8.46049289e-07 8.57104232e-07 -7.6666751e-07 8.57204232e-07 7.3868397e-07
+ 8.57304232e-07 -6.65596516e-07 8.57404232e-07 6.43597459e-07 8.57504232e-07 -5.76268889e-07 8.57604232e-07 5.59721194e-07 8.57704232e-07 -4.97617339e-07 8.57804232e-07 4.85996962e-07 8.57904232e-07 -4.28599301e-07 8.58004232e-07 4.21403053e-07
+ 8.58104232e-07 -3.68218431e-07 8.58204232e-07 3.64971765e-07 8.58304232e-07 -3.15538581e-07 8.58404232e-07 3.15800292e-07 8.58504232e-07 -2.69691964e-07 8.58604232e-07 2.73056533e-07 8.58704232e-07 -2.2988251e-07 8.58804232e-07 2.35978874e-07
+ 8.58904232e-07 -1.95381872e-07 8.59004232e-07 2.03872939e-07 8.59104232e-07 -1.65532531e-07 8.59204232e-07 1.76119e-07 8.59304232e-07 -1.39751474e-07 8.59404232e-07 1.52167858e-07 8.59504232e-07 -1.1752094e-07 8.59604232e-07 1.3153135e-07
+ 8.59704232e-07 -9.83820627e-08 8.59804232e-07 1.13778877e-07 8.59904232e-07 -8.19309294e-08 8.60004232e-07 9.8531214e-08 8.60104232e-07 -6.78117257e-08 8.60204232e-07 8.54545178e-08 8.60304232e-07 -5.57115593e-08 8.60404232e-07 7.42566393e-08
+ 8.60504232e-07 -4.5359055e-08 8.60604232e-07 6.46841334e-08 8.60704232e-07 -3.65163433e-08 8.60804232e-07 5.65134234e-08 8.60904232e-07 -2.89731026e-08 8.61004232e-07 4.95475203e-08 8.61104232e-07 -2.25458683e-08 8.61204232e-07 4.3615552e-08
+ 8.61304232e-07 -1.70756622e-08 8.61404232e-07 3.85696048e-08 8.61504232e-07 -1.24250063e-08 8.61604232e-07 3.42818967e-08 8.61704232e-07 -8.47524878e-09 8.61804232e-07 3.06422354e-08 8.61904232e-07 -5.1241329e-09 8.62004232e-07 2.75557194e-08
+ 8.62104232e-07 -2.28369379e-09 8.62204232e-07 2.494085e-08 8.62304232e-07 1.20663174e-10 8.62404232e-07 2.27293333e-08 8.62504232e-07 2.14064166e-09 8.62604232e-07 2.08840209e-08 8.62704232e-07 3.82602761e-09 8.62804232e-07 1.93450392e-08
+ 8.62904232e-07 5.23100624e-09 8.63004232e-07 1.80626871e-08 8.63104232e-07 6.40116757e-09 8.63204232e-07 1.69951489e-08 8.63304232e-07 7.37485339e-09 8.63404232e-07 1.61072773e-08 8.63504232e-07 8.18427445e-09 8.63604232e-07 1.53695615e-08
+ 8.63704232e-07 8.85646259e-09 8.63804232e-07 1.47572435e-08 8.63904232e-07 9.4140892e-09 8.64004232e-07 1.42496092e-08 8.64104232e-07 9.87609014e-09 8.64204232e-07 1.38293653e-08 8.64304232e-07 1.02579411e-08 8.64404232e-07 1.34824606e-08
+ 8.64504232e-07 1.05733336e-08 8.64604232e-07 1.31955877e-08 8.64704232e-07 1.08342035e-08 8.64804232e-07 1.29585628e-08 8.64904232e-07 1.1049393e-08 8.65004232e-07 1.27633174e-08 8.65104232e-07 1.12264359e-08 8.65204232e-07 1.26028726e-08
+ 8.65304232e-07 1.13717581e-08 8.65404232e-07 1.24713198e-08 8.65504232e-07 1.14908051e-08 8.65604232e-07 1.23635807e-08 8.65704232e-07 1.15882853e-08 8.65804232e-07 1.22755165e-08 8.65904232e-07 1.16676999e-08 8.66004232e-07 1.22039679e-08
+ 8.66104232e-07 1.17321324e-08 8.66204232e-07 1.21459758e-08 8.66304232e-07 1.17842887e-08 8.66404232e-07 1.20991124e-08 8.66504232e-07 1.18263538e-08 8.66604232e-07 1.20613944e-08 8.66704232e-07 1.18601353e-08 8.66804232e-07 1.20310981e-08
+ 8.66904232e-07 1.18872594e-08 8.67004232e-07 1.20070316e-08 8.67104232e-07 1.19085738e-08 8.67204232e-07 1.19880781e-08 8.67304232e-07 1.1925417e-08 8.67404232e-07 1.19731435e-08 8.67504232e-07 1.1938623e-08 8.67604232e-07 1.19615013e-08
+ 8.67704232e-07 1.19488514e-08 8.67804232e-07 1.19525492e-08 8.67904232e-07 1.19566547e-08 8.68004232e-07 1.19457785e-08 8.68104232e-07 1.19624982e-08 8.68204232e-07 1.19407656e-08 8.68304232e-07 1.19667684e-08 8.68404232e-07 1.19371593e-08
+ 8.68504232e-07 1.19697978e-08 8.68604232e-07 1.19346252e-08 8.68704232e-07 1.19718618e-08 8.68804232e-07 1.19330192e-08 8.68904232e-07 1.19730705e-08 8.69004232e-07 1.19321401e-08 8.69104232e-07 1.19736653e-08 8.69204232e-07 1.19317918e-08
+ 8.69304232e-07 1.19738028e-08 8.69404232e-07 1.19318361e-08 8.69504232e-07 1.1973595e-08 8.69604232e-07 1.19321918e-08 8.69704232e-07 1.1973111e-08 8.69804232e-07 1.19327847e-08 8.69904232e-07 1.19724274e-08 8.70004232e-07 1.19335432e-08
+ 8.70104232e-07 1.19716067e-08 8.70204232e-07 1.1934414e-08 8.70304232e-07 1.19706963e-08 8.70404232e-07 1.19353557e-08 8.70504232e-07 1.19697313e-08 8.70604232e-07 1.19363369e-08 8.70704232e-07 1.19687405e-08 8.70804232e-07 1.19373323e-08
+ 8.70904232e-07 1.19677451e-08 8.71004232e-07 1.19383236e-08 8.71104232e-07 1.19667617e-08 8.71204232e-07 1.19392961e-08 8.71304232e-07 1.19658027e-08 8.71404232e-07 1.19402395e-08 8.71504232e-07 1.19648765e-08 8.71604232e-07 1.1941147e-08
+ 8.71704232e-07 1.19639891e-08 8.71804232e-07 1.19420131e-08 8.71904232e-07 1.19631445e-08 8.72004232e-07 1.19428354e-08 8.72104232e-07 1.19623453e-08 8.72204232e-07 1.19436107e-08 8.72304232e-07 1.19615934e-08 8.72404232e-07 1.19443397e-08
+ 8.72504232e-07 1.19608878e-08 8.72604232e-07 1.19450219e-08 8.72704232e-07 1.19602288e-08 8.72804232e-07 1.19456583e-08 8.72904232e-07 1.19596146e-08 8.73004232e-07 1.19462507e-08 8.73104232e-07 1.19590441e-08 8.73204232e-07 1.19468001e-08
+ 8.73304232e-07 1.1958515e-08 8.73404232e-07 1.19473089e-08 8.73504232e-07 1.19580259e-08 8.73604232e-07 1.19477787e-08 8.73704232e-07 1.19575752e-08 8.73804232e-07 1.19482113e-08 8.73904232e-07 1.19571607e-08 8.74004232e-07 1.19486087e-08
+ 8.74104232e-07 1.19567795e-08 8.74204232e-07 1.19489735e-08 8.74304232e-07 1.19564303e-08 8.74404232e-07 1.1949308e-08 8.74504232e-07 1.19561108e-08 8.74604232e-07 1.19496138e-08 8.74704232e-07 1.1955818e-08 8.74804232e-07 1.19498936e-08
+ 8.74904232e-07 1.19555503e-08 8.75004232e-07 1.19501493e-08 8.75104232e-07 1.19553058e-08 8.75204232e-07 1.19503831e-08 8.75304232e-07 1.19550829e-08 8.75404232e-07 1.19505964e-08 8.75504232e-07 1.19548783e-08 8.75604232e-07 1.19507921e-08
+ 8.75704232e-07 1.19546915e-08 8.75804232e-07 1.19509708e-08 8.75904232e-07 1.19545207e-08 8.76004232e-07 1.19511337e-08 8.76104232e-07 1.19543651e-08 8.76204232e-07 1.1951282e-08 8.76304232e-07 1.19542242e-08 8.76404232e-07 1.19514164e-08
+ 8.76504232e-07 1.19540961e-08 8.76604232e-07 1.19515389e-08 8.76704232e-07 1.19539788e-08 8.76804232e-07 1.19516501e-08 8.76904232e-07 1.19538731e-08 8.77004232e-07 1.19517514e-08 8.77104232e-07 1.19537764e-08 8.77204232e-07 1.19518432e-08
+ 8.77304232e-07 1.19536883e-08 8.77404232e-07 1.19519276e-08 8.77504232e-07 1.19536083e-08 8.77604232e-07 1.19520037e-08 8.77704232e-07 1.19535355e-08 8.77804232e-07 1.19520732e-08 8.77904232e-07 1.19534692e-08 8.78004232e-07 1.19521367e-08
+ 8.78104232e-07 1.19534088e-08 8.78204232e-07 1.19521942e-08 8.78304232e-07 1.19533538e-08 8.78404232e-07 1.1952247e-08 8.78504232e-07 1.19533035e-08 8.78604232e-07 1.19522949e-08 8.78704232e-07 1.19532578e-08 8.78804232e-07 1.19523386e-08
+ 8.78904232e-07 1.19532158e-08 8.79004232e-07 1.19523784e-08 8.79104232e-07 1.19531782e-08 8.79204232e-07 1.19524149e-08 8.79304232e-07 1.19531433e-08 8.79404232e-07 1.19524479e-08 8.79504232e-07 1.19531118e-08 8.79604232e-07 1.19524782e-08
+ 8.79704232e-07 1.19530828e-08 8.79804232e-07 1.19525061e-08 8.79904232e-07 1.19530564e-08 8.80004232e-07 1.1952531e-08 8.80104232e-07 1.19530324e-08 8.80204232e-07 1.1952554e-08 8.80304232e-07 1.19530105e-08 8.80404232e-07 1.19525746e-08
+ 8.80504232e-07 1.19529909e-08 8.80604232e-07 1.19525937e-08 8.80704232e-07 1.19529724e-08 8.80804232e-07 1.19526111e-08 8.80904232e-07 1.19529559e-08 8.81004232e-07 1.19526271e-08 8.81104232e-07 1.1952941e-08 8.81204232e-07 1.19526412e-08
+ 8.81304232e-07 1.1952927e-08 8.81404232e-07 1.19526546e-08 8.81504232e-07 1.19529145e-08 8.81604232e-07 1.19526668e-08 8.81704232e-07 1.19529029e-08 8.81804232e-07 1.19526776e-08 8.81904232e-07 1.19528923e-08 8.82004232e-07 1.19526874e-08
+ 8.82104232e-07 1.19528829e-08 8.82204232e-07 1.19526967e-08 8.82304232e-07 1.19528742e-08 8.82404232e-07 1.1952705e-08 8.82504232e-07 1.19528661e-08 8.82604232e-07 1.19527124e-08 8.82704232e-07 1.1952859e-08 8.82804232e-07 1.19527194e-08
+ 8.82904232e-07 1.19528525e-08 8.83004232e-07 1.19527258e-08 8.83104232e-07 1.19528465e-08 8.83204232e-07 1.19527311e-08 8.83304232e-07 1.19528414e-08 8.83404232e-07 1.19527364e-08 8.83504232e-07 1.19528365e-08 8.83604232e-07 1.19527415e-08
+ 8.83704232e-07 1.19528318e-08 8.83804232e-07 1.19527457e-08 8.83904232e-07 1.19528277e-08 8.84004232e-07 1.19527493e-08 8.84104232e-07 1.19528241e-08 8.84204232e-07 1.19527531e-08 8.84304232e-07 1.19528209e-08 8.84404232e-07 1.19527559e-08
+ 8.84504232e-07 1.19528177e-08 8.84604232e-07 1.19527591e-08 8.84704232e-07 1.1952815e-08 8.84804232e-07 1.19527614e-08 8.84904232e-07 1.19528127e-08 8.85004232e-07 1.19527643e-08 8.85104232e-07 1.19528102e-08 8.85204232e-07 1.19527663e-08
+ 8.85304232e-07 1.19528082e-08 8.85404232e-07 1.19527684e-08 8.85504232e-07 1.19528061e-08 8.85604232e-07 1.19527703e-08 8.85704232e-07 1.19528042e-08 8.85804232e-07 1.19527717e-08 8.85904232e-07 1.19528026e-08 8.86004232e-07 1.19527734e-08
+ 8.86104232e-07 1.19528011e-08 8.86204232e-07 1.19527748e-08 8.86304232e-07 1.19528001e-08 8.86404232e-07 1.1952776e-08 8.86504232e-07 1.19527987e-08 8.86604232e-07 1.19527772e-08 8.86704232e-07 1.19527979e-08 8.86804232e-07 1.19527781e-08
+ 8.86904232e-07 1.19527971e-08 8.87004232e-07 1.19527788e-08 8.87104232e-07 1.19527962e-08 8.87204232e-07 1.19527798e-08 8.87304232e-07 1.19527953e-08 8.87404232e-07 1.19527808e-08 8.87504232e-07 1.19527946e-08 8.87604232e-07 1.19527812e-08
+ 8.87704232e-07 1.19527939e-08 8.87804232e-07 1.19527819e-08 8.87904232e-07 1.19527933e-08 8.88004232e-07 1.19527825e-08 8.88104232e-07 1.19527927e-08 8.88204232e-07 1.1952783e-08 8.88304232e-07 1.19527923e-08 8.88404232e-07 1.19527835e-08
+ 8.88504232e-07 1.19527919e-08 8.88604232e-07 1.19527838e-08 8.88704232e-07 1.19527913e-08 8.88804232e-07 1.19527843e-08 8.88904232e-07 1.19527911e-08 8.89004232e-07 1.19527845e-08 8.89104232e-07 1.19527908e-08 8.89204232e-07 1.19527846e-08
+ 8.89304232e-07 1.19527908e-08 8.89404232e-07 1.19527851e-08 8.89504232e-07 1.19527904e-08 8.89604232e-07 1.19527855e-08 8.89704232e-07 1.19527899e-08 8.89804232e-07 1.19527857e-08 8.89904232e-07 1.19527895e-08 8.90004232e-07 1.19527859e-08
+ 8.90104232e-07 1.19527896e-08 8.90204232e-07 1.19527862e-08 8.90304232e-07 1.19527894e-08 8.90404232e-07 1.19527862e-08 8.90504232e-07 1.19527892e-08 8.90604232e-07 1.19527863e-08 8.90704232e-07 1.19527893e-08 8.90804232e-07 1.19527866e-08
+ 8.90904232e-07 1.19527891e-08 8.91004232e-07 1.19527868e-08 8.91104232e-07 1.19527889e-08 8.91204232e-07 1.19527867e-08 8.91304232e-07 1.19527887e-08 8.91404232e-07 1.19527872e-08 8.91504232e-07 1.19527883e-08 8.91604232e-07 1.19527873e-08
+ 8.91704232e-07 1.19527882e-08 8.91804232e-07 1.19527873e-08 8.91904232e-07 1.19527884e-08 8.92004232e-07 1.19527872e-08 8.92104232e-07 1.19527884e-08 8.92204232e-07 1.19527875e-08 8.92304232e-07 1.19527883e-08 8.92404232e-07 1.19527874e-08
+ 8.92504232e-07 1.19527882e-08 8.92604232e-07 1.19527875e-08 8.92704232e-07 1.1952788e-08 8.92804232e-07 1.19527879e-08 8.92904232e-07 1.19527881e-08 8.93004232e-07 1.19527878e-08 8.93104232e-07 1.19527879e-08 8.93204232e-07 1.19527878e-08
+ 8.93304232e-07 1.1952788e-08 8.93404232e-07 1.19527875e-08 8.93504232e-07 1.19527881e-08 8.93604232e-07 1.19527878e-08 8.93704232e-07 1.1952788e-08 8.93804232e-07 1.19527877e-08 8.93904232e-07 1.19527881e-08 8.94004232e-07 1.19527876e-08
+ 8.94104232e-07 1.19527879e-08 8.94204232e-07 1.19527881e-08 8.94304232e-07 1.19527877e-08 8.94404232e-07 1.19527881e-08 8.94504232e-07 1.19527876e-08 8.94604232e-07 1.19527879e-08 8.94704232e-07 1.19527879e-08 8.94804232e-07 1.19527875e-08
+ 8.94904232e-07 1.19527879e-08 8.95004232e-07 1.19527879e-08 8.95104232e-07 1.19527876e-08 8.95204232e-07 1.1952788e-08 8.95304232e-07 1.19527882e-08 8.95404232e-07 1.19527876e-08 8.95504232e-07 1.19527879e-08 8.95604232e-07 1.19527878e-08
+ 8.95704232e-07 1.19527879e-08 8.95804232e-07 1.19527879e-08 8.95904232e-07 1.19527878e-08 8.96004232e-07 1.1952788e-08 8.96104232e-07 1.19527878e-08 8.96204232e-07 1.1952788e-08 8.96304232e-07 1.19527881e-08 8.96404232e-07 1.19527879e-08
+ 8.96504232e-07 1.19527879e-08 8.96604232e-07 1.19527877e-08 8.96704232e-07 1.19527879e-08 8.96804232e-07 1.1952788e-08 8.96904232e-07 1.19527881e-08 8.97004232e-07 1.19527877e-08 8.97104232e-07 1.19527882e-08 8.97204232e-07 1.19527875e-08
+ 8.97304232e-07 1.19527881e-08 8.97404232e-07 1.19527878e-08 8.97504232e-07 1.19527879e-08 8.97604232e-07 1.1952788e-08 8.97704232e-07 1.19527879e-08 8.97804232e-07 1.19527879e-08 8.97904232e-07 1.19527879e-08 8.98004232e-07 1.1952788e-08
+ 8.98104232e-07 1.19527878e-08 8.98204232e-07 1.1952788e-08 8.98304232e-07 1.19527877e-08 8.98404232e-07 1.19527882e-08 8.98504232e-07 1.19527878e-08 8.98604232e-07 1.19527883e-08 8.98704232e-07 1.19527877e-08 8.98804232e-07 1.1952788e-08
+ 8.98904232e-07 1.19527877e-08 8.99004232e-07 1.19527883e-08 8.99104232e-07 1.19527877e-08 8.99204232e-07 1.19527882e-08 8.99304232e-07 1.19527877e-08 8.99404232e-07 1.19527883e-08 8.99504232e-07 1.19527878e-08 8.99604232e-07 1.19527881e-08
+ 8.99704232e-07 1.19527878e-08 8.99804232e-07 1.19527879e-08 8.99904232e-07 1.19527877e-08 9e-07 1.19527882e-08 9.0001e-07 1.19897012e-08 9.0003e-07 1.17744015e-08 9.0007e-07 1.22290802e-08 9.0015e-07 1.16424027e-08
+ 9.0025e-07 1.22714108e-08 9.0035e-07 1.16453997e-08 9.0045e-07 1.22303623e-08 9.0055e-07 1.17276505e-08 9.0065e-07 1.18206769e-08 9.0075e-07 2.88720798e-08 9.0085e-07 -5.4410992e-07 9.00932051e-07 7.37313015e-06
+ 9.01e-07 -4.67316346e-05 9.01008488e-07 -5.13612331e-05 9.01025463e-07 -3.72346547e-05 9.01059414e-07 -3.10057984e-05 9.0109062e-07 0.000250461008 9.0114347e-07 0.00049480124 9.01199151e-07 0.00157091292 9.01299151e-07 -0.0175241145
+ 9.01399151e-07 0.171158646 9.01499151e-07 4.36372901 9.01599151e-07 5.20242883 9.01699151e-07 4.8824605 9.01799151e-07 5.06724446 9.01893327e-07 4.9583704 9.01993327e-07 5.0269427 9.02093327e-07 4.98189925
+ 9.02193327e-07 5.0121594 9.02293327e-07 4.99168783 9.02393327e-07 5.00564959 9.02493327e-07 4.99611607 9.02593327e-07 5.00265018 9.02693327e-07 4.99817445 9.02793327e-07 5.0012475 9.02893327e-07 4.99913996
+ 9.02993327e-07 5.00058806 9.03093327e-07 4.99959445 9.03193327e-07 5.0002773 9.03293327e-07 4.99980878 9.03393327e-07 5.00013066 9.03493327e-07 4.99990996 9.03593327e-07 5.00006141 9.03693327e-07 4.99995775
+ 9.03793327e-07 5.0000287 9.03893327e-07 4.99998031 9.03993327e-07 5.00001327 9.04093327e-07 4.99999095 9.04193327e-07 5.00000601 9.04293327e-07 4.99999594 9.04393327e-07 5.00000262 9.04493327e-07 4.99999825
+ 9.04593327e-07 5.00000105 9.04693327e-07 4.99999931 9.04793327e-07 5.00000035 9.04893327e-07 4.99999978 9.04993327e-07 5.00000005 9.05093327e-07 4.99999997 9.05193327e-07 4.99999993 9.05293327e-07 5.00000003
+ 9.05393327e-07 4.9999999 9.05493327e-07 5.00000005 9.05593327e-07 4.9999999 9.05693327e-07 5.00000004 9.05793327e-07 4.99999991 9.05893327e-07 5.00000002 9.05993327e-07 4.99999993 9.06093327e-07 5.00000001
+ 9.06193327e-07 4.99999994 9.06293327e-07 5.0 9.06393327e-07 4.99999995 9.06493327e-07 4.99999998 9.06593327e-07 4.99999996 9.06693327e-07 4.99999998 9.06793327e-07 4.99999997 9.06893327e-07 4.99999997
+ 9.06993327e-07 4.99999997 9.07093327e-07 4.99999997 9.07193327e-07 4.99999998 9.07293327e-07 4.99999996 9.07393327e-07 4.99999998 9.07493327e-07 4.99999996 9.07593327e-07 4.99999998 9.07693327e-07 4.99999996
+ 9.07793327e-07 4.99999998 9.07893327e-07 4.99999996 9.07993327e-07 4.99999998 9.08093327e-07 4.99999996 9.08193327e-07 4.99999998 9.08293327e-07 4.99999996 9.08393327e-07 4.99999998 9.08493327e-07 4.99999996
+ 9.08593327e-07 4.99999998 9.08693327e-07 4.99999996 9.08793327e-07 4.99999998 9.08893327e-07 4.99999996 9.08993327e-07 4.99999998 9.09093327e-07 4.99999996 9.09193327e-07 4.99999998 9.09293327e-07 4.99999997
+ 9.09393327e-07 4.99999998 9.09493327e-07 4.99999997 9.09593327e-07 4.99999998 9.09693327e-07 4.99999997 9.09793327e-07 4.99999998 9.09893327e-07 4.99999997 9.09993327e-07 4.99999998 9.10093327e-07 4.99999997
+ 9.10193327e-07 4.99999998 9.10293327e-07 4.99999997 9.10393327e-07 4.99999998 9.10493327e-07 4.99999997 9.10593327e-07 4.99999998 9.10693327e-07 4.99999997 9.10793327e-07 4.99999998 9.10893327e-07 4.99999997
+ 9.10993327e-07 4.99999997 9.11093327e-07 4.99999997 9.11193327e-07 4.99999997 9.11293327e-07 4.99999997 9.11393327e-07 4.99999997 9.11493327e-07 4.99999997 9.11593327e-07 4.99999997 9.11693327e-07 4.99999997
+ 9.11793327e-07 4.99999997 9.11893327e-07 4.99999997 9.11993327e-07 4.99999997 9.12093327e-07 4.99999997 9.12193327e-07 4.99999997 9.12293327e-07 4.99999997 9.12393327e-07 4.99999997 9.12493327e-07 4.99999997
+ 9.12593327e-07 4.99999997 9.12693327e-07 4.99999997 9.12793327e-07 4.99999997 9.12893327e-07 4.99999997 9.12993327e-07 4.99999997 9.13093327e-07 4.99999997 9.13193327e-07 4.99999997 9.13293327e-07 4.99999997
+ 9.13393327e-07 4.99999997 9.13493327e-07 4.99999997 9.13593327e-07 4.99999997 9.13693327e-07 4.99999997 9.13793327e-07 4.99999997 9.13893327e-07 4.99999997 9.13993327e-07 4.99999997 9.14093327e-07 4.99999997
+ 9.14193327e-07 4.99999997 9.14293327e-07 4.99999997 9.14393327e-07 4.99999997 9.14493327e-07 4.99999997 9.14593327e-07 4.99999997 9.14693327e-07 4.99999997 9.14793327e-07 4.99999997 9.14893327e-07 4.99999997
+ 9.14993327e-07 4.99999997 9.15093327e-07 4.99999997 9.15193327e-07 4.99999997 9.15293327e-07 4.99999997 9.15393327e-07 4.99999997 9.15493327e-07 4.99999997 9.15593327e-07 4.99999997 9.15693327e-07 4.99999997
+ 9.15793327e-07 4.99999997 9.15893327e-07 4.99999997 9.15993327e-07 4.99999997 9.16093327e-07 4.99999997 9.16193327e-07 4.99999997 9.16293327e-07 4.99999997 9.16393327e-07 4.99999997 9.16493327e-07 4.99999997
+ 9.16593327e-07 4.99999997 9.16693327e-07 4.99999997 9.16793327e-07 4.99999997 9.16893327e-07 4.99999997 9.16993327e-07 4.99999997 9.17093327e-07 4.99999997 9.17193327e-07 4.99999997 9.17293327e-07 4.99999997
+ 9.17393327e-07 4.99999997 9.17493327e-07 4.99999997 9.17593327e-07 4.99999997 9.17693327e-07 4.99999997 9.17793327e-07 4.99999997 9.17893327e-07 4.99999997 9.17993327e-07 4.99999997 9.18093327e-07 4.99999997
+ 9.18193327e-07 4.99999997 9.18293327e-07 4.99999997 9.18393327e-07 4.99999997 9.18493327e-07 4.99999997 9.18593327e-07 4.99999997 9.18693327e-07 4.99999997 9.18793327e-07 4.99999997 9.18893327e-07 4.99999997
+ 9.18993327e-07 4.99999997 9.19093327e-07 4.99999997 9.19193327e-07 4.99999997 9.19293327e-07 4.99999997 9.19393327e-07 4.99999997 9.19493327e-07 4.99999997 9.19593327e-07 4.99999997 9.19693327e-07 4.99999997
+ 9.19793327e-07 4.99999997 9.19893327e-07 4.99999997 9.19993327e-07 4.99999997 9.20093327e-07 4.99999997 9.20193327e-07 4.99999997 9.20293327e-07 4.99999997 9.20393327e-07 4.99999997 9.20493327e-07 4.99999997
+ 9.20593327e-07 4.99999997 9.20693327e-07 4.99999997 9.20793327e-07 4.99999997 9.20893327e-07 4.99999997 9.20993327e-07 4.99999997 9.21093327e-07 4.99999997 9.21193327e-07 4.99999997 9.21293327e-07 4.99999997
+ 9.21393327e-07 4.99999997 9.21493327e-07 4.99999997 9.21593327e-07 4.99999997 9.21693327e-07 4.99999997 9.21793327e-07 4.99999997 9.21893327e-07 4.99999997 9.21993327e-07 4.99999997 9.22093327e-07 4.99999997
+ 9.22193327e-07 4.99999997 9.22293327e-07 4.99999997 9.22393327e-07 4.99999997 9.22493327e-07 4.99999997 9.22593327e-07 4.99999997 9.22693327e-07 4.99999997 9.22793327e-07 4.99999997 9.22893327e-07 4.99999997
+ 9.22993327e-07 4.99999997 9.23093327e-07 4.99999997 9.23193327e-07 4.99999997 9.23293327e-07 4.99999997 9.23393327e-07 4.99999997 9.23493327e-07 4.99999997 9.23593327e-07 4.99999997 9.23693327e-07 4.99999997
+ 9.23793327e-07 4.99999997 9.23893327e-07 4.99999997 9.23993327e-07 4.99999997 9.24093327e-07 4.99999997 9.24193327e-07 4.99999997 9.24293327e-07 4.99999997 9.24393327e-07 4.99999997 9.24493327e-07 4.99999997
+ 9.24593327e-07 4.99999997 9.24693327e-07 4.99999997 9.24793327e-07 4.99999997 9.24893327e-07 4.99999997 9.24993327e-07 4.99999997 9.25093327e-07 4.99999997 9.25193327e-07 4.99999997 9.25293327e-07 4.99999997
+ 9.25393327e-07 4.99999997 9.25493327e-07 4.99999997 9.25593327e-07 4.99999997 9.25693327e-07 4.99999997 9.25793327e-07 4.99999997 9.25893327e-07 4.99999997 9.25993327e-07 4.99999997 9.26093327e-07 4.99999997
+ 9.26193327e-07 4.99999997 9.26293327e-07 4.99999997 9.26393327e-07 4.99999997 9.26493327e-07 4.99999997 9.26593327e-07 4.99999997 9.26693327e-07 4.99999997 9.26793327e-07 4.99999997 9.26893327e-07 4.99999997
+ 9.26993327e-07 4.99999997 9.27093327e-07 4.99999997 9.27193327e-07 4.99999997 9.27293327e-07 4.99999997 9.27393327e-07 4.99999997 9.27493327e-07 4.99999997 9.27593327e-07 4.99999997 9.27693327e-07 4.99999997
+ 9.27793327e-07 4.99999997 9.27893327e-07 4.99999997 9.27993327e-07 4.99999997 9.28093327e-07 4.99999997 9.28193327e-07 4.99999997 9.28293327e-07 4.99999997 9.28393327e-07 4.99999997 9.28493327e-07 4.99999997
+ 9.28593327e-07 4.99999997 9.28693327e-07 4.99999997 9.28793327e-07 4.99999997 9.28893327e-07 4.99999997 9.28993327e-07 4.99999997 9.29093327e-07 4.99999997 9.29193327e-07 4.99999997 9.29293327e-07 4.99999997
+ 9.29393327e-07 4.99999997 9.29493327e-07 4.99999997 9.29593327e-07 4.99999997 9.29693327e-07 4.99999997 9.29793327e-07 4.99999997 9.29893327e-07 4.99999997 9.29993327e-07 4.99999997 9.30093327e-07 4.99999997
+ 9.30193327e-07 4.99999997 9.30293327e-07 4.99999997 9.30393327e-07 4.99999997 9.30493327e-07 4.99999997 9.30593327e-07 4.99999997 9.30693327e-07 4.99999997 9.30793327e-07 4.99999997 9.30893327e-07 4.99999997
+ 9.30993327e-07 4.99999997 9.31093327e-07 4.99999997 9.31193327e-07 4.99999997 9.31293327e-07 4.99999997 9.31393327e-07 4.99999997 9.31493327e-07 4.99999997 9.31593327e-07 4.99999997 9.31693327e-07 4.99999997
+ 9.31793327e-07 4.99999997 9.31893327e-07 4.99999997 9.31993327e-07 4.99999997 9.32093327e-07 4.99999997 9.32193327e-07 4.99999997 9.32293327e-07 4.99999997 9.32393327e-07 4.99999997 9.32493327e-07 4.99999997
+ 9.32593327e-07 4.99999997 9.32693327e-07 4.99999997 9.32793327e-07 4.99999997 9.32893327e-07 4.99999997 9.32993327e-07 4.99999997 9.33093327e-07 4.99999997 9.33193327e-07 4.99999997 9.33293327e-07 4.99999997
+ 9.33393327e-07 4.99999997 9.33493327e-07 4.99999997 9.33593327e-07 4.99999997 9.33693327e-07 4.99999997 9.33793327e-07 4.99999997 9.33893327e-07 4.99999997 9.33993327e-07 4.99999997 9.34093327e-07 4.99999997
+ 9.34193327e-07 4.99999997 9.34293327e-07 4.99999997 9.34393327e-07 4.99999997 9.34493327e-07 4.99999997 9.34593327e-07 4.99999997 9.34693327e-07 4.99999997 9.34793327e-07 4.99999997 9.34893327e-07 4.99999997
+ 9.34993327e-07 4.99999997 9.35093327e-07 4.99999997 9.35193327e-07 4.99999997 9.35293327e-07 4.99999997 9.35393327e-07 4.99999997 9.35493327e-07 4.99999997 9.35593327e-07 4.99999997 9.35693327e-07 4.99999997
+ 9.35793327e-07 4.99999997 9.35893327e-07 4.99999997 9.35993327e-07 4.99999997 9.36093327e-07 4.99999997 9.36193327e-07 4.99999997 9.36293327e-07 4.99999997 9.36393327e-07 4.99999997 9.36493327e-07 4.99999997
+ 9.36593327e-07 4.99999997 9.36693327e-07 4.99999997 9.36793327e-07 4.99999997 9.36893327e-07 4.99999997 9.36993327e-07 4.99999997 9.37093327e-07 4.99999997 9.37193327e-07 4.99999997 9.37293327e-07 4.99999997
+ 9.37393327e-07 4.99999997 9.37493327e-07 4.99999997 9.37593327e-07 4.99999997 9.37693327e-07 4.99999997 9.37793327e-07 4.99999997 9.37893327e-07 4.99999997 9.37993327e-07 4.99999997 9.38093327e-07 4.99999997
+ 9.38193327e-07 4.99999997 9.38293327e-07 4.99999997 9.38393327e-07 4.99999997 9.38493327e-07 4.99999997 9.38593327e-07 4.99999997 9.38693327e-07 4.99999997 9.38793327e-07 4.99999997 9.38893327e-07 4.99999997
+ 9.38993327e-07 4.99999997 9.39093327e-07 4.99999997 9.39193327e-07 4.99999997 9.39293327e-07 4.99999997 9.39393327e-07 4.99999997 9.39493327e-07 4.99999997 9.39593327e-07 4.99999997 9.39693327e-07 4.99999997
+ 9.39793327e-07 4.99999997 9.39893327e-07 4.99999997 9.39993327e-07 4.99999997 9.40093327e-07 4.99999997 9.40193327e-07 4.99999997 9.40293327e-07 4.99999997 9.40393327e-07 4.99999997 9.40493327e-07 4.99999997
+ 9.40593327e-07 4.99999997 9.40693327e-07 4.99999997 9.40793327e-07 4.99999997 9.40893327e-07 4.99999997 9.40993327e-07 4.99999997 9.41093327e-07 4.99999997 9.41193327e-07 4.99999997 9.41293327e-07 4.99999997
+ 9.41393327e-07 4.99999997 9.41493327e-07 4.99999997 9.41593327e-07 4.99999997 9.41693327e-07 4.99999997 9.41793327e-07 4.99999997 9.41893327e-07 4.99999997 9.41993327e-07 4.99999997 9.42093327e-07 4.99999997
+ 9.42193327e-07 4.99999997 9.42293327e-07 4.99999997 9.42393327e-07 4.99999997 9.42493327e-07 4.99999997 9.42593327e-07 4.99999997 9.42693327e-07 4.99999997 9.42793327e-07 4.99999997 9.42893327e-07 4.99999997
+ 9.42993327e-07 4.99999997 9.43093327e-07 4.99999997 9.43193327e-07 4.99999997 9.43293327e-07 4.99999997 9.43393327e-07 4.99999997 9.43493327e-07 4.99999997 9.43593327e-07 4.99999997 9.43693327e-07 4.99999997
+ 9.43793327e-07 4.99999997 9.43893327e-07 4.99999997 9.43993327e-07 4.99999997 9.44093327e-07 4.99999997 9.44193327e-07 4.99999997 9.44293327e-07 4.99999997 9.44393327e-07 4.99999997 9.44493327e-07 4.99999997
+ 9.44593327e-07 4.99999997 9.44693327e-07 4.99999997 9.44793327e-07 4.99999997 9.44893327e-07 4.99999997 9.44993327e-07 4.99999997 9.45093327e-07 4.99999997 9.45193327e-07 4.99999997 9.45293327e-07 4.99999997
+ 9.45393327e-07 4.99999997 9.45493327e-07 4.99999997 9.45593327e-07 4.99999997 9.45693327e-07 4.99999997 9.45793327e-07 4.99999997 9.45893327e-07 4.99999997 9.45993327e-07 4.99999997 9.46093327e-07 4.99999997
+ 9.46193327e-07 4.99999997 9.46293327e-07 4.99999997 9.46393327e-07 4.99999997 9.46493327e-07 4.99999997 9.46593327e-07 4.99999997 9.46693327e-07 4.99999997 9.46793327e-07 4.99999997 9.46893327e-07 4.99999997
+ 9.46993327e-07 4.99999997 9.47093327e-07 4.99999997 9.47193327e-07 4.99999997 9.47293327e-07 4.99999997 9.47393327e-07 4.99999997 9.47493327e-07 4.99999997 9.47593327e-07 4.99999997 9.47693327e-07 4.99999997
+ 9.47793327e-07 4.99999997 9.47893327e-07 4.99999997 9.47993327e-07 4.99999997 9.48093327e-07 4.99999997 9.48193327e-07 4.99999997 9.48293327e-07 4.99999997 9.48393327e-07 4.99999997 9.48493327e-07 4.99999997
+ 9.48593327e-07 4.99999997 9.48693327e-07 4.99999997 9.48793327e-07 4.99999997 9.48893327e-07 4.99999997 9.48993327e-07 4.99999997 9.49093327e-07 4.99999997 9.49193327e-07 4.99999997 9.49293327e-07 4.99999997
+ 9.49393327e-07 4.99999997 9.49493327e-07 4.99999997 9.49593327e-07 4.99999997 9.49693327e-07 4.99999997 9.49793327e-07 4.99999997 9.49893327e-07 4.99999997 9.49993327e-07 4.99999997 9.50093327e-07 4.99999997
+ 9.50193327e-07 4.99999997 9.50293327e-07 4.99999997 9.50393327e-07 4.99999997 9.50493327e-07 4.99999997 9.50593327e-07 4.99999997 9.50693327e-07 4.99999997 9.50793327e-07 4.99999997 9.50893327e-07 4.99999997
+ 9.50993327e-07 4.99999997 9.51e-07 4.99999997 9.5101e-07 4.99999997 9.5103e-07 4.99999997 9.5107e-07 4.99999997 9.5115e-07 4.99999997 9.5125e-07 4.99999997 9.5135e-07 4.99999997
+ 9.5145e-07 4.99999997 9.5155e-07 4.99999997 9.5165e-07 4.99999997 9.5175e-07 4.99999997 9.5185e-07 4.99999997 9.51930828e-07 5.00000065 9.52e-07 5.00000149 9.52008608e-07 4.99999288
+ 9.52025825e-07 4.99997549 9.52060258e-07 4.99999257 9.52106188e-07 5.00004375 9.52150118e-07 5.00000856 9.5219811e-07 4.99994581 9.52255501e-07 5.00002983 9.52312176e-07 4.99999321 9.52404431e-07 5.00000355
+ 9.52490774e-07 5.00000011 9.52590774e-07 4.99999756 9.52690774e-07 5.00000329 9.52790774e-07 4.99999639 9.52890774e-07 5.0000034 9.52990774e-07 4.99999687 9.53090774e-07 5.00000266 9.53190774e-07 4.9999977
+ 9.53290774e-07 5.00000186 9.53390774e-07 4.99999842 9.53490774e-07 5.00000123 9.53590774e-07 4.99999895 9.53690774e-07 5.00000079 9.53790774e-07 4.99999931 9.53890774e-07 5.00000051 9.53990774e-07 4.99999954
+ 9.54090774e-07 5.00000033 9.54190774e-07 4.99999968 9.54290774e-07 5.00000021 9.54390774e-07 4.99999977 9.54490774e-07 5.00000014 9.54590774e-07 4.99999983 9.54690774e-07 5.00000009 9.54790774e-07 4.99999987
+ 9.54890774e-07 5.00000007 9.54990774e-07 4.99999989 9.55090774e-07 5.00000005 9.55190774e-07 4.99999991 9.55290774e-07 5.00000003 9.55390774e-07 4.99999992 9.55490774e-07 5.00000002 9.55590774e-07 4.99999993
+ 9.55690774e-07 5.00000001 9.55790774e-07 4.99999993 9.55890774e-07 5.00000001 9.55990774e-07 4.99999994 9.56090774e-07 5.0 9.56190774e-07 4.99999994 9.56290774e-07 5.0 9.56390774e-07 4.99999995
+ 9.56490774e-07 5.0 9.56590774e-07 4.99999995 9.56690774e-07 4.99999999 9.56790774e-07 4.99999995 9.56890774e-07 4.99999999 9.56990774e-07 4.99999996 9.57090774e-07 4.99999999 9.57190774e-07 4.99999996
+ 9.57290774e-07 4.99999999 9.57390774e-07 4.99999996 9.57490774e-07 4.99999998 9.57590774e-07 4.99999996 9.57690774e-07 4.99999998 9.57790774e-07 4.99999996 9.57890774e-07 4.99999998 9.57990774e-07 4.99999996
+ 9.58090774e-07 4.99999998 9.58190774e-07 4.99999997 9.58290774e-07 4.99999998 9.58390774e-07 4.99999997 9.58490774e-07 4.99999998 9.58590774e-07 4.99999997 9.58690774e-07 4.99999998 9.58790774e-07 4.99999997
+ 9.58890774e-07 4.99999998 9.58990774e-07 4.99999997 9.59090774e-07 4.99999998 9.59190774e-07 4.99999997 9.59290774e-07 4.99999997 9.59390774e-07 4.99999997 9.59490774e-07 4.99999997 9.59590774e-07 4.99999997
+ 9.59690774e-07 4.99999997 9.59790774e-07 4.99999997 9.59890774e-07 4.99999997 9.59990774e-07 4.99999997 9.60090774e-07 4.99999997 9.60190774e-07 4.99999997 9.60290774e-07 4.99999997 9.60390774e-07 4.99999997
+ 9.60490774e-07 4.99999997 9.60590774e-07 4.99999997 9.60690774e-07 4.99999997 9.60790774e-07 4.99999997 9.60890774e-07 4.99999997 9.60990774e-07 4.99999997 9.61090774e-07 4.99999997 9.61190774e-07 4.99999997
+ 9.61290774e-07 4.99999997 9.61390774e-07 4.99999997 9.61490774e-07 4.99999997 9.61590774e-07 4.99999997 9.61690774e-07 4.99999997 9.61790774e-07 4.99999997 9.61890774e-07 4.99999997 9.61990774e-07 4.99999997
+ 9.62090774e-07 4.99999997 9.62190774e-07 4.99999997 9.62290774e-07 4.99999997 9.62390774e-07 4.99999997 9.62490774e-07 4.99999997 9.62590774e-07 4.99999997 9.62690774e-07 4.99999997 9.62790774e-07 4.99999997
+ 9.62890774e-07 4.99999997 9.62990774e-07 4.99999997 9.63090774e-07 4.99999997 9.63190774e-07 4.99999997 9.63290774e-07 4.99999997 9.63390774e-07 4.99999997 9.63490774e-07 4.99999997 9.63590774e-07 4.99999997
+ 9.63690774e-07 4.99999997 9.63790774e-07 4.99999997 9.63890774e-07 4.99999997 9.63990774e-07 4.99999997 9.64090774e-07 4.99999997 9.64190774e-07 4.99999997 9.64290774e-07 4.99999997 9.64390774e-07 4.99999997
+ 9.64490774e-07 4.99999997 9.64590774e-07 4.99999997 9.64690774e-07 4.99999997 9.64790774e-07 4.99999997 9.64890774e-07 4.99999997 9.64990774e-07 4.99999997 9.65090774e-07 4.99999997 9.65190774e-07 4.99999997
+ 9.65290774e-07 4.99999997 9.65390774e-07 4.99999997 9.65490774e-07 4.99999997 9.65590774e-07 4.99999997 9.65690774e-07 4.99999997 9.65790774e-07 4.99999997 9.65890774e-07 4.99999997 9.65990774e-07 4.99999997
+ 9.66090774e-07 4.99999997 9.66190774e-07 4.99999997 9.66290774e-07 4.99999997 9.66390774e-07 4.99999997 9.66490774e-07 4.99999997 9.66590774e-07 4.99999997 9.66690774e-07 4.99999997 9.66790774e-07 4.99999997
+ 9.66890774e-07 4.99999997 9.66990774e-07 4.99999997 9.67090774e-07 4.99999997 9.67190774e-07 4.99999997 9.67290774e-07 4.99999997 9.67390774e-07 4.99999997 9.67490774e-07 4.99999997 9.67590774e-07 4.99999997
+ 9.67690774e-07 4.99999997 9.67790774e-07 4.99999997 9.67890774e-07 4.99999997 9.67990774e-07 4.99999997 9.68090774e-07 4.99999997 9.68190774e-07 4.99999997 9.68290774e-07 4.99999997 9.68390774e-07 4.99999997
+ 9.68490774e-07 4.99999997 9.68590774e-07 4.99999997 9.68690774e-07 4.99999997 9.68790774e-07 4.99999997 9.68890774e-07 4.99999997 9.68990774e-07 4.99999997 9.69090774e-07 4.99999997 9.69190774e-07 4.99999997
+ 9.69290774e-07 4.99999997 9.69390774e-07 4.99999997 9.69490774e-07 4.99999997 9.69590774e-07 4.99999997 9.69690774e-07 4.99999997 9.69790774e-07 4.99999997 9.69890774e-07 4.99999997 9.69990774e-07 4.99999997
+ 9.70090774e-07 4.99999997 9.70190774e-07 4.99999997 9.70290774e-07 4.99999997 9.70390774e-07 4.99999997 9.70490774e-07 4.99999997 9.70590774e-07 4.99999997 9.70690774e-07 4.99999997 9.70790774e-07 4.99999997
+ 9.70890774e-07 4.99999997 9.70990774e-07 4.99999997 9.71090774e-07 4.99999997 9.71190774e-07 4.99999997 9.71290774e-07 4.99999997 9.71390774e-07 4.99999997 9.71490774e-07 4.99999997 9.71590774e-07 4.99999997
+ 9.71690774e-07 4.99999997 9.71790774e-07 4.99999997 9.71890774e-07 4.99999997 9.71990774e-07 4.99999997 9.72090774e-07 4.99999997 9.72190774e-07 4.99999997 9.72290774e-07 4.99999997 9.72390774e-07 4.99999997
+ 9.72490774e-07 4.99999997 9.72590774e-07 4.99999997 9.72690774e-07 4.99999997 9.72790774e-07 4.99999997 9.72890774e-07 4.99999997 9.72990774e-07 4.99999997 9.73090774e-07 4.99999997 9.73190774e-07 4.99999997
+ 9.73290774e-07 4.99999997 9.73390774e-07 4.99999997 9.73490774e-07 4.99999997 9.73590774e-07 4.99999997 9.73690774e-07 4.99999997 9.73790774e-07 4.99999997 9.73890774e-07 4.99999997 9.73990774e-07 4.99999997
+ 9.74090774e-07 4.99999997 9.74190774e-07 4.99999997 9.74290774e-07 4.99999997 9.74390774e-07 4.99999997 9.74490774e-07 4.99999997 9.74590774e-07 4.99999997 9.74690774e-07 4.99999997 9.74790774e-07 4.99999997
+ 9.74890774e-07 4.99999997 9.74990774e-07 4.99999997 9.75090774e-07 4.99999997 9.75190774e-07 4.99999997 9.75290774e-07 4.99999997 9.75390774e-07 4.99999997 9.75490774e-07 4.99999997 9.75590774e-07 4.99999997
+ 9.75690774e-07 4.99999997 9.75790774e-07 4.99999997 9.75890774e-07 4.99999997 9.75990774e-07 4.99999997 9.76090774e-07 4.99999997 9.76190774e-07 4.99999997 9.76290774e-07 4.99999997 9.76390774e-07 4.99999997
+ 9.76490774e-07 4.99999997 9.76590774e-07 4.99999997 9.76690774e-07 4.99999997 9.76790774e-07 4.99999997 9.76890774e-07 4.99999997 9.76990774e-07 4.99999997 9.77090774e-07 4.99999997 9.77190774e-07 4.99999997
+ 9.77290774e-07 4.99999997 9.77390774e-07 4.99999997 9.77490774e-07 4.99999997 9.77590774e-07 4.99999997 9.77690774e-07 4.99999997 9.77790774e-07 4.99999997 9.77890774e-07 4.99999997 9.77990774e-07 4.99999997
+ 9.78090774e-07 4.99999997 9.78190774e-07 4.99999997 9.78290774e-07 4.99999997 9.78390774e-07 4.99999997 9.78490774e-07 4.99999997 9.78590774e-07 4.99999997 9.78690774e-07 4.99999997 9.78790774e-07 4.99999997
+ 9.78890774e-07 4.99999997 9.78990774e-07 4.99999997 9.79090774e-07 4.99999997 9.79190774e-07 4.99999997 9.79290774e-07 4.99999997 9.79390774e-07 4.99999997 9.79490774e-07 4.99999997 9.79590774e-07 4.99999997
+ 9.79690774e-07 4.99999997 9.79790774e-07 4.99999997 9.79890774e-07 4.99999997 9.79990774e-07 4.99999997 9.80090774e-07 4.99999997 9.80190774e-07 4.99999997 9.80290774e-07 4.99999997 9.80390774e-07 4.99999997
+ 9.80490774e-07 4.99999997 9.80590774e-07 4.99999997 9.80690774e-07 4.99999997 9.80790774e-07 4.99999997 9.80890774e-07 4.99999997 9.80990774e-07 4.99999997 9.81090774e-07 4.99999997 9.81190774e-07 4.99999997
+ 9.81290774e-07 4.99999997 9.81390774e-07 4.99999997 9.81490774e-07 4.99999997 9.81590774e-07 4.99999997 9.81690774e-07 4.99999997 9.81790774e-07 4.99999997 9.81890774e-07 4.99999997 9.81990774e-07 4.99999997
+ 9.82090774e-07 4.99999997 9.82190774e-07 4.99999997 9.82290774e-07 4.99999997 9.82390774e-07 4.99999997 9.82490774e-07 4.99999997 9.82590774e-07 4.99999997 9.82690774e-07 4.99999997 9.82790774e-07 4.99999997
+ 9.82890774e-07 4.99999997 9.82990774e-07 4.99999997 9.83090774e-07 4.99999997 9.83190774e-07 4.99999997 9.83290774e-07 4.99999997 9.83390774e-07 4.99999997 9.83490774e-07 4.99999997 9.83590774e-07 4.99999997
+ 9.83690774e-07 4.99999997 9.83790774e-07 4.99999997 9.83890774e-07 4.99999997 9.83990774e-07 4.99999997 9.84090774e-07 4.99999997 9.84190774e-07 4.99999997 9.84290774e-07 4.99999997 9.84390774e-07 4.99999997
+ 9.84490774e-07 4.99999997 9.84590774e-07 4.99999997 9.84690774e-07 4.99999997 9.84790774e-07 4.99999997 9.84890774e-07 4.99999997 9.84990774e-07 4.99999997 9.85090774e-07 4.99999997 9.85190774e-07 4.99999997
+ 9.85290774e-07 4.99999997 9.85390774e-07 4.99999997 9.85490774e-07 4.99999997 9.85590774e-07 4.99999997 9.85690774e-07 4.99999997 9.85790774e-07 4.99999997 9.85890774e-07 4.99999997 9.85990774e-07 4.99999997
+ 9.86090774e-07 4.99999997 9.86190774e-07 4.99999997 9.86290774e-07 4.99999997 9.86390774e-07 4.99999997 9.86490774e-07 4.99999997 9.86590774e-07 4.99999997 9.86690774e-07 4.99999997 9.86790774e-07 4.99999997
+ 9.86890774e-07 4.99999997 9.86990774e-07 4.99999997 9.87090774e-07 4.99999997 9.87190774e-07 4.99999997 9.87290774e-07 4.99999997 9.87390774e-07 4.99999997 9.87490774e-07 4.99999997 9.87590774e-07 4.99999997
+ 9.87690774e-07 4.99999997 9.87790774e-07 4.99999997 9.87890774e-07 4.99999997 9.87990774e-07 4.99999997 9.88090774e-07 4.99999997 9.88190774e-07 4.99999997 9.88290774e-07 4.99999997 9.88390774e-07 4.99999997
+ 9.88490774e-07 4.99999997 9.88590774e-07 4.99999997 9.88690774e-07 4.99999997 9.88790774e-07 4.99999997 9.88890774e-07 4.99999997 9.88990774e-07 4.99999997 9.89090774e-07 4.99999997 9.89190774e-07 4.99999997
+ 9.89290774e-07 4.99999997 9.89390774e-07 4.99999997 9.89490774e-07 4.99999997 9.89590774e-07 4.99999997 9.89690774e-07 4.99999997 9.89790774e-07 4.99999997 9.89890774e-07 4.99999997 9.89990774e-07 4.99999997
+ 9.90090774e-07 4.99999997 9.90190774e-07 4.99999997 9.90290774e-07 4.99999997 9.90390774e-07 4.99999997 9.90490774e-07 4.99999997 9.90590774e-07 4.99999997 9.90690774e-07 4.99999997 9.90790774e-07 4.99999997
+ 9.90890774e-07 4.99999997 9.90990774e-07 4.99999997 9.91090774e-07 4.99999997 9.91190774e-07 4.99999997 9.91290774e-07 4.99999997 9.91390774e-07 4.99999997 9.91490774e-07 4.99999997 9.91590774e-07 4.99999997
+ 9.91690774e-07 4.99999997 9.91790774e-07 4.99999997 9.91890774e-07 4.99999997 9.91990774e-07 4.99999997 9.92090774e-07 4.99999997 9.92190774e-07 4.99999997 9.92290774e-07 4.99999997 9.92390774e-07 4.99999997
+ 9.92490774e-07 4.99999997 9.92590774e-07 4.99999997 9.92690774e-07 4.99999997 9.92790774e-07 4.99999997 9.92890774e-07 4.99999997 9.92990774e-07 4.99999997 9.93090774e-07 4.99999997 9.93190774e-07 4.99999997
+ 9.93290774e-07 4.99999997 9.93390774e-07 4.99999997 9.93490774e-07 4.99999997 9.93590774e-07 4.99999997 9.93690774e-07 4.99999997 9.93790774e-07 4.99999997 9.93890774e-07 4.99999997 9.93990774e-07 4.99999997
+ 9.94090774e-07 4.99999997 9.94190774e-07 4.99999997 9.94290774e-07 4.99999997 9.94390774e-07 4.99999997 9.94490774e-07 4.99999997 9.94590774e-07 4.99999997 9.94690774e-07 4.99999997 9.94790774e-07 4.99999997
+ 9.94890774e-07 4.99999997 9.94990774e-07 4.99999997 9.95090774e-07 4.99999997 9.95190774e-07 4.99999997 9.95290774e-07 4.99999997 9.95390774e-07 4.99999997 9.95490774e-07 4.99999997 9.95590774e-07 4.99999997
+ 9.95690774e-07 4.99999997 9.95790774e-07 4.99999997 9.95890774e-07 4.99999997 9.95990774e-07 4.99999997 9.96090774e-07 4.99999997 9.96190774e-07 4.99999997 9.96290774e-07 4.99999997 9.96390774e-07 4.99999997
+ 9.96490774e-07 4.99999997 9.96590774e-07 4.99999997 9.96690774e-07 4.99999997 9.96790774e-07 4.99999997 9.96890774e-07 4.99999997 9.96990774e-07 4.99999997 9.97090774e-07 4.99999997 9.97190774e-07 4.99999997
+ 9.97290774e-07 4.99999997 9.97390774e-07 4.99999997 9.97490774e-07 4.99999997 9.97590774e-07 4.99999997 9.97690774e-07 4.99999997 9.97790774e-07 4.99999997 9.97890774e-07 4.99999997 9.97990774e-07 4.99999997
+ 9.98090774e-07 4.99999997 9.98190774e-07 4.99999997 9.98290774e-07 4.99999997 9.98390774e-07 4.99999997 9.98490774e-07 4.99999997 9.98590774e-07 4.99999997 9.98690774e-07 4.99999997 9.98790774e-07 4.99999997
+ 9.98890774e-07 4.99999997 9.98990774e-07 4.99999997 9.99090774e-07 4.99999997 9.99190774e-07 4.99999997 9.99290774e-07 4.99999997 9.99390774e-07 4.99999997 9.99490774e-07 4.99999997 9.99590774e-07 4.99999997
+ 9.99690774e-07 4.99999997 9.99790774e-07 4.99999997 9.99890774e-07 4.99999997 9.99990774e-07 4.99999997 1e-06 4.99999997 )

Vclkin4 in4 0 PWL( 0.0 1.19527881e-08 1e-12 1.23894446e-08 2e-12 1.24174266e-08 4e-12 1.21116663e-08 8e-12 1.13794303e-08 1.6e-11 1.18656753e-08 3.2e-11 1.22917884e-08 6.4e-11 1.1678974e-08
+ 1.28e-10 1.21533428e-08 2.28e-10 1.17980896e-08 3.28e-10 1.2069907e-08 4.28e-10 1.1863019e-08 5.28e-10 1.2027713e-08 6.28e-10 1.18447033e-08 7.28e-10 1.33402875e-08 8.17641203e-10 -3.51137717e-07
+ 8.87939724e-10 1.69691292e-06 9.63955785e-10 -5.72246145e-07 1e-09 -1.66556126e-05 1.00713579e-09 6.15865114e-06 1.02140738e-09 1.08591792e-05 1.04995055e-09 -1.72985475e-06 1.09557449e-09 9.85015735e-07 1.1454732e-09 -2.35135568e-06
+ 1.21884515e-09 1.93427741e-06 1.31884515e-09 -1.56725203e-06 1.41884515e-09 1.42053732e-06 1.51884515e-09 -1.29153738e-06 1.61884515e-09 1.24059975e-06 1.71884515e-09 -1.14817918e-06 1.81884515e-09 1.10462298e-06 1.91884515e-09 -1.01248979e-06
+ 2.01884515e-09 9.69196536e-07 2.11884515e-09 -8.79158158e-07 2.21884515e-09 8.39755508e-07 2.31884515e-09 -7.54990385e-07 2.41884515e-09 7.21675266e-07 2.51884515e-09 -6.43510101e-07 2.61884515e-09 6.16928946e-07 2.71884515e-09 -5.45534834e-07
+ 2.81884515e-09 5.2553402e-07 2.91884515e-09 -4.60540353e-07 3.01884515e-09 4.46615506e-07 3.11884515e-09 -3.87430672e-07 3.21884515e-09 3.78949005e-07 3.31884515e-09 -3.24915778e-07 3.41884515e-09 3.21223059e-07 3.51884515e-09 -2.71693049e-07
+ 3.61884515e-09 2.72164341e-07 3.71884515e-09 -2.25108271e-07 3.81884515e-09 2.32304069e-07 3.91884515e-09 -1.86991202e-07 4.01884515e-09 1.96862543e-07 4.11884515e-09 -1.54899068e-07 4.21884515e-09 1.66952856e-07 4.31884515e-09 -1.27839239e-07
+ 4.41884515e-09 1.41754699e-07 4.51884515e-09 -1.05062071e-07 4.61884515e-09 1.20558949e-07 4.71884515e-09 -8.59130108e-08 4.81884515e-09 1.02748528e-07 4.91884515e-09 -6.98318334e-08 5.01884515e-09 8.77996248e-08 5.11884515e-09 -5.63414924e-08
+ 5.21884515e-09 7.52653132e-08 5.31884515e-09 -4.5033854e-08 5.41884515e-09 6.47624625e-08 5.51884515e-09 -3.55618028e-08 5.61884515e-09 5.59670932e-08 5.71884515e-09 -2.76316835e-08 5.81884515e-09 4.8605104e-08 5.91884515e-09 -2.09952443e-08
+ 6.01884515e-09 4.24452808e-08 6.11884515e-09 -1.54294007e-08 6.21884515e-09 3.7280064e-08 6.31884515e-09 -1.0789148e-08 6.41884515e-09 3.29740449e-08 6.51884515e-09 -6.90923999e-09 6.61884515e-09 2.93742507e-08 6.71884515e-09 -3.665898e-09
+ 6.81884515e-09 2.63652905e-08 6.91884515e-09 -9.55089785e-10 7.01884515e-09 2.38505689e-08 7.11884515e-09 1.31027658e-09 7.21884515e-09 2.17662708e-08 7.31884515e-09 3.1886426e-09 7.41884515e-09 2.00484184e-08 7.51884515e-09 4.73720968e-09
+ 7.61884515e-09 1.86322537e-08 7.71884515e-09 6.01376088e-09 7.81884515e-09 1.74648971e-08 7.91884515e-09 7.06599182e-09 8.01884515e-09 1.65027064e-08 8.11884515e-09 7.93326302e-09 8.21884515e-09 1.57096708e-08 8.31884515e-09 8.64804753e-09
+ 8.41884515e-09 1.49587278e-08 8.51884515e-09 9.22329019e-09 8.61884515e-09 1.44312957e-08 8.71884515e-09 9.70221403e-09 8.81884515e-09 1.39963748e-08 8.91884515e-09 1.00971634e-08 9.01884515e-09 1.36377309e-08 9.11884515e-09 1.04228352e-08
+ 9.21884515e-09 1.33420031e-08 9.31884515e-09 1.0691369e-08 9.41884515e-09 1.30981648e-08 9.51884515e-09 1.09127822e-08 9.61884515e-09 1.28971152e-08 9.71884515e-09 1.10953403e-08 9.81884515e-09 1.27313488e-08 9.91884515e-09 1.12458588e-08
+ 1.00188451e-08 1.25946757e-08 1.01188451e-08 1.13699596e-08 1.02188451e-08 1.24819913e-08 1.03188451e-08 1.14722774e-08 1.04188451e-08 1.23890866e-08 1.05188451e-08 1.1556635e-08 1.06188451e-08 1.23124901e-08 1.07188451e-08 1.16261838e-08
+ 1.08188451e-08 1.224934e-08 1.09188451e-08 1.16835243e-08 1.10188451e-08 1.21972755e-08 1.11188451e-08 1.1730798e-08 1.12188451e-08 1.21543513e-08 1.13188451e-08 1.17697728e-08 1.14188451e-08 1.21189629e-08 1.15188451e-08 1.1801905e-08
+ 1.16188451e-08 1.20897873e-08 1.17188451e-08 1.18283959e-08 1.18188451e-08 1.20657338e-08 1.19188451e-08 1.18502358e-08 1.20188451e-08 1.20459034e-08 1.21188451e-08 1.18682418e-08 1.22188451e-08 1.20295547e-08 1.23188451e-08 1.18830861e-08
+ 1.24188451e-08 1.20160763e-08 1.25188451e-08 1.18953241e-08 1.26188451e-08 1.20049644e-08 1.27188451e-08 1.19054134e-08 1.28188451e-08 1.19958035e-08 1.29188451e-08 1.19137315e-08 1.30188451e-08 1.19882508e-08 1.31188451e-08 1.19205889e-08
+ 1.32188451e-08 1.19820247e-08 1.33188451e-08 1.19262425e-08 1.34188451e-08 1.1976891e-08 1.35188451e-08 1.19309038e-08 1.36188451e-08 1.1972659e-08 1.37188451e-08 1.19347462e-08 1.38188451e-08 1.19691702e-08 1.39188451e-08 1.19379137e-08
+ 1.40188451e-08 1.19662938e-08 1.41188451e-08 1.19405256e-08 1.42188451e-08 1.19639226e-08 1.43188451e-08 1.19426785e-08 1.44188451e-08 1.19619678e-08 1.45188451e-08 1.19444537e-08 1.46188451e-08 1.1960356e-08 1.47188451e-08 1.19459169e-08
+ 1.48188451e-08 1.19590272e-08 1.49188451e-08 1.19471234e-08 1.50188451e-08 1.19579321e-08 1.51188451e-08 1.1948118e-08 1.52188451e-08 1.19570286e-08 1.53188451e-08 1.19489383e-08 1.54188451e-08 1.1956284e-08 1.55188451e-08 1.19496142e-08
+ 1.56188451e-08 1.19556702e-08 1.57188451e-08 1.19501715e-08 1.58188451e-08 1.19551645e-08 1.59188451e-08 1.19506309e-08 1.60188451e-08 1.19547471e-08 1.61188451e-08 1.19510097e-08 1.62188451e-08 1.19544032e-08 1.63188451e-08 1.19513218e-08
+ 1.64188451e-08 1.19541198e-08 1.65188451e-08 1.19515793e-08 1.66188451e-08 1.19538859e-08 1.67188451e-08 1.19517918e-08 1.68188451e-08 1.19536933e-08 1.69188451e-08 1.19519666e-08 1.70188451e-08 1.19535342e-08 1.71188451e-08 1.19521106e-08
+ 1.72188451e-08 1.19534035e-08 1.73188451e-08 1.19522297e-08 1.74188451e-08 1.19532954e-08 1.75188451e-08 1.19523278e-08 1.76188451e-08 1.19532064e-08 1.77188451e-08 1.19524086e-08 1.78188451e-08 1.1953133e-08 1.79188451e-08 1.1952475e-08
+ 1.80188451e-08 1.19530727e-08 1.81188451e-08 1.19525299e-08 1.82188451e-08 1.19530228e-08 1.83188451e-08 1.19525753e-08 1.84188451e-08 1.19529817e-08 1.85188451e-08 1.19526127e-08 1.86188451e-08 1.19529475e-08 1.87188451e-08 1.19526435e-08
+ 1.88188451e-08 1.19529199e-08 1.89188451e-08 1.19526689e-08 1.90188451e-08 1.19528966e-08 1.91188451e-08 1.19526898e-08 1.92188451e-08 1.19528774e-08 1.93188451e-08 1.19527071e-08 1.94188451e-08 1.19528619e-08 1.95188451e-08 1.19527215e-08
+ 1.96188451e-08 1.19528488e-08 1.97188451e-08 1.19527334e-08 1.98188451e-08 1.19528382e-08 1.99188451e-08 1.19527427e-08 2e-08 1.19528287e-08 2.001e-08 4.54031335e-07 2.003e-08 -9.19688854e-07 2.007e-08 1.19439415e-07
+ 2.01e-08 1.33572873e-06 2.0108e-08 5.99959798e-06 2.0124e-08 9.93708622e-06 2.0156e-08 -8.6544918e-07 2.02150599e-08 -1.47787294e-05 2.02823902e-08 1.18571353e-05 2.03483061e-08 -9.63323815e-06 2.04483061e-08 1.67908448e-05
+ 2.05483061e-08 -2.08172021e-05 2.06483061e-08 2.06230284e-05 2.07483061e-08 -1.965003e-05 2.08483061e-08 1.83922363e-05 2.09483061e-08 -1.69351531e-05 2.10483061e-08 1.55120607e-05 2.11483061e-08 -1.40717308e-05 2.12483061e-08 1.27658979e-05
+ 2.13483061e-08 -1.14962806e-05 2.14483061e-08 1.03826023e-05 2.15483061e-08 -9.31242413e-06 2.16483061e-08 8.39272718e-06 2.17483061e-08 -7.50853974e-06 2.18483061e-08 6.76139193e-06 2.19483061e-08 -6.03770187e-06 2.20483061e-08 5.43648682e-06
+ 2.21483061e-08 -4.84666088e-06 2.22483061e-08 4.3659831e-06 2.23483061e-08 -3.88595196e-06 2.24483061e-08 3.50363252e-06 2.25483061e-08 -3.11284873e-06 2.26483061e-08 2.81025237e-06 2.27483061e-08 -2.49164944e-06 2.28483061e-08 2.25342153e-06
+ 2.29483061e-08 -1.99301809e-06 2.30483061e-08 1.80663484e-06 2.31483061e-08 -1.5930663e-06 2.32483061e-08 1.44837213e-06 2.33483061e-08 -1.27244403e-06 2.34483061e-08 1.16124557e-06 2.35483061e-08 -1.01554201e-06 2.36483061e-08 9.31224721e-07
+ 2.37483061e-08 -8.0977571e-07 2.38483061e-08 7.47023863e-07 2.39483061e-08 -6.45024483e-07 2.40483061e-08 5.99561945e-07 2.41483061e-08 -5.1315224e-07 2.42483061e-08 4.81544511e-07 2.43483061e-08 -4.07623885e-07 2.44483061e-08 3.87112686e-07
+ 2.45483061e-08 -3.23193719e-07 2.46483061e-08 3.1156849e-07 2.47483061e-08 -2.55658066e-07 2.48483061e-08 2.51147335e-07 2.49483061e-08 -2.0164823e-07 2.50483061e-08 2.02832493e-07 2.51483061e-08 -1.58465007e-07 2.52483061e-08 1.64207117e-07
+ 2.53483061e-08 -1.23946182e-07 2.54483061e-08 1.33335282e-07 2.55483061e-08 -9.63598259e-08 2.56483061e-08 1.08666353e-07 2.57483061e-08 -7.43188344e-08 2.58483061e-08 8.9538709e-08 2.59483061e-08 -5.62635895e-08 2.60483061e-08 7.36930547e-08
+ 2.61483061e-08 -4.22903585e-08 2.62483061e-08 6.10255795e-08 2.63483061e-08 -3.11379366e-08 2.64483061e-08 5.0913021e-08 2.65483061e-08 -2.22356416e-08 2.66483061e-08 4.2841942e-08 2.67483061e-08 -1.51314873e-08 2.68483061e-08 3.64016745e-08
+ 2.69483061e-08 -9.46309861e-09 2.70483061e-08 3.12639364e-08 2.71483061e-08 -4.94229727e-09 2.72483061e-08 2.71669083e-08 2.73483061e-08 -1.33743749e-09 2.74483061e-08 2.39001492e-08 2.75483061e-08 1.53673338e-09 2.76483061e-08 2.131567e-08
+ 2.77483061e-08 3.8110759e-09 2.78483061e-08 1.92848506e-08 2.79483061e-08 5.59808663e-09 2.80483061e-08 1.76899048e-08 2.81483061e-08 7.00089725e-09 2.82483061e-08 1.64384759e-08 2.83483061e-08 8.10098288e-09 2.84483061e-08 1.54577404e-08
+ 2.85483061e-08 8.96253552e-09 2.86483061e-08 1.45949781e-08 2.87483061e-08 9.62342941e-09 2.88483061e-08 1.40054847e-08 2.89483061e-08 1.01447451e-08 2.90483061e-08 1.35445587e-08 2.91483061e-08 1.05521442e-08 2.92483061e-08 1.31845844e-08
+ 2.93483061e-08 1.08701093e-08 2.94483061e-08 1.29038272e-08 2.95483061e-08 1.11177308e-08 2.96483061e-08 1.26856773e-08 2.97483061e-08 1.13100731e-08 2.98483061e-08 1.25159527e-08 2.99483061e-08 1.14597701e-08 3.00483061e-08 1.23840332e-08
+ 3.01483061e-08 1.15758833e-08 3.02483061e-08 1.2281875e-08 3.03483061e-08 1.16657727e-08 3.04483061e-08 1.22028316e-08 3.05483061e-08 1.1735211e-08 3.06483061e-08 1.21418779e-08 3.07483061e-08 1.17886773e-08 3.08483061e-08 1.20950147e-08
+ 3.09483061e-08 1.182972e-08 3.10483061e-08 1.20590998e-08 3.11483061e-08 1.18611207e-08 3.12483061e-08 1.20316695e-08 3.13483061e-08 1.18850622e-08 3.14483061e-08 1.20107931e-08 3.15483061e-08 1.19032426e-08 3.16483061e-08 1.19949838e-08
+ 3.17483061e-08 1.19169711e-08 3.18483061e-08 1.19830776e-08 3.19483061e-08 1.19272835e-08 3.20483061e-08 1.19741591e-08 3.21483061e-08 1.19349833e-08 3.22483061e-08 1.19675241e-08 3.23483061e-08 1.19406895e-08 3.24483061e-08 1.19626273e-08
+ 3.25483061e-08 1.19448805e-08 3.26483061e-08 1.19590505e-08 3.27483061e-08 1.19479229e-08 3.28483061e-08 1.19564725e-08 3.29483061e-08 1.19500996e-08 3.30483061e-08 1.19546419e-08 3.31483061e-08 1.19516317e-08 3.32483061e-08 1.19533671e-08
+ 3.33483061e-08 1.19526847e-08 3.34483061e-08 1.19525046e-08 3.35483061e-08 1.19533841e-08 3.36483061e-08 1.19519449e-08 3.37483061e-08 1.19538248e-08 3.38483061e-08 1.1951605e-08 3.39483061e-08 1.19540792e-08 3.40483061e-08 1.19514224e-08
+ 3.41483061e-08 1.19542017e-08 3.42483061e-08 1.19513499e-08 3.43483061e-08 1.19542333e-08 3.44483061e-08 1.19513524e-08 3.45483061e-08 1.19542029e-08 3.46483061e-08 1.1951405e-08 3.47483061e-08 1.1954133e-08 3.48483061e-08 1.19514887e-08
+ 3.49483061e-08 1.1954039e-08 3.50483061e-08 1.19515899e-08 3.51483061e-08 1.19539326e-08 3.52483061e-08 1.1951699e-08 3.53483061e-08 1.1953822e-08 3.54483061e-08 1.19518101e-08 3.55483061e-08 1.19537122e-08 3.56483061e-08 1.1951918e-08
+ 3.57483061e-08 1.19536067e-08 3.58483061e-08 1.19520204e-08 3.59483061e-08 1.19535076e-08 3.60483061e-08 1.19521155e-08 3.61483061e-08 1.19534164e-08 3.62483061e-08 1.19522029e-08 3.63483061e-08 1.19533335e-08 3.64483061e-08 1.19522813e-08
+ 3.65483061e-08 1.19532593e-08 3.66483061e-08 1.19523512e-08 3.67483061e-08 1.19531937e-08 3.68483061e-08 1.19524132e-08 3.69483061e-08 1.19531351e-08 3.70483061e-08 1.19524677e-08 3.71483061e-08 1.19530844e-08 3.72483061e-08 1.19525151e-08
+ 3.73483061e-08 1.19530401e-08 3.74483061e-08 1.19525561e-08 3.75483061e-08 1.19530021e-08 3.76483061e-08 1.19525916e-08 3.77483061e-08 1.19529695e-08 3.78483061e-08 1.1952622e-08 3.79483061e-08 1.19529412e-08 3.80483061e-08 1.19526479e-08
+ 3.81483061e-08 1.19529172e-08 3.82483061e-08 1.19526699e-08 3.83483061e-08 1.19528968e-08 3.84483061e-08 1.19526888e-08 3.85483061e-08 1.19528794e-08 3.86483061e-08 1.19527047e-08 3.87483061e-08 1.19528648e-08 3.88483061e-08 1.19527181e-08
+ 3.89483061e-08 1.19528523e-08 3.90483061e-08 1.19527296e-08 3.91483061e-08 1.19528421e-08 3.92483061e-08 1.1952739e-08 3.93483061e-08 1.19528334e-08 3.94483061e-08 1.19527473e-08 3.95483061e-08 1.19528257e-08 3.96483061e-08 1.19527539e-08
+ 3.97483061e-08 1.19528197e-08 3.98483061e-08 1.19527598e-08 3.99483061e-08 1.19528144e-08 4.00483061e-08 1.19527646e-08 4.01483061e-08 1.195281e-08 4.02483061e-08 1.19527686e-08 4.03483061e-08 1.19528064e-08 4.04483061e-08 1.19527718e-08
+ 4.05483061e-08 1.19528034e-08 4.06483061e-08 1.19527747e-08 4.07483061e-08 1.19528007e-08 4.08483061e-08 1.1952777e-08 4.09483061e-08 1.19527989e-08 4.10483061e-08 1.19527788e-08 4.11483061e-08 1.19527969e-08 4.12483061e-08 1.19527805e-08
+ 4.13483061e-08 1.19527955e-08 4.14483061e-08 1.19527818e-08 4.15483061e-08 1.19527941e-08 4.16483061e-08 1.19527831e-08 4.17483061e-08 1.1952793e-08 4.18483061e-08 1.1952784e-08 4.19483061e-08 1.19527921e-08 4.20483061e-08 1.19527849e-08
+ 4.21483061e-08 1.19527913e-08 4.22483061e-08 1.19527856e-08 4.23483061e-08 1.1952791e-08 4.24483061e-08 1.1952786e-08 4.25483061e-08 1.19527902e-08 4.26483061e-08 1.19527864e-08 4.27483061e-08 1.19527899e-08 4.28483061e-08 1.19527866e-08
+ 4.29483061e-08 1.19527896e-08 4.30483061e-08 1.19527871e-08 4.31483061e-08 1.19527896e-08 4.32483061e-08 1.19527872e-08 4.33483061e-08 1.19527892e-08 4.34483061e-08 1.19527873e-08 4.35483061e-08 1.19527893e-08 4.36483061e-08 1.19527873e-08
+ 4.37483061e-08 1.19527891e-08 4.38483061e-08 1.19527875e-08 4.39483061e-08 1.19527891e-08 4.40483061e-08 1.19527876e-08 4.41483061e-08 1.19527888e-08 4.42483061e-08 1.19527878e-08 4.43483061e-08 1.19527887e-08 4.44483061e-08 1.19527879e-08
+ 4.45483061e-08 1.1952789e-08 4.46483061e-08 1.19527877e-08 4.47483061e-08 1.19527888e-08 4.48483061e-08 1.19527877e-08 4.49483061e-08 1.19527891e-08 4.50483061e-08 1.19527876e-08 4.51483061e-08 1.19527889e-08 4.52483061e-08 1.19527877e-08
+ 4.53483061e-08 1.19527888e-08 4.54483061e-08 1.19527878e-08 4.55483061e-08 1.1952789e-08 4.56483061e-08 1.19527876e-08 4.57483061e-08 1.19527888e-08 4.58483061e-08 1.19527879e-08 4.59483061e-08 1.19527889e-08 4.60483061e-08 1.19527877e-08
+ 4.61483061e-08 1.19527888e-08 4.62483061e-08 1.19527878e-08 4.63483061e-08 1.1952789e-08 4.64483061e-08 1.19527878e-08 4.65483061e-08 1.1952789e-08 4.66483061e-08 1.19527878e-08 4.67483061e-08 1.1952789e-08 4.68483061e-08 1.19527879e-08
+ 4.69483061e-08 1.19527889e-08 4.70483061e-08 1.1952788e-08 4.71483061e-08 1.19527888e-08 4.72483061e-08 1.19527878e-08 4.73483061e-08 1.19527888e-08 4.74483061e-08 1.19527881e-08 4.75483061e-08 1.19527887e-08 4.76483061e-08 1.1952788e-08
+ 4.77483061e-08 1.19527885e-08 4.78483061e-08 1.19527878e-08 4.79483061e-08 1.19527886e-08 4.80483061e-08 1.19527879e-08 4.81483061e-08 1.19527886e-08 4.82483061e-08 1.19527881e-08 4.83483061e-08 1.19527887e-08 4.84483061e-08 1.1952788e-08
+ 4.85483061e-08 1.19527887e-08 4.86483061e-08 1.19527879e-08 4.87483061e-08 1.19527886e-08 4.88483061e-08 1.19527881e-08 4.89483061e-08 1.19527887e-08 4.90483061e-08 1.1952788e-08 4.91483061e-08 1.19527888e-08 4.92483061e-08 1.19527879e-08
+ 4.93483061e-08 1.19527888e-08 4.94483061e-08 1.19527878e-08 4.95483061e-08 1.19527889e-08 4.96483061e-08 1.19527878e-08 4.97483061e-08 1.1952789e-08 4.98483061e-08 1.19527876e-08 4.99483061e-08 1.1952789e-08 5.00483061e-08 1.19527877e-08
+ 5.01483061e-08 1.19527891e-08 5.02483061e-08 1.19527877e-08 5.03483061e-08 1.19527891e-08 5.04483061e-08 1.19527876e-08 5.05483061e-08 1.1952789e-08 5.06483061e-08 1.19527876e-08 5.07483061e-08 1.1952789e-08 5.08483061e-08 1.19527878e-08
+ 5.09483061e-08 1.1952789e-08 5.1e-08 1.19527875e-08 5.101e-08 1.19392991e-08 5.103e-08 1.20184647e-08 5.107e-08 1.18497342e-08 5.115e-08 1.20699984e-08 5.125e-08 1.18320609e-08 5.135e-08 1.20670217e-08
+ 5.145e-08 1.18546077e-08 5.155e-08 1.20278828e-08 5.165e-08 1.19035409e-08 5.175e-08 1.1973316e-08 5.185e-08 1.19649727e-08 5.19308282e-08 1.89258373e-07 5.2e-08 2.60151236e-07 5.20086083e-08 -7.14363737e-06
+ 5.2025825e-08 -6.95176104e-06 5.20602584e-08 1.22749827e-05 5.21061808e-08 -2.31708097e-07 5.21500808e-08 -6.86343727e-06 5.21980262e-08 -7.31793064e-07 5.22553803e-08 5.62213537e-06 5.23120186e-08 -4.8074731e-06 5.24042316e-08 3.76475686e-06
+ 5.25042316e-08 -3.03544165e-06 5.26042316e-08 2.49411106e-06 5.27042316e-08 -2.00984843e-06 5.28042316e-08 1.66794373e-06 5.29042316e-08 -1.35001926e-06 5.30042316e-08 1.14114027e-06 5.31042316e-08 -9.29894509e-07 5.32042316e-08 8.04845249e-07
+ 5.33042316e-08 -6.60306738e-07 5.34042316e-08 5.87542323e-07 5.35042316e-08 -4.84637649e-07 5.36042316e-08 4.4459476e-07 5.37042316e-08 -3.67852556e-07 5.38042316e-08 3.48473083e-07 5.39042316e-08 -2.88325344e-07 5.40042316e-08 2.82115808e-07
+ 5.41042316e-08 -2.32624698e-07 5.42042316e-08 2.34943424e-07 5.43042316e-08 -1.92413165e-07 5.44042316e-08 2.00347253e-07 5.45042316e-08 -1.62432568e-07 5.46042316e-08 1.74124235e-07 5.47042316e-08 -1.39330015e-07 5.48042316e-08 1.53591658e-07
+ 5.49042316e-08 -1.2095803e-07 5.50042316e-08 1.37022712e-07 5.51042316e-08 -1.0592632e-07 5.52042316e-08 1.23292891e-07 5.53042316e-08 -9.33235999e-08 5.54042316e-08 1.11659789e-07 5.55042316e-08 -8.25434371e-08 5.56042316e-08 1.01625211e-07
+ 5.57042316e-08 -7.31746015e-08 5.58042316e-08 9.2846256e-08 5.59042316e-08 -6.49299889e-08 5.60042316e-08 8.50824931e-08 5.61042316e-08 -5.76076953e-08 5.62042316e-08 7.81618226e-08 5.63042316e-08 -5.10595458e-08 5.64042316e-08 7.19558248e-08
+ 5.65042316e-08 -4.51736107e-08 5.66042316e-08 6.63661036e-08 5.67042316e-08 -3.98628736e-08 5.68042316e-08 6.1315114e-08 5.69042316e-08 -3.50580536e-08 5.70042316e-08 5.67411617e-08 5.71042316e-08 -3.07043376e-08 5.72042316e-08 5.25949753e-08
+ 5.73042316e-08 -2.67565805e-08 5.74042316e-08 4.88340739e-08 5.75042316e-08 -2.31741426e-08 5.76042316e-08 4.54196842e-08 5.77042316e-08 -1.99203326e-08 5.78042316e-08 4.23178497e-08 5.79042316e-08 -1.69644787e-08 5.80042316e-08 3.94999291e-08
+ 5.81042316e-08 -1.42788637e-08 5.82042316e-08 3.69391616e-08 5.83042316e-08 -1.18376721e-08 5.84042316e-08 3.46109255e-08 5.85042316e-08 -9.61771707e-09 5.86042316e-08 3.2493336e-08 5.87042316e-08 -7.59832e-09 5.88042316e-08 3.05667707e-08
+ 5.89042316e-08 -5.7607481e-09 5.90042316e-08 2.88133344e-08 5.91042316e-08 -4.08805068e-09 5.92042316e-08 2.72170516e-08 5.93042316e-08 -2.56516575e-09 5.94042316e-08 2.57636961e-08 5.95042316e-08 -1.17864715e-09 5.96042316e-08 2.44405289e-08
+ 5.97042316e-08 8.30635283e-11 5.98042316e-08 2.32370241e-08 5.99042316e-08 1.22373989e-09 6.00042316e-08 2.21552592e-08 6.01042316e-08 2.24987651e-09 6.02042316e-08 2.11816668e-08 6.03042316e-08 3.17381954e-09 6.04042316e-08 2.03046547e-08
+ 6.05042316e-08 4.00645458e-09 6.06042316e-08 1.95139946e-08 6.07042316e-08 4.75739864e-09 6.08042316e-08 1.88006402e-08 6.09042316e-08 5.43516571e-09 6.10042316e-08 1.81565751e-08 6.11042316e-08 6.0473061e-09 6.12042316e-08 1.75746841e-08
+ 6.13042316e-08 6.6005276e-09 6.14042316e-08 1.70486417e-08 6.15042316e-08 7.10079767e-09 6.16042316e-08 1.65728156e-08 6.17042316e-08 7.55343396e-09 6.18042316e-08 1.61421844e-08 6.19042316e-08 7.96317995e-09 6.20042316e-08 1.57522654e-08
+ 6.21042316e-08 8.33427238e-09 6.22042316e-08 1.53990533e-08 6.23042316e-08 8.6704984e-09 6.24042316e-08 1.50789661e-08 6.25042316e-08 8.97524777e-09 6.26042316e-08 1.47887982e-08 6.27042316e-08 9.25154531e-09 6.28042316e-08 1.45257079e-08
+ 6.29042316e-08 9.50205054e-09 6.30042316e-08 1.4287196e-08 6.31042316e-08 9.72913938e-09 6.32042316e-08 1.40709807e-08 6.33042316e-08 9.93499988e-09 6.34042316e-08 1.3874989e-08 6.35042316e-08 1.01215867e-08 6.36042316e-08 1.36973622e-08
+ 6.37042316e-08 1.02906836e-08 6.38042316e-08 1.35363784e-08 6.39042316e-08 1.04439535e-08 6.40042316e-08 1.33906269e-08 6.41042316e-08 1.05823832e-08 6.42042316e-08 1.32591181e-08 6.43042316e-08 1.07073398e-08 6.44042316e-08 1.31401034e-08
+ 6.45042316e-08 1.08210732e-08 6.46042316e-08 1.30313816e-08 6.47042316e-08 1.09248979e-08 6.48042316e-08 1.29323184e-08 6.49042316e-08 1.10193644e-08 6.50042316e-08 1.28422571e-08 6.51042316e-08 1.11052355e-08 6.52042316e-08 1.27603821e-08
+ 6.53042316e-08 1.11832529e-08 6.54042316e-08 1.26860943e-08 6.55042316e-08 1.12539986e-08 6.56042316e-08 1.26184633e-08 6.57042316e-08 1.13187881e-08 6.58042316e-08 1.2556781e-08 6.59042316e-08 1.13772567e-08 6.60042316e-08 1.25012838e-08
+ 6.61042316e-08 1.14300049e-08 6.62042316e-08 1.24511002e-08 6.63042316e-08 1.14777794e-08 6.64042316e-08 1.24056e-08 6.65042316e-08 1.15211252e-08 6.66042316e-08 1.23642986e-08 6.67042316e-08 1.15604834e-08 6.68042316e-08 1.23267886e-08
+ 6.69042316e-08 1.15962348e-08 6.70042316e-08 1.22927119e-08 6.71042316e-08 1.16287152e-08 6.72042316e-08 1.22617511e-08 6.73042316e-08 1.16582681e-08 6.74042316e-08 1.22334815e-08 6.75042316e-08 1.16852742e-08 6.76042316e-08 1.22077809e-08
+ 6.77042316e-08 1.17097037e-08 6.78042316e-08 1.21845376e-08 6.79042316e-08 1.17318351e-08 6.80042316e-08 1.21634536e-08 6.81042316e-08 1.17519279e-08 6.82042316e-08 1.21443018e-08 6.83042316e-08 1.17701857e-08 6.84042316e-08 1.21268952e-08
+ 6.85042316e-08 1.17867817e-08 6.86042316e-08 1.21110708e-08 6.87042316e-08 1.18018708e-08 6.88042316e-08 1.20966832e-08 6.89042316e-08 1.18155888e-08 6.90042316e-08 1.20836038e-08 6.91042316e-08 1.18280601e-08 6.92042316e-08 1.20717127e-08
+ 6.93042316e-08 1.18393979e-08 6.94042316e-08 1.20609019e-08 6.95042316e-08 1.1849706e-08 6.96042316e-08 1.20510733e-08 6.97042316e-08 1.18590776e-08 6.98042316e-08 1.20421373e-08 6.99042316e-08 1.18675976e-08 7.00042316e-08 1.20340134e-08
+ 7.01042316e-08 1.1875344e-08 7.02042316e-08 1.20266282e-08 7.03042316e-08 1.18823859e-08 7.04042316e-08 1.20199133e-08 7.05042316e-08 1.18887879e-08 7.06042316e-08 1.20138091e-08 7.07042316e-08 1.18946082e-08 7.08042316e-08 1.20082595e-08
+ 7.09042316e-08 1.18998998e-08 7.10042316e-08 1.20032143e-08 7.11042316e-08 1.19047101e-08 7.12042316e-08 1.19986273e-08 7.13042316e-08 1.19090842e-08 7.14042316e-08 1.19944567e-08 7.15042316e-08 1.19130606e-08 7.16042316e-08 1.19906658e-08
+ 7.17042316e-08 1.19166753e-08 7.18042316e-08 1.19872193e-08 7.19042316e-08 1.19199609e-08 7.20042316e-08 1.19840864e-08 7.21042316e-08 1.19229479e-08 7.22042316e-08 1.19812386e-08 7.23042316e-08 1.19256631e-08 7.24042316e-08 1.19786499e-08
+ 7.25042316e-08 1.19281313e-08 7.26042316e-08 1.19762963e-08 7.27042316e-08 1.19303752e-08 7.28042316e-08 1.1974157e-08 7.29042316e-08 1.19324154e-08 7.30042316e-08 1.19722117e-08 7.31042316e-08 1.19342695e-08 7.32042316e-08 1.19704439e-08
+ 7.33042316e-08 1.19359556e-08 7.34042316e-08 1.19688364e-08 7.35042316e-08 1.19374882e-08 7.36042316e-08 1.19673751e-08 7.37042316e-08 1.19388816e-08 7.38042316e-08 1.19660468e-08 7.39042316e-08 1.19401479e-08 7.40042316e-08 1.19648392e-08
+ 7.41042316e-08 1.19412992e-08 7.42042316e-08 1.19637417e-08 7.43042316e-08 1.1942346e-08 7.44042316e-08 1.19627437e-08 7.45042316e-08 1.19432972e-08 7.46042316e-08 1.19618364e-08 7.47042316e-08 1.19441622e-08 7.48042316e-08 1.19610119e-08
+ 7.49042316e-08 1.19449487e-08 7.50042316e-08 1.19602623e-08 7.51042316e-08 1.19456633e-08 7.52042316e-08 1.19595806e-08 7.53042316e-08 1.1946313e-08 7.54042316e-08 1.19589612e-08 7.55042316e-08 1.19469037e-08 7.56042316e-08 1.19583982e-08
+ 7.57042316e-08 1.19474406e-08 7.58042316e-08 1.19578862e-08 7.59042316e-08 1.19479288e-08 7.60042316e-08 1.19574207e-08 7.61042316e-08 1.19483725e-08 7.62042316e-08 1.19569974e-08 7.63042316e-08 1.19487758e-08 7.64042316e-08 1.19566131e-08
+ 7.65042316e-08 1.19491426e-08 7.66042316e-08 1.19562633e-08 7.67042316e-08 1.19494762e-08 7.68042316e-08 1.19559453e-08 7.69042316e-08 1.19497792e-08 7.70042316e-08 1.19556563e-08 7.71042316e-08 1.19500546e-08 7.72042316e-08 1.19553937e-08
+ 7.73042316e-08 1.19503053e-08 7.74042316e-08 1.1955155e-08 7.75042316e-08 1.19505328e-08 7.76042316e-08 1.19549377e-08 7.77042316e-08 1.19507396e-08 7.78042316e-08 1.19547406e-08 7.79042316e-08 1.19509277e-08 7.80042316e-08 1.1954561e-08
+ 7.81042316e-08 1.1951099e-08 7.82042316e-08 1.19543981e-08 7.83042316e-08 1.19512544e-08 7.84042316e-08 1.19542503e-08 7.85042316e-08 1.19513952e-08 7.86042316e-08 1.19541155e-08 7.87042316e-08 1.19515237e-08 7.88042316e-08 1.19539933e-08
+ 7.89042316e-08 1.19516399e-08 7.90042316e-08 1.19538824e-08 7.91042316e-08 1.19517458e-08 7.92042316e-08 1.19537817e-08 7.93042316e-08 1.19518415e-08 7.94042316e-08 1.19536904e-08 7.95042316e-08 1.19519286e-08 7.96042316e-08 1.19536075e-08
+ 7.97042316e-08 1.19520075e-08 7.98042316e-08 1.1953532e-08 7.99042316e-08 1.19520794e-08 8.00042316e-08 1.19534641e-08 8.01042316e-08 1.19521444e-08 8.02042316e-08 1.19534019e-08 8.03042316e-08 1.19522035e-08 8.04042316e-08 1.19533455e-08
+ 8.05042316e-08 1.19522574e-08 8.06042316e-08 1.19532938e-08 8.07042316e-08 1.19523063e-08 8.08042316e-08 1.19532477e-08 8.09042316e-08 1.19523502e-08 8.10042316e-08 1.19532053e-08 8.11042316e-08 1.1952391e-08 8.12042316e-08 1.19531671e-08
+ 8.13042316e-08 1.19524272e-08 8.14042316e-08 1.19531327e-08 8.15042316e-08 1.195246e-08 8.16042316e-08 1.19531013e-08 8.17042316e-08 1.19524899e-08 8.18042316e-08 1.19530723e-08 8.19042316e-08 1.19525173e-08 8.20042316e-08 1.19530465e-08
+ 8.21042316e-08 1.1952542e-08 8.22042316e-08 1.1953023e-08 8.23042316e-08 1.19525646e-08 8.24042316e-08 1.19530016e-08 8.25042316e-08 1.1952585e-08 8.26042316e-08 1.1952982e-08 8.27042316e-08 1.19526034e-08 8.28042316e-08 1.19529643e-08
+ 8.29042316e-08 1.19526203e-08 8.30042316e-08 1.19529483e-08 8.31042316e-08 1.1952636e-08 8.32042316e-08 1.19529336e-08 8.33042316e-08 1.19526497e-08 8.34042316e-08 1.19529203e-08 8.35042316e-08 1.19526625e-08 8.36042316e-08 1.19529083e-08
+ 8.37042316e-08 1.1952674e-08 8.38042316e-08 1.19528973e-08 8.39042316e-08 1.19526847e-08 8.40042316e-08 1.19528872e-08 8.41042316e-08 1.1952694e-08 8.42042316e-08 1.19528781e-08 8.43042316e-08 1.19527024e-08 8.44042316e-08 1.195287e-08
+ 8.45042316e-08 1.19527104e-08 8.46042316e-08 1.19528628e-08 8.47042316e-08 1.19527172e-08 8.48042316e-08 1.19528561e-08 8.49042316e-08 1.19527239e-08 8.50042316e-08 1.19528496e-08 8.51042316e-08 1.19527297e-08 8.52042316e-08 1.19528442e-08
+ 8.53042316e-08 1.19527353e-08 8.54042316e-08 1.1952839e-08 8.55042316e-08 1.19527398e-08 8.56042316e-08 1.19528344e-08 8.57042316e-08 1.19527441e-08 8.58042316e-08 1.19528302e-08 8.59042316e-08 1.19527483e-08 8.60042316e-08 1.19528265e-08
+ 8.61042316e-08 1.1952752e-08 8.62042316e-08 1.19528227e-08 8.63042316e-08 1.19527555e-08 8.64042316e-08 1.19528197e-08 8.65042316e-08 1.19527586e-08 8.66042316e-08 1.19528166e-08 8.67042316e-08 1.19527612e-08 8.68042316e-08 1.19528139e-08
+ 8.69042316e-08 1.19527637e-08 8.70042316e-08 1.19528119e-08 8.71042316e-08 1.1952766e-08 8.72042316e-08 1.19528096e-08 8.73042316e-08 1.1952768e-08 8.74042316e-08 1.19528077e-08 8.75042316e-08 1.195277e-08 8.76042316e-08 1.1952806e-08
+ 8.77042316e-08 1.19527715e-08 8.78042316e-08 1.19528044e-08 8.79042316e-08 1.19527731e-08 8.80042316e-08 1.19528028e-08 8.81042316e-08 1.19527745e-08 8.82042316e-08 1.19528013e-08 8.83042316e-08 1.19527758e-08 8.84042316e-08 1.19528002e-08
+ 8.85042316e-08 1.1952777e-08 8.86042316e-08 1.19527993e-08 8.87042316e-08 1.19527781e-08 8.88042316e-08 1.19527981e-08 8.89042316e-08 1.19527789e-08 8.90042316e-08 1.19527973e-08 8.91042316e-08 1.19527795e-08 8.92042316e-08 1.19527964e-08
+ 8.93042316e-08 1.19527807e-08 8.94042316e-08 1.19527957e-08 8.95042316e-08 1.19527812e-08 8.96042316e-08 1.19527949e-08 8.97042316e-08 1.19527822e-08 8.98042316e-08 1.19527941e-08 8.99042316e-08 1.19527826e-08 9.00042316e-08 1.19527935e-08
+ 9.01042316e-08 1.19527831e-08 9.02042316e-08 1.19527931e-08 9.03042316e-08 1.19527837e-08 9.04042316e-08 1.19527928e-08 9.05042316e-08 1.1952784e-08 9.06042316e-08 1.19527922e-08 9.07042316e-08 1.19527846e-08 9.08042316e-08 1.1952792e-08
+ 9.09042316e-08 1.19527847e-08 9.10042316e-08 1.19527916e-08 9.11042316e-08 1.1952785e-08 9.12042316e-08 1.19527916e-08 9.13042316e-08 1.19527853e-08 9.14042316e-08 1.19527912e-08 9.15042316e-08 1.19527858e-08 9.16042316e-08 1.1952791e-08
+ 9.17042316e-08 1.19527859e-08 9.18042316e-08 1.19527906e-08 9.19042316e-08 1.19527861e-08 9.20042316e-08 1.19527903e-08 9.21042316e-08 1.19527864e-08 9.22042316e-08 1.19527902e-08 9.23042316e-08 1.19527866e-08 9.24042316e-08 1.19527901e-08
+ 9.25042316e-08 1.19527868e-08 9.26042316e-08 1.19527899e-08 9.27042316e-08 1.19527868e-08 9.28042316e-08 1.19527898e-08 9.29042316e-08 1.19527868e-08 9.30042316e-08 1.19527898e-08 9.31042316e-08 1.1952787e-08 9.32042316e-08 1.19527895e-08
+ 9.33042316e-08 1.19527869e-08 9.34042316e-08 1.19527897e-08 9.35042316e-08 1.1952787e-08 9.36042316e-08 1.19527897e-08 9.37042316e-08 1.19527871e-08 9.38042316e-08 1.19527895e-08 9.39042316e-08 1.19527873e-08 9.40042316e-08 1.19527893e-08
+ 9.41042316e-08 1.19527875e-08 9.42042316e-08 1.1952789e-08 9.43042316e-08 1.19527874e-08 9.44042316e-08 1.1952789e-08 9.45042316e-08 1.19527875e-08 9.46042316e-08 1.19527891e-08 9.47042316e-08 1.19527877e-08 9.48042316e-08 1.19527888e-08
+ 9.49042316e-08 1.19527878e-08 9.50042316e-08 1.19527886e-08 9.51042316e-08 1.19527878e-08 9.52042316e-08 1.19527887e-08 9.53042316e-08 1.19527878e-08 9.54042316e-08 1.19527888e-08 9.55042316e-08 1.19527877e-08 9.56042316e-08 1.19527889e-08
+ 9.57042316e-08 1.1952788e-08 9.58042316e-08 1.19527888e-08 9.59042316e-08 1.19527878e-08 9.60042316e-08 1.19527885e-08 9.61042316e-08 1.19527878e-08 9.62042316e-08 1.19527885e-08 9.63042316e-08 1.19527878e-08 9.64042316e-08 1.19527886e-08
+ 9.65042316e-08 1.19527882e-08 9.66042316e-08 1.19527886e-08 9.67042316e-08 1.19527881e-08 9.68042316e-08 1.19527887e-08 9.69042316e-08 1.19527881e-08 9.70042316e-08 1.19527888e-08 9.71042316e-08 1.19527882e-08 9.72042316e-08 1.19527885e-08
+ 9.73042316e-08 1.19527883e-08 9.74042316e-08 1.19527884e-08 9.75042316e-08 1.19527881e-08 9.76042316e-08 1.19527882e-08 9.77042316e-08 1.1952788e-08 9.78042316e-08 1.19527883e-08 9.79042316e-08 1.1952788e-08 9.80042316e-08 1.19527883e-08
+ 9.81042316e-08 1.1952788e-08 9.82042316e-08 1.19527883e-08 9.83042316e-08 1.1952788e-08 9.84042316e-08 1.19527883e-08 9.85042316e-08 1.19527879e-08 9.86042316e-08 1.19527884e-08 9.87042316e-08 1.19527879e-08 9.88042316e-08 1.19527884e-08
+ 9.89042316e-08 1.19527879e-08 9.90042316e-08 1.19527884e-08 9.91042316e-08 1.19527879e-08 9.92042316e-08 1.19527885e-08 9.93042316e-08 1.19527879e-08 9.94042316e-08 1.19527884e-08 9.95042316e-08 1.19527879e-08 9.96042316e-08 1.19527885e-08
+ 9.97042316e-08 1.19527878e-08 9.98042316e-08 1.19527885e-08 9.99042316e-08 1.1952788e-08 1e-07 1.19527887e-08 1.0001e-07 1.19843157e-08 1.0003e-07 1.17984604e-08 1.0007e-07 1.2192678e-08 1.0015e-07 1.16828425e-08
+ 1.0025e-07 1.22306964e-08 1.0035e-07 1.16831308e-08 1.0045e-07 1.21985944e-08 1.0055e-07 1.17500971e-08 1.0065e-07 1.18572505e-08 1.0075e-07 2.60724813e-08 1.0085e-07 -6.68242726e-07 1.00932051e-07 4.41896813e-06
+ 1.01e-07 -1.00694179e-05 1.01008488e-07 -1.02957209e-05 1.01025463e-07 4.64439514e-06 1.01059414e-07 6.17767808e-06 1.0109062e-07 3.02645003e-06 1.0114347e-07 -2.66952664e-07 1.01199151e-07 8.0803544e-06 1.01299151e-07 -3.08581739e-05
+ 1.01399151e-07 0.000140233009 1.01499151e-07 -0.000220926504 1.01599151e-07 0.000209325087 1.01699151e-07 -0.000302115401 1.01799151e-07 0.000382343756 1.01893117e-07 -0.000382660074 1.01993117e-07 0.000390002872 1.02093117e-07 -0.00038322251
+ 1.02193117e-07 0.000370033687 1.02293117e-07 -0.000351833758 1.02393117e-07 0.000330885424 1.02493117e-07 -0.000308234189 1.02593117e-07 0.000285448498 1.02693117e-07 -0.000262835121 1.02793117e-07 0.000241355801 1.02893117e-07 -0.000220866106
+ 1.02993117e-07 0.000201938945 1.03093117e-07 -0.000184229611 1.03193117e-07 0.000168099169 1.03293117e-07 -0.000153146898 1.03393117e-07 0.000139624338 1.03493117e-07 -0.000127141006 1.03593117e-07 0.000115892869 1.03693117e-07 -0.000105523311
+ 1.03793117e-07 9.61985944e-05 1.03893117e-07 -8.76011855e-05 1.03993117e-07 7.98800579e-05 1.04093117e-07 -7.2754336e-05 1.04193117e-07 6.63618384e-05 1.04293117e-07 -6.04535358e-05 1.04393117e-07 5.51593269e-05 1.04493117e-07 -5.02569369e-05
+ 1.04593117e-07 4.58702337e-05 1.04693117e-07 -4.17990937e-05 1.04793117e-07 3.81625873e-05 1.04893117e-07 -3.47788243e-05 1.04993117e-07 3.17629641e-05 1.05093117e-07 -2.89481014e-05 1.05193117e-07 2.64461661e-05 1.05293117e-07 -2.41025714e-05
+ 1.05393117e-07 2.20265626e-05 1.05493117e-07 -2.00736917e-05 1.05593117e-07 1.83509654e-05 1.05693117e-07 -1.67222914e-05 1.05793117e-07 1.52928075e-05 1.05893117e-07 -1.39333182e-05 1.05993117e-07 1.27473992e-05 1.06093117e-07 -1.16115549e-05
+ 1.06193117e-07 1.06280554e-05 1.06293117e-07 -9.67812186e-06 1.06393117e-07 8.86293251e-06 1.06493117e-07 -8.06761573e-06 1.06593117e-07 7.39243728e-06 1.06693117e-07 -6.68331516e-06 1.06793117e-07 6.17335834e-06 1.06893117e-07 -5.57478631e-06
+ 1.06993117e-07 5.15354516e-06 1.07093117e-07 -4.65033415e-06 1.07193117e-07 4.30299237e-06 1.07293117e-07 -3.87926558e-06 1.07393117e-07 3.59349993e-06 1.07493117e-07 -3.23603174e-06 1.07593117e-07 3.00158461e-06 1.07693117e-07 -2.69935978e-06
+ 1.07793117e-07 2.50769152e-06 1.07893117e-07 -2.25153441e-06 1.07993117e-07 2.1089765e-06 1.08093117e-07 -1.87566961e-06 1.08193117e-07 1.76168627e-06 1.08293117e-07 -1.56308438e-06 1.08393117e-07 1.47197494e-06 1.08493117e-07 -1.30232738e-06
+ 1.08593117e-07 1.23028425e-06 1.08693117e-07 -1.08478071e-06 1.08793117e-07 1.02863478e-06 1.08893117e-07 -9.03267173e-07 1.08993117e-07 8.60377678e-07 1.09093117e-07 -7.51805599e-07 1.09193117e-07 7.19972287e-07 1.09293117e-07 -6.25411135e-07
+ 1.09393117e-07 6.02800373e-07 1.09493117e-07 -5.19928465e-07 1.09593117e-07 5.05011231e-07 1.09693117e-07 -4.31892402e-07 1.09793117e-07 4.23394e-07 1.09893117e-07 -3.58413241e-07 1.09993117e-07 3.55270146e-07 1.10093117e-07 -2.97080227e-07
+ 1.10193117e-07 2.98405669e-07 1.10293117e-07 -2.45882941e-07 1.10393117e-07 2.50937343e-07 1.10493117e-07 -2.0314448e-07 1.10593117e-07 2.1131093e-07 1.10693117e-07 -1.67465823e-07 1.10793117e-07 1.7822958e-07 1.10893117e-07 -1.3767959e-07
+ 1.10993117e-07 1.50611157e-07 1.11093117e-07 -1.12811646e-07 1.11193117e-07 1.27552605e-07 1.11293117e-07 -9.20490655e-08 1.11393117e-07 1.08300333e-07 1.11493117e-07 -7.47149043e-08 1.11593117e-07 9.22283551e-08 1.11693117e-07 -6.02462155e-08
+ 1.11793117e-07 7.88150193e-08 1.11893117e-07 -4.81705203e-08 1.11993117e-07 6.76201229e-08 1.12093117e-07 -3.80921457e-08 1.12193117e-07 5.8276667e-08 1.12293117e-07 -2.96803156e-08 1.12393117e-07 5.04780957e-08 1.12493117e-07 -2.26592329e-08
+ 1.12593117e-07 4.39688022e-08 1.12693117e-07 -1.67988287e-08 1.12793117e-07 3.85355268e-08 1.12893117e-07 -1.18935464e-08 1.12993117e-07 3.39879655e-08 1.13093117e-07 -7.81334442e-09 1.13193117e-07 3.02048422e-08 1.13293117e-07 -4.407159e-09
+ 1.13393117e-07 2.70468237e-08 1.13493117e-07 -1.56378385e-09 1.13593117e-07 2.44105963e-08 1.13693117e-07 8.09806638e-10 1.13793117e-07 2.22204477e-08 1.13893117e-07 2.78229173e-09 1.13993117e-07 2.04173205e-08 1.14093117e-07 4.40704434e-09
+ 1.14193117e-07 1.89320684e-08 1.14293117e-07 5.74538023e-09 1.14393117e-07 1.77086319e-08 1.14493117e-07 6.84780377e-09 1.14593117e-07 1.67008505e-08 1.14693117e-07 7.75590589e-09 1.14793117e-07 1.58707073e-08 1.14893117e-07 8.50394116e-09
+ 1.14993117e-07 1.50886834e-08 1.15093117e-07 9.10616932e-09 1.15193117e-07 1.45368225e-08 1.15293117e-07 9.60716226e-09 1.15393117e-07 1.40819625e-08 1.15493117e-07 1.00201277e-08 1.15593117e-07 1.37070384e-08 1.15693117e-07 1.03605111e-08
+ 1.15793117e-07 1.33980156e-08 1.15893117e-07 1.06410608e-08 1.15993117e-07 1.3143318e-08 1.16093117e-07 1.08722873e-08 1.16193117e-07 1.29334015e-08 1.16293117e-07 1.10628563e-08 1.16393117e-07 1.27603986e-08 1.16493117e-07 1.12199106e-08
+ 1.16593117e-07 1.26178241e-08 1.16693117e-07 1.13493387e-08 1.16793117e-07 1.25003314e-08 1.16893117e-07 1.14559949e-08 1.16993117e-07 1.24035135e-08 1.17093117e-07 1.15438805e-08 1.17193117e-07 1.23237376e-08 1.17293117e-07 1.16162935e-08
+ 1.17393117e-07 1.22580092e-08 1.17493117e-07 1.16759534e-08 1.17593117e-07 1.22038587e-08 1.17693117e-07 1.17251016e-08 1.17793117e-07 1.21592517e-08 1.17893117e-07 1.17655863e-08 1.17993117e-07 1.21225097e-08 1.18093117e-07 1.17989305e-08
+ 1.18193117e-07 1.20922499e-08 1.18293117e-07 1.18263899e-08 1.18393117e-07 1.20673331e-08 1.18493117e-07 1.18489988e-08 1.18593117e-07 1.20468191e-08 1.18693117e-07 1.18676109e-08 1.18793117e-07 1.20299337e-08 1.18893117e-07 1.1882929e-08
+ 1.18993117e-07 1.20160384e-08 1.19093117e-07 1.18955329e-08 1.19193117e-07 1.20046068e-08 1.19293117e-07 1.19058997e-08 1.19393117e-07 1.19952064e-08 1.19493117e-07 1.19144241e-08 1.19593117e-07 1.19874772e-08 1.19693117e-07 1.19214318e-08
+ 1.19793117e-07 1.19811245e-08 1.19893117e-07 1.19271895e-08 1.19993117e-07 1.19759066e-08 1.20093117e-07 1.19319174e-08 1.20193117e-07 1.19716233e-08 1.20293117e-07 1.19357973e-08 1.20393117e-07 1.19681095e-08 1.20493117e-07 1.19389791e-08
+ 1.20593117e-07 1.19652286e-08 1.20693117e-07 1.19415871e-08 1.20793117e-07 1.19628679e-08 1.20893117e-07 1.19437232e-08 1.20993117e-07 1.1960936e-08 1.21093117e-07 1.19454703e-08 1.21193117e-07 1.19593564e-08 1.21293117e-07 1.19468978e-08
+ 1.21393117e-07 1.19580661e-08 1.21493117e-07 1.19480633e-08 1.21593117e-07 1.1957014e-08 1.21693117e-07 1.19490133e-08 1.21793117e-07 1.19561572e-08 1.21893117e-07 1.19497862e-08 1.21993117e-07 1.19554599e-08 1.22093117e-07 1.19504143e-08
+ 1.22193117e-07 1.19548942e-08 1.22293117e-07 1.19509235e-08 1.22393117e-07 1.1954436e-08 1.22493117e-07 1.19513358e-08 1.22593117e-07 1.19540655e-08 1.22693117e-07 1.19516682e-08 1.22793117e-07 1.1953767e-08 1.22893117e-07 1.1951936e-08
+ 1.22993117e-07 1.19535271e-08 1.23093117e-07 1.19521507e-08 1.23193117e-07 1.19533349e-08 1.23293117e-07 1.19523225e-08 1.23393117e-07 1.19531821e-08 1.23493117e-07 1.19524589e-08 1.23593117e-07 1.19530608e-08 1.23693117e-07 1.19525667e-08
+ 1.23793117e-07 1.1952965e-08 1.23893117e-07 1.19526511e-08 1.23993117e-07 1.19528906e-08 1.24093117e-07 1.19527166e-08 1.24193117e-07 1.19528329e-08 1.24293117e-07 1.19527673e-08 1.24393117e-07 1.19527886e-08 1.24493117e-07 1.1952806e-08
+ 1.24593117e-07 1.19527553e-08 1.24693117e-07 1.19528344e-08 1.24793117e-07 1.19527306e-08 1.24893117e-07 1.19528555e-08 1.24993117e-07 1.1952713e-08 1.25093117e-07 1.195287e-08 1.25193117e-07 1.19527006e-08 1.25293117e-07 1.19528804e-08
+ 1.25393117e-07 1.19526928e-08 1.25493117e-07 1.19528863e-08 1.25593117e-07 1.19526884e-08 1.25693117e-07 1.19528893e-08 1.25793117e-07 1.19526865e-08 1.25893117e-07 1.19528901e-08 1.25993117e-07 1.19526864e-08 1.26093117e-07 1.19528897e-08
+ 1.26193117e-07 1.19526881e-08 1.26293117e-07 1.1952887e-08 1.26393117e-07 1.19526909e-08 1.26493117e-07 1.19528837e-08 1.26593117e-07 1.19526944e-08 1.26693117e-07 1.195288e-08 1.26793117e-07 1.19526989e-08 1.26893117e-07 1.19528756e-08
+ 1.26993117e-07 1.19527034e-08 1.27093117e-07 1.19528711e-08 1.27193117e-07 1.19527079e-08 1.27293117e-07 1.19528664e-08 1.27393117e-07 1.19527124e-08 1.27493117e-07 1.19528618e-08 1.27593117e-07 1.19527173e-08 1.27693117e-07 1.1952857e-08
+ 1.27793117e-07 1.19527221e-08 1.27893117e-07 1.19528522e-08 1.27993117e-07 1.19527266e-08 1.28093117e-07 1.19528479e-08 1.28193117e-07 1.19527309e-08 1.28293117e-07 1.19528437e-08 1.28393117e-07 1.19527353e-08 1.28493117e-07 1.19528394e-08
+ 1.28593117e-07 1.19527391e-08 1.28693117e-07 1.19528357e-08 1.28793117e-07 1.19527425e-08 1.28893117e-07 1.19528323e-08 1.28993117e-07 1.19527461e-08 1.29093117e-07 1.19528289e-08 1.29193117e-07 1.19527496e-08 1.29293117e-07 1.19528256e-08
+ 1.29393117e-07 1.19527523e-08 1.29493117e-07 1.19528228e-08 1.29593117e-07 1.19527553e-08 1.29693117e-07 1.195282e-08 1.29793117e-07 1.19527582e-08 1.29893117e-07 1.19528173e-08 1.29993117e-07 1.19527604e-08 1.30093117e-07 1.19528149e-08
+ 1.30193117e-07 1.19527625e-08 1.30293117e-07 1.19528127e-08 1.30393117e-07 1.19527648e-08 1.30493117e-07 1.19528107e-08 1.30593117e-07 1.19527666e-08 1.30693117e-07 1.19528089e-08 1.30793117e-07 1.19527683e-08 1.30893117e-07 1.19528072e-08
+ 1.30993117e-07 1.19527702e-08 1.31093117e-07 1.19528055e-08 1.31193117e-07 1.19527717e-08 1.31293117e-07 1.19528039e-08 1.31393117e-07 1.19527733e-08 1.31493117e-07 1.19528025e-08 1.31593117e-07 1.19527745e-08 1.31693117e-07 1.19528012e-08
+ 1.31793117e-07 1.1952776e-08 1.31893117e-07 1.19528001e-08 1.31993117e-07 1.19527769e-08 1.32093117e-07 1.19527992e-08 1.32193117e-07 1.19527779e-08 1.32293117e-07 1.19527984e-08 1.32393117e-07 1.19527786e-08 1.32493117e-07 1.19527974e-08
+ 1.32593117e-07 1.19527793e-08 1.32693117e-07 1.19527967e-08 1.32793117e-07 1.19527803e-08 1.32893117e-07 1.19527958e-08 1.32993117e-07 1.19527811e-08 1.33093117e-07 1.19527952e-08 1.33193117e-07 1.19527817e-08 1.33293117e-07 1.19527945e-08
+ 1.33393117e-07 1.19527823e-08 1.33493117e-07 1.19527942e-08 1.33593117e-07 1.19527827e-08 1.33693117e-07 1.19527935e-08 1.33793117e-07 1.19527834e-08 1.33893117e-07 1.19527932e-08 1.33993117e-07 1.19527837e-08 1.34093117e-07 1.19527929e-08
+ 1.34193117e-07 1.1952784e-08 1.34293117e-07 1.19527924e-08 1.34393117e-07 1.19527844e-08 1.34493117e-07 1.19527921e-08 1.34593117e-07 1.19527845e-08 1.34693117e-07 1.19527918e-08 1.34793117e-07 1.19527847e-08 1.34893117e-07 1.19527914e-08
+ 1.34993117e-07 1.19527853e-08 1.35093117e-07 1.19527915e-08 1.35193117e-07 1.19527854e-08 1.35293117e-07 1.19527911e-08 1.35393117e-07 1.19527857e-08 1.35493117e-07 1.19527909e-08 1.35593117e-07 1.19527859e-08 1.35693117e-07 1.19527906e-08
+ 1.35793117e-07 1.19527862e-08 1.35893117e-07 1.19527905e-08 1.35993117e-07 1.19527865e-08 1.36093117e-07 1.19527902e-08 1.36193117e-07 1.19527864e-08 1.36293117e-07 1.19527902e-08 1.36393117e-07 1.19527868e-08 1.36493117e-07 1.19527897e-08
+ 1.36593117e-07 1.19527868e-08 1.36693117e-07 1.19527898e-08 1.36793117e-07 1.19527869e-08 1.36893117e-07 1.19527898e-08 1.36993117e-07 1.19527869e-08 1.37093117e-07 1.19527899e-08 1.37193117e-07 1.1952787e-08 1.37293117e-07 1.19527896e-08
+ 1.37393117e-07 1.19527871e-08 1.37493117e-07 1.19527896e-08 1.37593117e-07 1.19527872e-08 1.37693117e-07 1.19527893e-08 1.37793117e-07 1.19527872e-08 1.37893117e-07 1.19527892e-08 1.37993117e-07 1.19527872e-08 1.38093117e-07 1.19527892e-08
+ 1.38193117e-07 1.19527872e-08 1.38293117e-07 1.19527892e-08 1.38393117e-07 1.19527872e-08 1.38493117e-07 1.19527893e-08 1.38593117e-07 1.19527872e-08 1.38693117e-07 1.19527891e-08 1.38793117e-07 1.19527873e-08 1.38893117e-07 1.19527893e-08
+ 1.38993117e-07 1.19527876e-08 1.39093117e-07 1.19527891e-08 1.39193117e-07 1.19527876e-08 1.39293117e-07 1.1952789e-08 1.39393117e-07 1.19527876e-08 1.39493117e-07 1.19527889e-08 1.39593117e-07 1.19527877e-08 1.39693117e-07 1.19527891e-08
+ 1.39793117e-07 1.19527876e-08 1.39893117e-07 1.19527891e-08 1.39993117e-07 1.19527876e-08 1.40093117e-07 1.19527889e-08 1.40193117e-07 1.19527878e-08 1.40293117e-07 1.19527889e-08 1.40393117e-07 1.1952788e-08 1.40493117e-07 1.19527889e-08
+ 1.40593117e-07 1.19527878e-08 1.40693117e-07 1.19527888e-08 1.40793117e-07 1.19527878e-08 1.40893117e-07 1.1952789e-08 1.40993117e-07 1.19527879e-08 1.41093117e-07 1.1952789e-08 1.41193117e-07 1.19527879e-08 1.41293117e-07 1.1952789e-08
+ 1.41393117e-07 1.19527878e-08 1.41493117e-07 1.1952789e-08 1.41593117e-07 1.19527879e-08 1.41693117e-07 1.1952789e-08 1.41793117e-07 1.19527878e-08 1.41893117e-07 1.1952789e-08 1.41993117e-07 1.19527879e-08 1.42093117e-07 1.19527889e-08
+ 1.42193117e-07 1.19527877e-08 1.42293117e-07 1.19527887e-08 1.42393117e-07 1.1952788e-08 1.42493117e-07 1.19527888e-08 1.42593117e-07 1.1952788e-08 1.42693117e-07 1.19527888e-08 1.42793117e-07 1.1952788e-08 1.42893117e-07 1.19527889e-08
+ 1.42993117e-07 1.19527879e-08 1.43093117e-07 1.19527888e-08 1.43193117e-07 1.19527878e-08 1.43293117e-07 1.19527886e-08 1.43393117e-07 1.19527883e-08 1.43493117e-07 1.19527885e-08 1.43593117e-07 1.19527879e-08 1.43693117e-07 1.19527883e-08
+ 1.43793117e-07 1.1952788e-08 1.43893117e-07 1.19527883e-08 1.43993117e-07 1.1952788e-08 1.44093117e-07 1.19527881e-08 1.44193117e-07 1.1952788e-08 1.44293117e-07 1.19527883e-08 1.44393117e-07 1.19527881e-08 1.44493117e-07 1.19527882e-08
+ 1.44593117e-07 1.19527881e-08 1.44693117e-07 1.19527882e-08 1.44793117e-07 1.19527882e-08 1.44893117e-07 1.19527883e-08 1.44993117e-07 1.19527879e-08 1.45093117e-07 1.19527882e-08 1.45193117e-07 1.1952788e-08 1.45293117e-07 1.19527883e-08
+ 1.45393117e-07 1.19527881e-08 1.45493117e-07 1.19527882e-08 1.45593117e-07 1.19527881e-08 1.45693117e-07 1.19527882e-08 1.45793117e-07 1.19527881e-08 1.45893117e-07 1.19527882e-08 1.45993117e-07 1.19527881e-08 1.46093117e-07 1.19527881e-08
+ 1.46193117e-07 1.19527883e-08 1.46293117e-07 1.19527881e-08 1.46393117e-07 1.19527883e-08 1.46493117e-07 1.19527881e-08 1.46593117e-07 1.1952788e-08 1.46693117e-07 1.19527883e-08 1.46793117e-07 1.19527881e-08 1.46893117e-07 1.19527883e-08
+ 1.46993117e-07 1.1952788e-08 1.47093117e-07 1.19527882e-08 1.47193117e-07 1.19527881e-08 1.47293117e-07 1.19527883e-08 1.47393117e-07 1.1952788e-08 1.47493117e-07 1.19527882e-08 1.47593117e-07 1.19527881e-08 1.47693117e-07 1.19527883e-08
+ 1.47793117e-07 1.1952788e-08 1.47893117e-07 1.19527882e-08 1.47993117e-07 1.19527881e-08 1.48093117e-07 1.19527883e-08 1.48193117e-07 1.1952788e-08 1.48293117e-07 1.19527882e-08 1.48393117e-07 1.19527881e-08 1.48493117e-07 1.19527883e-08
+ 1.48593117e-07 1.1952788e-08 1.48693117e-07 1.19527882e-08 1.48793117e-07 1.19527881e-08 1.48893117e-07 1.19527882e-08 1.48993117e-07 1.1952788e-08 1.49093117e-07 1.19527883e-08 1.49193117e-07 1.19527881e-08 1.49293117e-07 1.19527882e-08
+ 1.49393117e-07 1.1952788e-08 1.49493117e-07 1.19527884e-08 1.49593117e-07 1.1952788e-08 1.49693117e-07 1.19527883e-08 1.49793117e-07 1.19527881e-08 1.49893117e-07 1.19527881e-08 1.49993117e-07 1.19527881e-08 1.50093117e-07 1.19527882e-08
+ 1.50193117e-07 1.19527881e-08 1.50293117e-07 1.19527883e-08 1.50393117e-07 1.19527881e-08 1.50493117e-07 1.19527883e-08 1.50593117e-07 1.1952788e-08 1.50693117e-07 1.19527883e-08 1.50793117e-07 1.19527881e-08 1.50893117e-07 1.19527883e-08
+ 1.50993117e-07 1.1952788e-08 1.51e-07 1.19527885e-08 1.5101e-07 1.19399425e-08 1.5103e-07 1.2015012e-08 1.5107e-07 1.18559373e-08 1.5115e-07 1.2062103e-08 1.5125e-07 1.18410984e-08 1.5135e-07 1.20574879e-08
+ 1.5145e-07 1.18638218e-08 1.5155e-07 1.20197038e-08 1.5165e-07 1.19101577e-08 1.5175e-07 1.19686133e-08 1.5185e-07 1.19674861e-08 1.51930828e-07 1.83418271e-07 1.52e-07 1.06002511e-07 1.52008608e-07 -6.35218177e-06
+ 1.52025825e-07 -6.40058772e-06 1.52060258e-07 9.75152889e-06 1.52106188e-07 5.28436065e-06 1.52150118e-07 -1.51923821e-05 1.5219811e-07 6.42631694e-06 1.52255501e-07 9.57203275e-07 1.52312176e-07 -1.57312897e-06 1.52404431e-07 1.13651066e-06
+ 1.52490774e-07 -1.00481012e-06 1.52590774e-07 9.71177181e-07 1.52690774e-07 -8.68538702e-07 1.52790774e-07 8.16800246e-07 1.52890774e-07 -7.24280335e-07 1.52990774e-07 6.88959109e-07 1.53090774e-07 -6.14045776e-07 1.53190774e-07 5.94780994e-07
+ 1.53290774e-07 -5.33636397e-07 1.53390774e-07 5.25524356e-07 1.53490774e-07 -4.73280576e-07 1.53590774e-07 4.72031482e-07 1.53690774e-07 -4.25080802e-07 1.53790774e-07 4.27831273e-07 1.53890774e-07 -3.83949754e-07 1.53990774e-07 3.89044558e-07
+ 1.54090774e-07 -3.47015132e-07 1.54190774e-07 3.53600162e-07 1.54290774e-07 -3.1283798e-07 1.54390774e-07 3.20535389e-07 1.54490774e-07 -2.8080758e-07 1.54590774e-07 2.89489066e-07 1.54690774e-07 -2.50736593e-07 1.54790774e-07 2.60387935e-07
+ 1.54890774e-07 -2.22622727e-07 1.54990774e-07 2.33268483e-07 1.55090774e-07 -1.96518922e-07 1.55190774e-07 2.08184555e-07 1.55290774e-07 -1.72469417e-07 1.55390774e-07 1.85164419e-07 1.55490774e-07 -1.5048341e-07 1.55590774e-07 1.64197736e-07
+ 1.55690774e-07 -1.30531136e-07 1.55790774e-07 1.45236105e-07 1.55890774e-07 -1.12546679e-07 1.55990774e-07 1.28198009e-07 1.56090774e-07 -9.64348403e-08 1.56190774e-07 1.12976722e-07 1.56290774e-07 -8.20793923e-08 1.56390774e-07 9.94488437e-08
+ 1.56490774e-07 -6.93518937e-08 1.56590774e-07 8.74824824e-08 1.56690774e-07 -5.81181588e-08 1.56790774e-07 7.69424794e-08 1.56890774e-07 -4.82432685e-08 1.56990774e-07 6.76957126e-08 1.57090774e-07 -3.95973242e-08 1.57190774e-07 5.96159857e-08
+ 1.57290774e-07 -3.20580606e-08 1.57390774e-07 5.25831339e-08 1.57490774e-07 -2.55059897e-08 1.57590774e-07 4.64804555e-08 1.57690774e-07 -1.98288805e-08 1.57790774e-07 4.12001345e-08 1.57890774e-07 -1.49233718e-08 1.57990774e-07 3.6643288e-08
+ 1.58090774e-07 -1.06953085e-08 1.58190774e-07 3.27206463e-08 1.58290774e-07 -7.06022138e-09 1.58390774e-07 2.93522183e-08 1.58490774e-07 -3.94248906e-09 1.58590774e-07 2.6466716e-08 1.58690774e-07 -1.27504032e-09 1.58790774e-07 2.40009079e-08
+ 1.58890774e-07 9.95289573e-10 1.58990774e-07 2.19106553e-08 1.59090774e-07 2.91105623e-09 1.59190774e-07 2.01553628e-08 1.59290774e-07 4.51844337e-09 1.59390774e-07 1.86842277e-08 1.59490774e-07 5.864113e-09 1.59590774e-07 1.7454049e-08
+ 1.59690774e-07 6.98801472e-09 1.59790774e-07 1.64279171e-08 1.59890774e-07 7.92425447e-09 1.59990774e-07 1.55742663e-08 1.60090774e-07 8.70207323e-09 1.60190774e-07 1.48660349e-08 1.60290774e-07 9.34648151e-09 1.60390774e-07 1.42801325e-08
+ 1.60490774e-07 9.87878085e-09 1.60590774e-07 1.3796919e-08 1.60690774e-07 1.03170683e-08 1.60790774e-07 1.33997285e-08 1.60890774e-07 1.06766847e-08 1.60990774e-07 1.3074447e-08 1.61090774e-07 1.09706078e-08 1.61190774e-07 1.2809147e-08
+ 1.61290774e-07 1.1209796e-08 1.61390774e-07 1.25937661e-08 1.61490774e-07 1.14034843e-08 1.61590774e-07 1.24198311e-08 1.61690774e-07 1.15594432e-08 1.61790774e-07 1.22802219e-08 1.61890774e-07 1.16841978e-08 1.61990774e-07 1.21689479e-08
+ 1.62090774e-07 1.17832445e-08 1.62190774e-07 1.20809862e-08 1.62290774e-07 1.1861163e-08 1.62390774e-07 1.20121623e-08 1.62490774e-07 1.19217604e-08 1.62590774e-07 1.19589891e-08 1.62690774e-07 1.19682517e-08 1.62790774e-07 1.19184985e-08
+ 1.62890774e-07 1.2003359e-08 1.62990774e-07 1.188822e-08 1.63090774e-07 1.20293076e-08 1.63190774e-07 1.18661521e-08 1.63290774e-07 1.20479006e-08 1.63390774e-07 1.1850666e-08 1.63490774e-07 1.20606126e-08 1.63590774e-07 1.18404268e-08
+ 1.63690774e-07 1.20686533e-08 1.63790774e-07 1.18343362e-08 1.63890774e-07 1.20729633e-08 1.63990774e-07 1.18315274e-08 1.64090774e-07 1.20748436e-08 1.64190774e-07 1.18303351e-08 1.64290774e-07 1.20749986e-08 1.64390774e-07 1.18314627e-08
+ 1.64490774e-07 1.20727056e-08 1.64590774e-07 1.18346066e-08 1.64690774e-07 1.20689997e-08 1.64790774e-07 1.18387731e-08 1.64890774e-07 1.20644194e-08 1.64990774e-07 1.18436918e-08 1.65090774e-07 1.20592334e-08 1.65190774e-07 1.18490817e-08
+ 1.65290774e-07 1.20536923e-08 1.65390774e-07 1.18547565e-08 1.65490774e-07 1.20478497e-08 1.65590774e-07 1.18607562e-08 1.65690774e-07 1.20418228e-08 1.65790774e-07 1.18666814e-08 1.65890774e-07 1.20360293e-08 1.65990774e-07 1.18723594e-08
+ 1.66090774e-07 1.20304547e-08 1.66190774e-07 1.18778331e-08 1.66290774e-07 1.20250876e-08 1.66390774e-07 1.18830881e-08 1.66490774e-07 1.20199485e-08 1.66590774e-07 1.18881072e-08 1.66690774e-07 1.2015053e-08 1.66790774e-07 1.18928766e-08
+ 1.66890774e-07 1.20104109e-08 1.66990774e-07 1.18973895e-08 1.67090774e-07 1.20060287e-08 1.67190774e-07 1.190164e-08 1.67290774e-07 1.20019106e-08 1.67390774e-07 1.19056273e-08 1.67490774e-07 1.1998053e-08 1.67590774e-07 1.19093543e-08
+ 1.67690774e-07 1.19944559e-08 1.67790774e-07 1.1912825e-08 1.67890774e-07 1.19911087e-08 1.67990774e-07 1.19160522e-08 1.68090774e-07 1.19879979e-08 1.68190774e-07 1.19190487e-08 1.68290774e-07 1.19851126e-08 1.68390774e-07 1.19218422e-08
+ 1.68490774e-07 1.19823897e-08 1.68590774e-07 1.1924464e-08 1.68690774e-07 1.19799095e-08 1.68790774e-07 1.19268165e-08 1.68890774e-07 1.19776573e-08 1.68990774e-07 1.19289794e-08 1.69090774e-07 1.19755767e-08 1.69190774e-07 1.1930985e-08
+ 1.69290774e-07 1.19736411e-08 1.69390774e-07 1.19328468e-08 1.69490774e-07 1.19718586e-08 1.69590774e-07 1.19345518e-08 1.69690774e-07 1.19702252e-08 1.69790774e-07 1.19361179e-08 1.69890774e-07 1.19687256e-08 1.69990774e-07 1.19375515e-08
+ 1.70090774e-07 1.19673548e-08 1.70190774e-07 1.19388629e-08 1.70290774e-07 1.19660999e-08 1.70390774e-07 1.19400645e-08 1.70490774e-07 1.19649493e-08 1.70590774e-07 1.19411661e-08 1.70690774e-07 1.19638948e-08 1.70790774e-07 1.19421753e-08
+ 1.70890774e-07 1.19629286e-08 1.70990774e-07 1.19431002e-08 1.71090774e-07 1.1962044e-08 1.71190774e-07 1.19439458e-08 1.71290774e-07 1.1961235e-08 1.71390774e-07 1.19447196e-08 1.71490774e-07 1.19604953e-08 1.71590774e-07 1.19454269e-08
+ 1.71690774e-07 1.19598197e-08 1.71790774e-07 1.19460721e-08 1.71890774e-07 1.19592031e-08 1.71990774e-07 1.19466613e-08 1.72090774e-07 1.19586405e-08 1.72190774e-07 1.19471981e-08 1.72290774e-07 1.19581276e-08 1.72390774e-07 1.19476889e-08
+ 1.72490774e-07 1.19576588e-08 1.72590774e-07 1.19481366e-08 1.72690774e-07 1.19572314e-08 1.72790774e-07 1.19485446e-08 1.72890774e-07 1.19568415e-08 1.72990774e-07 1.19489171e-08 1.73090774e-07 1.19564856e-08 1.73190774e-07 1.19492572e-08
+ 1.73290774e-07 1.19561605e-08 1.73390774e-07 1.19495682e-08 1.73490774e-07 1.19558634e-08 1.73590774e-07 1.19498513e-08 1.73690774e-07 1.19555937e-08 1.73790774e-07 1.19501088e-08 1.73890774e-07 1.19553474e-08 1.73990774e-07 1.19503443e-08
+ 1.74090774e-07 1.19551221e-08 1.74190774e-07 1.19505598e-08 1.74290774e-07 1.1954916e-08 1.74390774e-07 1.19507568e-08 1.74490774e-07 1.19547276e-08 1.74590774e-07 1.19509369e-08 1.74690774e-07 1.19545555e-08 1.74790774e-07 1.19511014e-08
+ 1.74890774e-07 1.1954398e-08 1.74990774e-07 1.19512519e-08 1.75090774e-07 1.19542541e-08 1.75190774e-07 1.19513894e-08 1.75290774e-07 1.1954123e-08 1.75390774e-07 1.19515147e-08 1.75490774e-07 1.19540033e-08 1.75590774e-07 1.19516285e-08
+ 1.75690774e-07 1.19538951e-08 1.75790774e-07 1.19517321e-08 1.75890774e-07 1.19537961e-08 1.75990774e-07 1.19518266e-08 1.76090774e-07 1.19537054e-08 1.76190774e-07 1.19519137e-08 1.76290774e-07 1.19536226e-08 1.76390774e-07 1.19519931e-08
+ 1.76490774e-07 1.19535465e-08 1.76590774e-07 1.19520655e-08 1.76690774e-07 1.19534773e-08 1.76790774e-07 1.19521314e-08 1.76890774e-07 1.19534144e-08 1.76990774e-07 1.19521917e-08 1.77090774e-07 1.19533567e-08 1.77190774e-07 1.19522465e-08
+ 1.77290774e-07 1.19533046e-08 1.77390774e-07 1.19522966e-08 1.77490774e-07 1.19532571e-08 1.77590774e-07 1.19523421e-08 1.77690774e-07 1.19532133e-08 1.77790774e-07 1.19523835e-08 1.77890774e-07 1.19531737e-08 1.77990774e-07 1.19524212e-08
+ 1.78090774e-07 1.19531379e-08 1.78190774e-07 1.19524555e-08 1.78290774e-07 1.1953105e-08 1.78390774e-07 1.19524866e-08 1.78490774e-07 1.19530755e-08 1.78590774e-07 1.19525148e-08 1.78690774e-07 1.19530485e-08 1.78790774e-07 1.19525405e-08
+ 1.78890774e-07 1.19530244e-08 1.78990774e-07 1.19525634e-08 1.79090774e-07 1.19530023e-08 1.79190774e-07 1.19525844e-08 1.79290774e-07 1.19529825e-08 1.79390774e-07 1.19526031e-08 1.79490774e-07 1.19529646e-08 1.79590774e-07 1.19526204e-08
+ 1.79690774e-07 1.19529481e-08 1.79790774e-07 1.19526362e-08 1.79890774e-07 1.19529332e-08 1.79990774e-07 1.19526501e-08 1.80090774e-07 1.19529197e-08 1.80190774e-07 1.19526631e-08 1.80290774e-07 1.19529075e-08 1.80390774e-07 1.19526747e-08
+ 1.80490774e-07 1.19528963e-08 1.80590774e-07 1.19526854e-08 1.80690774e-07 1.19528863e-08 1.80790774e-07 1.1952695e-08 1.80890774e-07 1.19528772e-08 1.80990774e-07 1.19527035e-08 1.81090774e-07 1.1952869e-08 1.81190774e-07 1.19527115e-08
+ 1.81290774e-07 1.19528619e-08 1.81390774e-07 1.19527184e-08 1.81490774e-07 1.1952855e-08 1.81590774e-07 1.19527248e-08 1.81690774e-07 1.19528489e-08 1.81790774e-07 1.19527304e-08 1.81890774e-07 1.19528434e-08 1.81990774e-07 1.1952736e-08
+ 1.82090774e-07 1.19528385e-08 1.82190774e-07 1.19527407e-08 1.82290774e-07 1.19528338e-08 1.82390774e-07 1.19527451e-08 1.82490774e-07 1.19528294e-08 1.82590774e-07 1.1952749e-08 1.82690774e-07 1.19528259e-08 1.82790774e-07 1.19527526e-08
+ 1.82890774e-07 1.19528223e-08 1.82990774e-07 1.19527557e-08 1.83090774e-07 1.19528194e-08 1.83190774e-07 1.19527588e-08 1.83290774e-07 1.19528165e-08 1.83390774e-07 1.19527615e-08 1.83490774e-07 1.19528138e-08 1.83590774e-07 1.19527637e-08
+ 1.83690774e-07 1.19528119e-08 1.83790774e-07 1.19527659e-08 1.83890774e-07 1.19528098e-08 1.83990774e-07 1.19527681e-08 1.84090774e-07 1.19528076e-08 1.84190774e-07 1.19527698e-08 1.84290774e-07 1.19528059e-08 1.84390774e-07 1.19527714e-08
+ 1.84490774e-07 1.19528044e-08 1.84590774e-07 1.1952773e-08 1.84690774e-07 1.1952803e-08 1.84790774e-07 1.19527743e-08 1.84890774e-07 1.19528015e-08 1.84990774e-07 1.19527756e-08 1.85090774e-07 1.19528004e-08 1.85190774e-07 1.19527767e-08
+ 1.85290774e-07 1.19527994e-08 1.85390774e-07 1.19527779e-08 1.85490774e-07 1.19527985e-08 1.85590774e-07 1.19527787e-08 1.85690774e-07 1.19527974e-08 1.85790774e-07 1.19527794e-08 1.85890774e-07 1.19527966e-08 1.85990774e-07 1.19527802e-08
+ 1.86090774e-07 1.19527959e-08 1.86190774e-07 1.19527811e-08 1.86290774e-07 1.19527951e-08 1.86390774e-07 1.1952782e-08 1.86490774e-07 1.19527945e-08 1.86590774e-07 1.19527821e-08 1.86690774e-07 1.1952794e-08 1.86790774e-07 1.19527827e-08
+ 1.86890774e-07 1.19527934e-08 1.86990774e-07 1.19527833e-08 1.87090774e-07 1.19527932e-08 1.87190774e-07 1.19527837e-08 1.87290774e-07 1.19527928e-08 1.87390774e-07 1.19527838e-08 1.87490774e-07 1.19527925e-08 1.87590774e-07 1.19527841e-08
+ 1.87690774e-07 1.19527923e-08 1.87790774e-07 1.19527845e-08 1.87890774e-07 1.19527921e-08 1.87990774e-07 1.19527847e-08 1.88090774e-07 1.19527917e-08 1.88190774e-07 1.1952785e-08 1.88290774e-07 1.19527915e-08 1.88390774e-07 1.19527853e-08
+ 1.88490774e-07 1.19527913e-08 1.88590774e-07 1.19527857e-08 1.88690774e-07 1.19527911e-08 1.88790774e-07 1.19527857e-08 1.88890774e-07 1.19527905e-08 1.88990774e-07 1.1952786e-08 1.89090774e-07 1.19527906e-08 1.89190774e-07 1.19527863e-08
+ 1.89290774e-07 1.195279e-08 1.89390774e-07 1.19527864e-08 1.89490774e-07 1.19527903e-08 1.89590774e-07 1.19527866e-08 1.89690774e-07 1.19527896e-08 1.89790774e-07 1.19527868e-08 1.89890774e-07 1.19527898e-08 1.89990774e-07 1.19527869e-08
+ 1.90090774e-07 1.19527897e-08 1.90190774e-07 1.1952787e-08 1.90290774e-07 1.19527896e-08 1.90390774e-07 1.19527871e-08 1.90490774e-07 1.19527896e-08 1.90590774e-07 1.1952787e-08 1.90690774e-07 1.19527896e-08 1.90790774e-07 1.19527872e-08
+ 1.90890774e-07 1.19527894e-08 1.90990774e-07 1.19527873e-08 1.91090774e-07 1.19527893e-08 1.91190774e-07 1.19527874e-08 1.91290774e-07 1.19527891e-08 1.91390774e-07 1.19527875e-08 1.91490774e-07 1.19527892e-08 1.91590774e-07 1.19527877e-08
+ 1.91690774e-07 1.1952789e-08 1.91790774e-07 1.19527876e-08 1.91890774e-07 1.19527889e-08 1.91990774e-07 1.19527877e-08 1.92090774e-07 1.19527888e-08 1.92190774e-07 1.19527879e-08 1.92290774e-07 1.19527889e-08 1.92390774e-07 1.19527878e-08
+ 1.92490774e-07 1.19527887e-08 1.92590774e-07 1.1952788e-08 1.92690774e-07 1.19527889e-08 1.92790774e-07 1.19527879e-08 1.92890774e-07 1.19527888e-08 1.92990774e-07 1.19527879e-08 1.93090774e-07 1.19527889e-08 1.93190774e-07 1.19527879e-08
+ 1.93290774e-07 1.19527889e-08 1.93390774e-07 1.19527877e-08 1.93490774e-07 1.19527885e-08 1.93590774e-07 1.19527878e-08 1.93690774e-07 1.19527886e-08 1.93790774e-07 1.1952788e-08 1.93890774e-07 1.19527888e-08 1.93990774e-07 1.1952788e-08
+ 1.94090774e-07 1.19527889e-08 1.94190774e-07 1.1952788e-08 1.94290774e-07 1.19527888e-08 1.94390774e-07 1.19527879e-08 1.94490774e-07 1.19527886e-08 1.94590774e-07 1.1952788e-08 1.94690774e-07 1.19527889e-08 1.94790774e-07 1.1952788e-08
+ 1.94890774e-07 1.19527888e-08 1.94990774e-07 1.19527881e-08 1.95090774e-07 1.19527887e-08 1.95190774e-07 1.19527879e-08 1.95290774e-07 1.19527886e-08 1.95390774e-07 1.1952788e-08 1.95490774e-07 1.19527888e-08 1.95590774e-07 1.19527881e-08
+ 1.95690774e-07 1.19527887e-08 1.95790774e-07 1.19527881e-08 1.95890774e-07 1.19527888e-08 1.95990774e-07 1.19527881e-08 1.96090774e-07 1.19527885e-08 1.96190774e-07 1.19527883e-08 1.96290774e-07 1.19527884e-08 1.96390774e-07 1.1952788e-08
+ 1.96490774e-07 1.19527882e-08 1.96590774e-07 1.1952788e-08 1.96690774e-07 1.19527883e-08 1.96790774e-07 1.19527879e-08 1.96890774e-07 1.19527884e-08 1.96990774e-07 1.1952788e-08 1.97090774e-07 1.19527883e-08 1.97190774e-07 1.1952788e-08
+ 1.97290774e-07 1.19527884e-08 1.97390774e-07 1.1952788e-08 1.97490774e-07 1.19527884e-08 1.97590774e-07 1.1952788e-08 1.97690774e-07 1.19527883e-08 1.97790774e-07 1.1952788e-08 1.97890774e-07 1.19527884e-08 1.97990774e-07 1.19527879e-08
+ 1.98090774e-07 1.19527884e-08 1.98190774e-07 1.1952788e-08 1.98290774e-07 1.19527882e-08 1.98390774e-07 1.1952788e-08 1.98490774e-07 1.19527884e-08 1.98590774e-07 1.1952788e-08 1.98690774e-07 1.19527883e-08 1.98790774e-07 1.1952788e-08
+ 1.98890774e-07 1.19527884e-08 1.98990774e-07 1.19527881e-08 1.99090774e-07 1.19527883e-08 1.99190774e-07 1.19527881e-08 1.99290774e-07 1.19527885e-08 1.99390774e-07 1.19527879e-08 1.99490774e-07 1.19527885e-08 1.99590774e-07 1.19527879e-08
+ 1.99690774e-07 1.19527885e-08 1.99790774e-07 1.19527879e-08 1.99890774e-07 1.19527884e-08 1.99990774e-07 1.1952788e-08 2e-07 1.19527885e-08 2.0001e-07 1.19810074e-08 2.0003e-07 1.18152688e-08 2.0007e-07 1.21656675e-08
+ 2.0015e-07 1.1714175e-08 2.0025e-07 1.21973737e-08 2.0035e-07 1.17166001e-08 2.0045e-07 1.21670031e-08 2.0055e-07 1.1777596e-08 2.0065e-07 1.18484742e-08 2.0075e-07 2.53191128e-08 2.0085e-07 -4.04759482e-07
+ 2.00932239e-07 6.49708168e-06 2.01e-07 -4.94343878e-05 2.01008502e-07 -5.0992026e-05 2.01025505e-07 -4.39145059e-05 2.01059511e-07 -1.62206912e-05 2.01090728e-07 0.000285043155 2.01143656e-07 0.000513849787 2.01199398e-07 0.00155348227
+ 2.01276452e-07 -0.0180250591 2.01342062e-07 -0.00339007548 2.01411951e-07 3.25710063 2.01487979e-07 4.90275261 2.01566956e-07 5.02684152 2.01643585e-07 4.98988775 2.01743585e-07 5.00539209 2.01843585e-07 4.99682771
+ 2.01943585e-07 5.00195612 2.02043585e-07 4.99873104 2.02143585e-07 5.00083562 2.02243585e-07 4.99943657 2.02343585e-07 5.00037969 2.02443585e-07 4.99974066 2.02543585e-07 5.00017605 2.02643585e-07 4.99987923
+ 2.02743585e-07 5.00008215 2.02843585e-07 4.99994356 2.02943585e-07 5.00003839 2.03043585e-07 4.9999736 2.03143585e-07 5.00001792 2.03243585e-07 4.99998767 2.03343585e-07 5.00000832 2.03443585e-07 4.99999427
+ 2.03543585e-07 5.00000382 2.03643585e-07 4.99999736 2.03743585e-07 5.00000171 2.03843585e-07 4.99999881 2.03943585e-07 5.00000073 2.04043585e-07 4.99999949 2.04143585e-07 5.00000027 2.04243585e-07 4.9999998
+ 2.04343585e-07 5.00000006 2.04443585e-07 4.99999994 2.04543585e-07 4.99999996 2.04643585e-07 5.0 2.04743585e-07 4.99999993 2.04843585e-07 5.00000002 2.04943585e-07 4.99999992 2.05043585e-07 5.00000003
+ 2.05143585e-07 4.99999992 2.05243585e-07 5.00000003 2.05343585e-07 4.99999992 2.05443585e-07 5.00000002 2.05543585e-07 4.99999993 2.05643585e-07 5.00000001 2.05743585e-07 4.99999993 2.05843585e-07 5.00000001
+ 2.05943585e-07 4.99999994 2.06043585e-07 5.0 2.06143585e-07 4.99999994 2.06243585e-07 5.0 2.06343585e-07 4.99999995 2.06443585e-07 4.99999999 2.06543585e-07 4.99999995 2.06643585e-07 4.99999999
+ 2.06743585e-07 4.99999996 2.06843585e-07 4.99999999 2.06943585e-07 4.99999996 2.07043585e-07 4.99999998 2.07143585e-07 4.99999996 2.07243585e-07 4.99999998 2.07343585e-07 4.99999996 2.07443585e-07 4.99999998
+ 2.07543585e-07 4.99999996 2.07643585e-07 4.99999998 2.07743585e-07 4.99999997 2.07843585e-07 4.99999998 2.07943585e-07 4.99999997 2.08043585e-07 4.99999998 2.08143585e-07 4.99999997 2.08243585e-07 4.99999998
+ 2.08343585e-07 4.99999997 2.08443585e-07 4.99999998 2.08543585e-07 4.99999997 2.08643585e-07 4.99999997 2.08743585e-07 4.99999997 2.08843585e-07 4.99999997 2.08943585e-07 4.99999997 2.09043585e-07 4.99999997
+ 2.09143585e-07 4.99999997 2.09243585e-07 4.99999997 2.09343585e-07 4.99999997 2.09443585e-07 4.99999997 2.09543585e-07 4.99999997 2.09643585e-07 4.99999997 2.09743585e-07 4.99999997 2.09843585e-07 4.99999997
+ 2.09943585e-07 4.99999997 2.10043585e-07 4.99999997 2.10143585e-07 4.99999997 2.10243585e-07 4.99999997 2.10343585e-07 4.99999997 2.10443585e-07 4.99999997 2.10543585e-07 4.99999997 2.10643585e-07 4.99999997
+ 2.10743585e-07 4.99999997 2.10843585e-07 4.99999997 2.10943585e-07 4.99999997 2.11043585e-07 4.99999997 2.11143585e-07 4.99999997 2.11243585e-07 4.99999997 2.11343585e-07 4.99999997 2.11443585e-07 4.99999997
+ 2.11543585e-07 4.99999997 2.11643585e-07 4.99999997 2.11743585e-07 4.99999997 2.11843585e-07 4.99999997 2.11943585e-07 4.99999997 2.12043585e-07 4.99999997 2.12143585e-07 4.99999997 2.12243585e-07 4.99999997
+ 2.12343585e-07 4.99999997 2.12443585e-07 4.99999997 2.12543585e-07 4.99999997 2.12643585e-07 4.99999997 2.12743585e-07 4.99999997 2.12843585e-07 4.99999997 2.12943585e-07 4.99999997 2.13043585e-07 4.99999997
+ 2.13143585e-07 4.99999997 2.13243585e-07 4.99999997 2.13343585e-07 4.99999997 2.13443585e-07 4.99999997 2.13543585e-07 4.99999997 2.13643585e-07 4.99999997 2.13743585e-07 4.99999997 2.13843585e-07 4.99999997
+ 2.13943585e-07 4.99999997 2.14043585e-07 4.99999997 2.14143585e-07 4.99999997 2.14243585e-07 4.99999997 2.14343585e-07 4.99999997 2.14443585e-07 4.99999997 2.14543585e-07 4.99999997 2.14643585e-07 4.99999997
+ 2.14743585e-07 4.99999997 2.14843585e-07 4.99999997 2.14943585e-07 4.99999997 2.15043585e-07 4.99999997 2.15143585e-07 4.99999997 2.15243585e-07 4.99999997 2.15343585e-07 4.99999997 2.15443585e-07 4.99999997
+ 2.15543585e-07 4.99999997 2.15643585e-07 4.99999997 2.15743585e-07 4.99999997 2.15843585e-07 4.99999997 2.15943585e-07 4.99999997 2.16043585e-07 4.99999997 2.16143585e-07 4.99999997 2.16243585e-07 4.99999997
+ 2.16343585e-07 4.99999997 2.16443585e-07 4.99999997 2.16543585e-07 4.99999997 2.16643585e-07 4.99999997 2.16743585e-07 4.99999997 2.16843585e-07 4.99999997 2.16943585e-07 4.99999997 2.17043585e-07 4.99999997
+ 2.17143585e-07 4.99999997 2.17243585e-07 4.99999997 2.17343585e-07 4.99999997 2.17443585e-07 4.99999997 2.17543585e-07 4.99999997 2.17643585e-07 4.99999997 2.17743585e-07 4.99999997 2.17843585e-07 4.99999997
+ 2.17943585e-07 4.99999997 2.18043585e-07 4.99999997 2.18143585e-07 4.99999997 2.18243585e-07 4.99999997 2.18343585e-07 4.99999997 2.18443585e-07 4.99999997 2.18543585e-07 4.99999997 2.18643585e-07 4.99999997
+ 2.18743585e-07 4.99999997 2.18843585e-07 4.99999997 2.18943585e-07 4.99999997 2.19043585e-07 4.99999997 2.19143585e-07 4.99999997 2.19243585e-07 4.99999997 2.19343585e-07 4.99999997 2.19443585e-07 4.99999997
+ 2.19543585e-07 4.99999997 2.19643585e-07 4.99999997 2.19743585e-07 4.99999997 2.19843585e-07 4.99999997 2.19943585e-07 4.99999997 2.20043585e-07 4.99999997 2.20143585e-07 4.99999997 2.20243585e-07 4.99999997
+ 2.20343585e-07 4.99999997 2.20443585e-07 4.99999997 2.20543585e-07 4.99999997 2.20643585e-07 4.99999997 2.20743585e-07 4.99999997 2.20843585e-07 4.99999997 2.20943585e-07 4.99999997 2.21043585e-07 4.99999997
+ 2.21143585e-07 4.99999997 2.21243585e-07 4.99999997 2.21343585e-07 4.99999997 2.21443585e-07 4.99999997 2.21543585e-07 4.99999997 2.21643585e-07 4.99999997 2.21743585e-07 4.99999997 2.21843585e-07 4.99999997
+ 2.21943585e-07 4.99999997 2.22043585e-07 4.99999997 2.22143585e-07 4.99999997 2.22243585e-07 4.99999997 2.22343585e-07 4.99999997 2.22443585e-07 4.99999997 2.22543585e-07 4.99999997 2.22643585e-07 4.99999997
+ 2.22743585e-07 4.99999997 2.22843585e-07 4.99999997 2.22943585e-07 4.99999997 2.23043585e-07 4.99999997 2.23143585e-07 4.99999997 2.23243585e-07 4.99999997 2.23343585e-07 4.99999997 2.23443585e-07 4.99999997
+ 2.23543585e-07 4.99999997 2.23643585e-07 4.99999997 2.23743585e-07 4.99999997 2.23843585e-07 4.99999997 2.23943585e-07 4.99999997 2.24043585e-07 4.99999997 2.24143585e-07 4.99999997 2.24243585e-07 4.99999997
+ 2.24343585e-07 4.99999997 2.24443585e-07 4.99999997 2.24543585e-07 4.99999997 2.24643585e-07 4.99999997 2.24743585e-07 4.99999997 2.24843585e-07 4.99999997 2.24943585e-07 4.99999997 2.25043585e-07 4.99999997
+ 2.25143585e-07 4.99999997 2.25243585e-07 4.99999997 2.25343585e-07 4.99999997 2.25443585e-07 4.99999997 2.25543585e-07 4.99999997 2.25643585e-07 4.99999997 2.25743585e-07 4.99999997 2.25843585e-07 4.99999997
+ 2.25943585e-07 4.99999997 2.26043585e-07 4.99999997 2.26143585e-07 4.99999997 2.26243585e-07 4.99999997 2.26343585e-07 4.99999997 2.26443585e-07 4.99999997 2.26543585e-07 4.99999997 2.26643585e-07 4.99999997
+ 2.26743585e-07 4.99999997 2.26843585e-07 4.99999997 2.26943585e-07 4.99999997 2.27043585e-07 4.99999997 2.27143585e-07 4.99999997 2.27243585e-07 4.99999997 2.27343585e-07 4.99999997 2.27443585e-07 4.99999997
+ 2.27543585e-07 4.99999997 2.27643585e-07 4.99999997 2.27743585e-07 4.99999997 2.27843585e-07 4.99999997 2.27943585e-07 4.99999997 2.28043585e-07 4.99999997 2.28143585e-07 4.99999997 2.28243585e-07 4.99999997
+ 2.28343585e-07 4.99999997 2.28443585e-07 4.99999997 2.28543585e-07 4.99999997 2.28643585e-07 4.99999997 2.28743585e-07 4.99999997 2.28843585e-07 4.99999997 2.28943585e-07 4.99999997 2.29043585e-07 4.99999997
+ 2.29143585e-07 4.99999997 2.29243585e-07 4.99999997 2.29343585e-07 4.99999997 2.29443585e-07 4.99999997 2.29543585e-07 4.99999997 2.29643585e-07 4.99999997 2.29743585e-07 4.99999997 2.29843585e-07 4.99999997
+ 2.29943585e-07 4.99999997 2.30043585e-07 4.99999997 2.30143585e-07 4.99999997 2.30243585e-07 4.99999997 2.30343585e-07 4.99999997 2.30443585e-07 4.99999997 2.30543585e-07 4.99999997 2.30643585e-07 4.99999997
+ 2.30743585e-07 4.99999997 2.30843585e-07 4.99999997 2.30943585e-07 4.99999997 2.31043585e-07 4.99999997 2.31143585e-07 4.99999997 2.31243585e-07 4.99999997 2.31343585e-07 4.99999997 2.31443585e-07 4.99999997
+ 2.31543585e-07 4.99999997 2.31643585e-07 4.99999997 2.31743585e-07 4.99999997 2.31843585e-07 4.99999997 2.31943585e-07 4.99999997 2.32043585e-07 4.99999997 2.32143585e-07 4.99999997 2.32243585e-07 4.99999997
+ 2.32343585e-07 4.99999997 2.32443585e-07 4.99999997 2.32543585e-07 4.99999997 2.32643585e-07 4.99999997 2.32743585e-07 4.99999997 2.32843585e-07 4.99999997 2.32943585e-07 4.99999997 2.33043585e-07 4.99999997
+ 2.33143585e-07 4.99999997 2.33243585e-07 4.99999997 2.33343585e-07 4.99999997 2.33443585e-07 4.99999997 2.33543585e-07 4.99999997 2.33643585e-07 4.99999997 2.33743585e-07 4.99999997 2.33843585e-07 4.99999997
+ 2.33943585e-07 4.99999997 2.34043585e-07 4.99999997 2.34143585e-07 4.99999997 2.34243585e-07 4.99999997 2.34343585e-07 4.99999997 2.34443585e-07 4.99999997 2.34543585e-07 4.99999997 2.34643585e-07 4.99999997
+ 2.34743585e-07 4.99999997 2.34843585e-07 4.99999997 2.34943585e-07 4.99999997 2.35043585e-07 4.99999997 2.35143585e-07 4.99999997 2.35243585e-07 4.99999997 2.35343585e-07 4.99999997 2.35443585e-07 4.99999997
+ 2.35543585e-07 4.99999997 2.35643585e-07 4.99999997 2.35743585e-07 4.99999997 2.35843585e-07 4.99999997 2.35943585e-07 4.99999997 2.36043585e-07 4.99999997 2.36143585e-07 4.99999997 2.36243585e-07 4.99999997
+ 2.36343585e-07 4.99999997 2.36443585e-07 4.99999997 2.36543585e-07 4.99999997 2.36643585e-07 4.99999997 2.36743585e-07 4.99999997 2.36843585e-07 4.99999997 2.36943585e-07 4.99999997 2.37043585e-07 4.99999997
+ 2.37143585e-07 4.99999997 2.37243585e-07 4.99999997 2.37343585e-07 4.99999997 2.37443585e-07 4.99999997 2.37543585e-07 4.99999997 2.37643585e-07 4.99999997 2.37743585e-07 4.99999997 2.37843585e-07 4.99999997
+ 2.37943585e-07 4.99999997 2.38043585e-07 4.99999997 2.38143585e-07 4.99999997 2.38243585e-07 4.99999997 2.38343585e-07 4.99999997 2.38443585e-07 4.99999997 2.38543585e-07 4.99999997 2.38643585e-07 4.99999997
+ 2.38743585e-07 4.99999997 2.38843585e-07 4.99999997 2.38943585e-07 4.99999997 2.39043585e-07 4.99999997 2.39143585e-07 4.99999997 2.39243585e-07 4.99999997 2.39343585e-07 4.99999997 2.39443585e-07 4.99999997
+ 2.39543585e-07 4.99999997 2.39643585e-07 4.99999997 2.39743585e-07 4.99999997 2.39843585e-07 4.99999997 2.39943585e-07 4.99999997 2.40043585e-07 4.99999997 2.40143585e-07 4.99999997 2.40243585e-07 4.99999997
+ 2.40343585e-07 4.99999997 2.40443585e-07 4.99999997 2.40543585e-07 4.99999997 2.40643585e-07 4.99999997 2.40743585e-07 4.99999997 2.40843585e-07 4.99999997 2.40943585e-07 4.99999997 2.41043585e-07 4.99999997
+ 2.41143585e-07 4.99999997 2.41243585e-07 4.99999997 2.41343585e-07 4.99999997 2.41443585e-07 4.99999997 2.41543585e-07 4.99999997 2.41643585e-07 4.99999997 2.41743585e-07 4.99999997 2.41843585e-07 4.99999997
+ 2.41943585e-07 4.99999997 2.42043585e-07 4.99999997 2.42143585e-07 4.99999997 2.42243585e-07 4.99999997 2.42343585e-07 4.99999997 2.42443585e-07 4.99999997 2.42543585e-07 4.99999997 2.42643585e-07 4.99999997
+ 2.42743585e-07 4.99999997 2.42843585e-07 4.99999997 2.42943585e-07 4.99999997 2.43043585e-07 4.99999997 2.43143585e-07 4.99999997 2.43243585e-07 4.99999997 2.43343585e-07 4.99999997 2.43443585e-07 4.99999997
+ 2.43543585e-07 4.99999997 2.43643585e-07 4.99999997 2.43743585e-07 4.99999997 2.43843585e-07 4.99999997 2.43943585e-07 4.99999997 2.44043585e-07 4.99999997 2.44143585e-07 4.99999997 2.44243585e-07 4.99999997
+ 2.44343585e-07 4.99999997 2.44443585e-07 4.99999997 2.44543585e-07 4.99999997 2.44643585e-07 4.99999997 2.44743585e-07 4.99999997 2.44843585e-07 4.99999997 2.44943585e-07 4.99999997 2.45043585e-07 4.99999997
+ 2.45143585e-07 4.99999997 2.45243585e-07 4.99999997 2.45343585e-07 4.99999997 2.45443585e-07 4.99999997 2.45543585e-07 4.99999997 2.45643585e-07 4.99999997 2.45743585e-07 4.99999997 2.45843585e-07 4.99999997
+ 2.45943585e-07 4.99999997 2.46043585e-07 4.99999997 2.46143585e-07 4.99999997 2.46243585e-07 4.99999997 2.46343585e-07 4.99999997 2.46443585e-07 4.99999997 2.46543585e-07 4.99999997 2.46643585e-07 4.99999997
+ 2.46743585e-07 4.99999997 2.46843585e-07 4.99999997 2.46943585e-07 4.99999997 2.47043585e-07 4.99999997 2.47143585e-07 4.99999997 2.47243585e-07 4.99999997 2.47343585e-07 4.99999997 2.47443585e-07 4.99999997
+ 2.47543585e-07 4.99999997 2.47643585e-07 4.99999997 2.47743585e-07 4.99999997 2.47843585e-07 4.99999997 2.47943585e-07 4.99999997 2.48043585e-07 4.99999997 2.48143585e-07 4.99999997 2.48243585e-07 4.99999997
+ 2.48343585e-07 4.99999997 2.48443585e-07 4.99999997 2.48543585e-07 4.99999997 2.48643585e-07 4.99999997 2.48743585e-07 4.99999997 2.48843585e-07 4.99999997 2.48943585e-07 4.99999997 2.49043585e-07 4.99999997
+ 2.49143585e-07 4.99999997 2.49243585e-07 4.99999997 2.49343585e-07 4.99999997 2.49443585e-07 4.99999997 2.49543585e-07 4.99999997 2.49643585e-07 4.99999997 2.49743585e-07 4.99999997 2.49843585e-07 4.99999997
+ 2.49943585e-07 4.99999997 2.50043585e-07 4.99999997 2.50143585e-07 4.99999997 2.50243585e-07 4.99999997 2.50343585e-07 4.99999997 2.50443585e-07 4.99999997 2.50543585e-07 4.99999997 2.50643585e-07 4.99999997
+ 2.50743585e-07 4.99999997 2.50843585e-07 4.99999997 2.50943585e-07 4.99999997 2.51e-07 4.99999997 2.5101e-07 4.99999997 2.5103e-07 4.99999997 2.5107e-07 4.99999997 2.5115e-07 4.99999997
+ 2.5125e-07 4.99999997 2.5135e-07 4.99999997 2.5145e-07 4.99999997 2.5155e-07 4.99999997 2.5165e-07 4.99999997 2.5175e-07 4.99999997 2.5185e-07 4.99999997 2.51930828e-07 5.00000127
+ 2.52e-07 5.00000077 2.52008608e-07 4.99998869 2.52025825e-07 4.99996401 2.52060258e-07 5.00000369 2.52106181e-07 5.00005267 2.52150081e-07 4.99998208 2.52198026e-07 4.9999678 2.5225538e-07 5.00001892
+ 2.52312019e-07 4.99999862 2.52404231e-07 5.00000003 2.52504231e-07 5.00000076 2.52604231e-07 4.99999856 2.52704231e-07 5.00000151 2.52804231e-07 4.99999846 2.52904231e-07 5.00000136 2.53004231e-07 4.99999873
+ 2.53104231e-07 5.00000105 2.53204231e-07 4.99999904 2.53304231e-07 5.00000077 2.53404231e-07 4.99999929 2.53504231e-07 5.00000056 2.53604231e-07 4.99999946 2.53704231e-07 5.00000041 2.53804231e-07 4.99999959
+ 2.53904231e-07 5.00000031 2.54004231e-07 4.99999967 2.54104231e-07 5.00000024 2.54204231e-07 4.99999973 2.54304231e-07 5.00000019 2.54404231e-07 4.99999977 2.54504231e-07 5.00000015 2.54604231e-07 4.99999981
+ 2.54704231e-07 5.00000013 2.54804231e-07 4.99999983 2.54904231e-07 5.0000001 2.55004231e-07 4.99999985 2.55104231e-07 5.00000009 2.55204231e-07 4.99999987 2.55304231e-07 5.00000007 2.55404231e-07 4.99999988
+ 2.55504231e-07 5.00000006 2.55604231e-07 4.99999989 2.55704231e-07 5.00000005 2.55804231e-07 4.9999999 2.55904231e-07 5.00000004 2.56004231e-07 4.99999991 2.56104231e-07 5.00000003 2.56204231e-07 4.99999992
+ 2.56304231e-07 5.00000003 2.56404231e-07 4.99999992 2.56504231e-07 5.00000002 2.56604231e-07 4.99999993 2.56704231e-07 5.00000001 2.56804231e-07 4.99999993 2.56904231e-07 5.00000001 2.57004231e-07 4.99999994
+ 2.57104231e-07 5.0 2.57204231e-07 4.99999994 2.57304231e-07 5.0 2.57404231e-07 4.99999994 2.57504231e-07 5.0 2.57604231e-07 4.99999995 2.57704231e-07 4.99999999 2.57804231e-07 4.99999995
+ 2.57904231e-07 4.99999999 2.58004231e-07 4.99999995 2.58104231e-07 4.99999999 2.58204231e-07 4.99999996 2.58304231e-07 4.99999999 2.58404231e-07 4.99999996 2.58504231e-07 4.99999999 2.58604231e-07 4.99999996
+ 2.58704231e-07 4.99999998 2.58804231e-07 4.99999996 2.58904231e-07 4.99999998 2.59004231e-07 4.99999996 2.59104231e-07 4.99999998 2.59204231e-07 4.99999996 2.59304231e-07 4.99999998 2.59404231e-07 4.99999996
+ 2.59504231e-07 4.99999998 2.59604231e-07 4.99999996 2.59704231e-07 4.99999998 2.59804231e-07 4.99999997 2.59904231e-07 4.99999998 2.60004231e-07 4.99999997 2.60104231e-07 4.99999998 2.60204231e-07 4.99999997
+ 2.60304231e-07 4.99999998 2.60404231e-07 4.99999997 2.60504231e-07 4.99999998 2.60604231e-07 4.99999997 2.60704231e-07 4.99999998 2.60804231e-07 4.99999997 2.60904231e-07 4.99999998 2.61004231e-07 4.99999997
+ 2.61104231e-07 4.99999998 2.61204231e-07 4.99999997 2.61304231e-07 4.99999997 2.61404231e-07 4.99999997 2.61504231e-07 4.99999997 2.61604231e-07 4.99999997 2.61704231e-07 4.99999997 2.61804231e-07 4.99999997
+ 2.61904231e-07 4.99999997 2.62004231e-07 4.99999997 2.62104231e-07 4.99999997 2.62204231e-07 4.99999997 2.62304231e-07 4.99999997 2.62404231e-07 4.99999997 2.62504231e-07 4.99999997 2.62604231e-07 4.99999997
+ 2.62704231e-07 4.99999997 2.62804231e-07 4.99999997 2.62904231e-07 4.99999997 2.63004231e-07 4.99999997 2.63104231e-07 4.99999997 2.63204231e-07 4.99999997 2.63304231e-07 4.99999997 2.63404231e-07 4.99999997
+ 2.63504231e-07 4.99999997 2.63604231e-07 4.99999997 2.63704231e-07 4.99999997 2.63804231e-07 4.99999997 2.63904231e-07 4.99999997 2.64004231e-07 4.99999997 2.64104231e-07 4.99999997 2.64204231e-07 4.99999997
+ 2.64304231e-07 4.99999997 2.64404231e-07 4.99999997 2.64504231e-07 4.99999997 2.64604231e-07 4.99999997 2.64704231e-07 4.99999997 2.64804231e-07 4.99999997 2.64904231e-07 4.99999997 2.65004231e-07 4.99999997
+ 2.65104231e-07 4.99999997 2.65204231e-07 4.99999997 2.65304231e-07 4.99999997 2.65404231e-07 4.99999997 2.65504231e-07 4.99999997 2.65604231e-07 4.99999997 2.65704231e-07 4.99999997 2.65804231e-07 4.99999997
+ 2.65904231e-07 4.99999997 2.66004231e-07 4.99999997 2.66104231e-07 4.99999997 2.66204231e-07 4.99999997 2.66304231e-07 4.99999997 2.66404231e-07 4.99999997 2.66504231e-07 4.99999997 2.66604231e-07 4.99999997
+ 2.66704231e-07 4.99999997 2.66804231e-07 4.99999997 2.66904231e-07 4.99999997 2.67004231e-07 4.99999997 2.67104231e-07 4.99999997 2.67204231e-07 4.99999997 2.67304231e-07 4.99999997 2.67404231e-07 4.99999997
+ 2.67504231e-07 4.99999997 2.67604231e-07 4.99999997 2.67704231e-07 4.99999997 2.67804231e-07 4.99999997 2.67904231e-07 4.99999997 2.68004231e-07 4.99999997 2.68104231e-07 4.99999997 2.68204231e-07 4.99999997
+ 2.68304231e-07 4.99999997 2.68404231e-07 4.99999997 2.68504231e-07 4.99999997 2.68604231e-07 4.99999997 2.68704231e-07 4.99999997 2.68804231e-07 4.99999997 2.68904231e-07 4.99999997 2.69004231e-07 4.99999997
+ 2.69104231e-07 4.99999997 2.69204231e-07 4.99999997 2.69304231e-07 4.99999997 2.69404231e-07 4.99999997 2.69504231e-07 4.99999997 2.69604231e-07 4.99999997 2.69704231e-07 4.99999997 2.69804231e-07 4.99999997
+ 2.69904231e-07 4.99999997 2.70004231e-07 4.99999997 2.70104231e-07 4.99999997 2.70204231e-07 4.99999997 2.70304231e-07 4.99999997 2.70404231e-07 4.99999997 2.70504231e-07 4.99999997 2.70604231e-07 4.99999997
+ 2.70704231e-07 4.99999997 2.70804231e-07 4.99999997 2.70904231e-07 4.99999997 2.71004231e-07 4.99999997 2.71104231e-07 4.99999997 2.71204231e-07 4.99999997 2.71304231e-07 4.99999997 2.71404231e-07 4.99999997
+ 2.71504231e-07 4.99999997 2.71604231e-07 4.99999997 2.71704231e-07 4.99999997 2.71804231e-07 4.99999997 2.71904231e-07 4.99999997 2.72004231e-07 4.99999997 2.72104231e-07 4.99999997 2.72204231e-07 4.99999997
+ 2.72304231e-07 4.99999997 2.72404231e-07 4.99999997 2.72504231e-07 4.99999997 2.72604231e-07 4.99999997 2.72704231e-07 4.99999997 2.72804231e-07 4.99999997 2.72904231e-07 4.99999997 2.73004231e-07 4.99999997
+ 2.73104231e-07 4.99999997 2.73204231e-07 4.99999997 2.73304231e-07 4.99999997 2.73404231e-07 4.99999997 2.73504231e-07 4.99999997 2.73604231e-07 4.99999997 2.73704231e-07 4.99999997 2.73804231e-07 4.99999997
+ 2.73904231e-07 4.99999997 2.74004231e-07 4.99999997 2.74104231e-07 4.99999997 2.74204231e-07 4.99999997 2.74304231e-07 4.99999997 2.74404231e-07 4.99999997 2.74504231e-07 4.99999997 2.74604231e-07 4.99999997
+ 2.74704231e-07 4.99999997 2.74804231e-07 4.99999997 2.74904231e-07 4.99999997 2.75004231e-07 4.99999997 2.75104231e-07 4.99999997 2.75204231e-07 4.99999997 2.75304231e-07 4.99999997 2.75404231e-07 4.99999997
+ 2.75504231e-07 4.99999997 2.75604231e-07 4.99999997 2.75704231e-07 4.99999997 2.75804231e-07 4.99999997 2.75904231e-07 4.99999997 2.76004231e-07 4.99999997 2.76104231e-07 4.99999997 2.76204231e-07 4.99999997
+ 2.76304231e-07 4.99999997 2.76404231e-07 4.99999997 2.76504231e-07 4.99999997 2.76604231e-07 4.99999997 2.76704231e-07 4.99999997 2.76804231e-07 4.99999997 2.76904231e-07 4.99999997 2.77004231e-07 4.99999997
+ 2.77104231e-07 4.99999997 2.77204231e-07 4.99999997 2.77304231e-07 4.99999997 2.77404231e-07 4.99999997 2.77504231e-07 4.99999997 2.77604231e-07 4.99999997 2.77704231e-07 4.99999997 2.77804231e-07 4.99999997
+ 2.77904231e-07 4.99999997 2.78004231e-07 4.99999997 2.78104231e-07 4.99999997 2.78204231e-07 4.99999997 2.78304231e-07 4.99999997 2.78404231e-07 4.99999997 2.78504231e-07 4.99999997 2.78604231e-07 4.99999997
+ 2.78704231e-07 4.99999997 2.78804231e-07 4.99999997 2.78904231e-07 4.99999997 2.79004231e-07 4.99999997 2.79104231e-07 4.99999997 2.79204231e-07 4.99999997 2.79304231e-07 4.99999997 2.79404231e-07 4.99999997
+ 2.79504231e-07 4.99999997 2.79604231e-07 4.99999997 2.79704231e-07 4.99999997 2.79804231e-07 4.99999997 2.79904231e-07 4.99999997 2.80004231e-07 4.99999997 2.80104231e-07 4.99999997 2.80204231e-07 4.99999997
+ 2.80304231e-07 4.99999997 2.80404231e-07 4.99999997 2.80504231e-07 4.99999997 2.80604231e-07 4.99999997 2.80704231e-07 4.99999997 2.80804231e-07 4.99999997 2.80904231e-07 4.99999997 2.81004231e-07 4.99999997
+ 2.81104231e-07 4.99999997 2.81204231e-07 4.99999997 2.81304231e-07 4.99999997 2.81404231e-07 4.99999997 2.81504231e-07 4.99999997 2.81604231e-07 4.99999997 2.81704231e-07 4.99999997 2.81804231e-07 4.99999997
+ 2.81904231e-07 4.99999997 2.82004231e-07 4.99999997 2.82104231e-07 4.99999997 2.82204231e-07 4.99999997 2.82304231e-07 4.99999997 2.82404231e-07 4.99999997 2.82504231e-07 4.99999997 2.82604231e-07 4.99999997
+ 2.82704231e-07 4.99999997 2.82804231e-07 4.99999997 2.82904231e-07 4.99999997 2.83004231e-07 4.99999997 2.83104231e-07 4.99999997 2.83204231e-07 4.99999997 2.83304231e-07 4.99999997 2.83404231e-07 4.99999997
+ 2.83504231e-07 4.99999997 2.83604231e-07 4.99999997 2.83704231e-07 4.99999997 2.83804231e-07 4.99999997 2.83904231e-07 4.99999997 2.84004231e-07 4.99999997 2.84104231e-07 4.99999997 2.84204231e-07 4.99999997
+ 2.84304231e-07 4.99999997 2.84404231e-07 4.99999997 2.84504231e-07 4.99999997 2.84604231e-07 4.99999997 2.84704231e-07 4.99999997 2.84804231e-07 4.99999997 2.84904231e-07 4.99999997 2.85004231e-07 4.99999997
+ 2.85104231e-07 4.99999997 2.85204231e-07 4.99999997 2.85304231e-07 4.99999997 2.85404231e-07 4.99999997 2.85504231e-07 4.99999997 2.85604231e-07 4.99999997 2.85704231e-07 4.99999997 2.85804231e-07 4.99999997
+ 2.85904231e-07 4.99999997 2.86004231e-07 4.99999997 2.86104231e-07 4.99999997 2.86204231e-07 4.99999997 2.86304231e-07 4.99999997 2.86404231e-07 4.99999997 2.86504231e-07 4.99999997 2.86604231e-07 4.99999997
+ 2.86704231e-07 4.99999997 2.86804231e-07 4.99999997 2.86904231e-07 4.99999997 2.87004231e-07 4.99999997 2.87104231e-07 4.99999997 2.87204231e-07 4.99999997 2.87304231e-07 4.99999997 2.87404231e-07 4.99999997
+ 2.87504231e-07 4.99999997 2.87604231e-07 4.99999997 2.87704231e-07 4.99999997 2.87804231e-07 4.99999997 2.87904231e-07 4.99999997 2.88004231e-07 4.99999997 2.88104231e-07 4.99999997 2.88204231e-07 4.99999997
+ 2.88304231e-07 4.99999997 2.88404231e-07 4.99999997 2.88504231e-07 4.99999997 2.88604231e-07 4.99999997 2.88704231e-07 4.99999997 2.88804231e-07 4.99999997 2.88904231e-07 4.99999997 2.89004231e-07 4.99999997
+ 2.89104231e-07 4.99999997 2.89204231e-07 4.99999997 2.89304231e-07 4.99999997 2.89404231e-07 4.99999997 2.89504231e-07 4.99999997 2.89604231e-07 4.99999997 2.89704231e-07 4.99999997 2.89804231e-07 4.99999997
+ 2.89904231e-07 4.99999997 2.90004231e-07 4.99999997 2.90104231e-07 4.99999997 2.90204231e-07 4.99999997 2.90304231e-07 4.99999997 2.90404231e-07 4.99999997 2.90504231e-07 4.99999997 2.90604231e-07 4.99999997
+ 2.90704231e-07 4.99999997 2.90804231e-07 4.99999997 2.90904231e-07 4.99999997 2.91004231e-07 4.99999997 2.91104231e-07 4.99999997 2.91204231e-07 4.99999997 2.91304231e-07 4.99999997 2.91404231e-07 4.99999997
+ 2.91504231e-07 4.99999997 2.91604231e-07 4.99999997 2.91704231e-07 4.99999997 2.91804231e-07 4.99999997 2.91904231e-07 4.99999997 2.92004231e-07 4.99999997 2.92104231e-07 4.99999997 2.92204231e-07 4.99999997
+ 2.92304231e-07 4.99999997 2.92404231e-07 4.99999997 2.92504231e-07 4.99999997 2.92604231e-07 4.99999997 2.92704231e-07 4.99999997 2.92804231e-07 4.99999997 2.92904231e-07 4.99999997 2.93004231e-07 4.99999997
+ 2.93104231e-07 4.99999997 2.93204231e-07 4.99999997 2.93304231e-07 4.99999997 2.93404231e-07 4.99999997 2.93504231e-07 4.99999997 2.93604231e-07 4.99999997 2.93704231e-07 4.99999997 2.93804231e-07 4.99999997
+ 2.93904231e-07 4.99999997 2.94004231e-07 4.99999997 2.94104231e-07 4.99999997 2.94204231e-07 4.99999997 2.94304231e-07 4.99999997 2.94404231e-07 4.99999997 2.94504231e-07 4.99999997 2.94604231e-07 4.99999997
+ 2.94704231e-07 4.99999997 2.94804231e-07 4.99999997 2.94904231e-07 4.99999997 2.95004231e-07 4.99999997 2.95104231e-07 4.99999997 2.95204231e-07 4.99999997 2.95304231e-07 4.99999997 2.95404231e-07 4.99999997
+ 2.95504231e-07 4.99999997 2.95604231e-07 4.99999997 2.95704231e-07 4.99999997 2.95804231e-07 4.99999997 2.95904231e-07 4.99999997 2.96004231e-07 4.99999997 2.96104231e-07 4.99999997 2.96204231e-07 4.99999997
+ 2.96304231e-07 4.99999997 2.96404231e-07 4.99999997 2.96504231e-07 4.99999997 2.96604231e-07 4.99999997 2.96704231e-07 4.99999997 2.96804231e-07 4.99999997 2.96904231e-07 4.99999997 2.97004231e-07 4.99999997
+ 2.97104231e-07 4.99999997 2.97204231e-07 4.99999997 2.97304231e-07 4.99999997 2.97404231e-07 4.99999997 2.97504231e-07 4.99999997 2.97604231e-07 4.99999997 2.97704231e-07 4.99999997 2.97804231e-07 4.99999997
+ 2.97904231e-07 4.99999997 2.98004231e-07 4.99999997 2.98104231e-07 4.99999997 2.98204231e-07 4.99999997 2.98304231e-07 4.99999997 2.98404231e-07 4.99999997 2.98504231e-07 4.99999997 2.98604231e-07 4.99999997
+ 2.98704231e-07 4.99999997 2.98804231e-07 4.99999997 2.98904231e-07 4.99999997 2.99004231e-07 4.99999997 2.99104231e-07 4.99999997 2.99204231e-07 4.99999997 2.99304231e-07 4.99999997 2.99404231e-07 4.99999997
+ 2.99504231e-07 4.99999997 2.99604231e-07 4.99999997 2.99704231e-07 4.99999997 2.99804231e-07 4.99999997 2.99904231e-07 4.99999997 3e-07 4.99999997 3.0001e-07 4.99999997 3.0003e-07 4.99999997
+ 3.0007e-07 4.99999997 3.0015e-07 4.99999997 3.0025e-07 4.99999997 3.0035e-07 4.99999997 3.0045e-07 4.99999997 3.0055e-07 4.99999997 3.0065e-07 4.99999997 3.0075e-07 5.00000001
+ 3.0085e-07 4.99999814 3.00931988e-07 5.00001158 3.01e-07 4.99997651 3.01008484e-07 4.99997816 3.01025451e-07 4.99999556 3.01059385e-07 5.00001851 3.01090588e-07 5.00001181 3.01143428e-07 5.00000049
+ 3.011991e-07 5.00001369 3.012991e-07 4.99978337 3.013991e-07 5.00014046 3.014991e-07 5.00032641 3.01578678e-07 4.99987228 3.01663998e-07 4.99960593 3.01763998e-07 5.00049059 3.01858547e-07 4.99953494
+ 3.01958547e-07 5.000381 3.02058547e-07 4.99971267 3.02158547e-07 5.00020063 3.02258547e-07 4.99986803 3.02358547e-07 5.00007856 3.02458547e-07 4.99995925 3.02558547e-07 5.00001358 3.02658547e-07 5.00000443
+ 3.02758547e-07 4.99998371 3.02858547e-07 5.00002377 3.02958547e-07 4.99997188 3.03058547e-07 5.0000303 3.03158547e-07 4.99996886 3.03258547e-07 5.00003095 3.03358547e-07 4.99996972 3.03458547e-07 5.00002911
+ 3.03558547e-07 4.99997213 3.03658547e-07 5.00002639 3.03758547e-07 4.99997499 3.03858547e-07 5.0000235 3.03958547e-07 4.99997783 3.04058547e-07 5.00002075 3.04158547e-07 4.99998047 3.04258547e-07 5.00001824
+ 3.04358547e-07 4.99998284 3.04458547e-07 5.000016 3.04558547e-07 4.99998495 3.04658547e-07 5.00001403 3.04758547e-07 4.99998681 3.04858547e-07 5.00001229 3.04958547e-07 4.99998843 3.05058547e-07 5.00001077
+ 3.05158547e-07 4.99998986 3.05258547e-07 5.00000943 3.05358547e-07 4.99999111 3.05458547e-07 5.00000826 3.05558547e-07 4.99999221 3.05658547e-07 5.00000724 3.05758547e-07 4.99999317 3.05858547e-07 5.00000634
+ 3.05958547e-07 4.99999401 3.06058547e-07 5.00000555 3.06158547e-07 4.99999474 3.06258547e-07 5.00000486 3.06358547e-07 4.99999539 3.06458547e-07 5.00000426 3.06558547e-07 4.99999595 3.06658547e-07 5.00000373
+ 3.06758547e-07 4.99999645 3.06858547e-07 5.00000327 3.06958547e-07 4.99999688 3.07058547e-07 5.00000286 3.07158547e-07 4.99999727 3.07258547e-07 5.00000251 3.07358547e-07 4.9999976 3.07458547e-07 5.00000219
+ 3.07558547e-07 4.99999789 3.07658547e-07 5.00000192 3.07758547e-07 4.99999815 3.07858547e-07 5.00000168 3.07958547e-07 4.99999837 3.08058547e-07 5.00000147 3.08158547e-07 4.99999857 3.08258547e-07 5.00000128
+ 3.08358547e-07 4.99999874 3.08458547e-07 5.00000112 3.08558547e-07 4.99999889 3.08658547e-07 5.00000098 3.08758547e-07 4.99999903 3.08858547e-07 5.00000086 3.08958547e-07 4.99999914 3.09058547e-07 5.00000075
+ 3.09158547e-07 4.99999925 3.09258547e-07 5.00000065 3.09358547e-07 4.99999934 3.09458547e-07 5.00000057 3.09558547e-07 4.99999941 3.09658547e-07 5.00000049 3.09758547e-07 4.99999948 3.09858547e-07 5.00000043
+ 3.09958547e-07 4.99999954 3.10058547e-07 5.00000037 3.10158547e-07 4.9999996 3.10258547e-07 5.00000032 3.10358547e-07 4.99999964 3.10458547e-07 5.00000028 3.10558547e-07 4.99999968 3.10658547e-07 5.00000024
+ 3.10758547e-07 4.99999972 3.10858547e-07 5.00000021 3.10958547e-07 4.99999975 3.11058547e-07 5.00000018 3.11158547e-07 4.99999977 3.11258547e-07 5.00000015 3.11358547e-07 4.9999998 3.11458547e-07 5.00000013
+ 3.11558547e-07 4.99999982 3.11658547e-07 5.00000011 3.11758547e-07 4.99999984 3.11858547e-07 5.00000009 3.11958547e-07 4.99999986 3.12058547e-07 5.00000008 3.12158547e-07 4.99999987 3.12258547e-07 5.00000006
+ 3.12358547e-07 4.99999988 3.12458547e-07 5.00000005 3.12558547e-07 4.99999989 3.12658547e-07 5.00000004 3.12758547e-07 4.9999999 3.12858547e-07 5.00000003 3.12958547e-07 4.99999991 3.13058547e-07 5.00000003
+ 3.13158547e-07 4.99999992 3.13258547e-07 5.00000002 3.13358547e-07 4.99999993 3.13458547e-07 5.00000001 3.13558547e-07 4.99999993 3.13658547e-07 5.00000001 3.13758547e-07 4.99999994 3.13858547e-07 5.0
+ 3.13958547e-07 4.99999994 3.14058547e-07 5.0 3.14158547e-07 4.99999995 3.14258547e-07 5.0 3.14358547e-07 4.99999995 3.14458547e-07 4.99999999 3.14558547e-07 4.99999995 3.14658547e-07 4.99999999
+ 3.14758547e-07 4.99999995 3.14858547e-07 4.99999999 3.14958547e-07 4.99999996 3.15058547e-07 4.99999999 3.15158547e-07 4.99999996 3.15258547e-07 4.99999998 3.15358547e-07 4.99999996 3.15458547e-07 4.99999998
+ 3.15558547e-07 4.99999996 3.15658547e-07 4.99999998 3.15758547e-07 4.99999996 3.15858547e-07 4.99999998 3.15958547e-07 4.99999996 3.16058547e-07 4.99999998 3.16158547e-07 4.99999997 3.16258547e-07 4.99999998
+ 3.16358547e-07 4.99999997 3.16458547e-07 4.99999998 3.16558547e-07 4.99999997 3.16658547e-07 4.99999998 3.16758547e-07 4.99999997 3.16858547e-07 4.99999998 3.16958547e-07 4.99999997 3.17058547e-07 4.99999998
+ 3.17158547e-07 4.99999997 3.17258547e-07 4.99999998 3.17358547e-07 4.99999997 3.17458547e-07 4.99999998 3.17558547e-07 4.99999997 3.17658547e-07 4.99999997 3.17758547e-07 4.99999997 3.17858547e-07 4.99999997
+ 3.17958547e-07 4.99999997 3.18058547e-07 4.99999997 3.18158547e-07 4.99999997 3.18258547e-07 4.99999997 3.18358547e-07 4.99999997 3.18458547e-07 4.99999997 3.18558547e-07 4.99999997 3.18658547e-07 4.99999997
+ 3.18758547e-07 4.99999997 3.18858547e-07 4.99999997 3.18958547e-07 4.99999997 3.19058547e-07 4.99999997 3.19158547e-07 4.99999997 3.19258547e-07 4.99999997 3.19358547e-07 4.99999997 3.19458547e-07 4.99999997
+ 3.19558547e-07 4.99999997 3.19658547e-07 4.99999997 3.19758547e-07 4.99999997 3.19858547e-07 4.99999997 3.19958547e-07 4.99999997 3.20058547e-07 4.99999997 3.20158547e-07 4.99999997 3.20258547e-07 4.99999997
+ 3.20358547e-07 4.99999997 3.20458547e-07 4.99999997 3.20558547e-07 4.99999997 3.20658547e-07 4.99999997 3.20758547e-07 4.99999997 3.20858547e-07 4.99999997 3.20958547e-07 4.99999997 3.21058547e-07 4.99999997
+ 3.21158547e-07 4.99999997 3.21258547e-07 4.99999997 3.21358547e-07 4.99999997 3.21458547e-07 4.99999997 3.21558547e-07 4.99999997 3.21658547e-07 4.99999997 3.21758547e-07 4.99999997 3.21858547e-07 4.99999997
+ 3.21958547e-07 4.99999997 3.22058547e-07 4.99999997 3.22158547e-07 4.99999997 3.22258547e-07 4.99999997 3.22358547e-07 4.99999997 3.22458547e-07 4.99999997 3.22558547e-07 4.99999997 3.22658547e-07 4.99999997
+ 3.22758547e-07 4.99999997 3.22858547e-07 4.99999997 3.22958547e-07 4.99999997 3.23058547e-07 4.99999997 3.23158547e-07 4.99999997 3.23258547e-07 4.99999997 3.23358547e-07 4.99999997 3.23458547e-07 4.99999997
+ 3.23558547e-07 4.99999997 3.23658547e-07 4.99999997 3.23758547e-07 4.99999997 3.23858547e-07 4.99999997 3.23958547e-07 4.99999997 3.24058547e-07 4.99999997 3.24158547e-07 4.99999997 3.24258547e-07 4.99999997
+ 3.24358547e-07 4.99999997 3.24458547e-07 4.99999997 3.24558547e-07 4.99999997 3.24658547e-07 4.99999997 3.24758547e-07 4.99999997 3.24858547e-07 4.99999997 3.24958547e-07 4.99999997 3.25058547e-07 4.99999997
+ 3.25158547e-07 4.99999997 3.25258547e-07 4.99999997 3.25358547e-07 4.99999997 3.25458547e-07 4.99999997 3.25558547e-07 4.99999997 3.25658547e-07 4.99999997 3.25758547e-07 4.99999997 3.25858547e-07 4.99999997
+ 3.25958547e-07 4.99999997 3.26058547e-07 4.99999997 3.26158547e-07 4.99999997 3.26258547e-07 4.99999997 3.26358547e-07 4.99999997 3.26458547e-07 4.99999997 3.26558547e-07 4.99999997 3.26658547e-07 4.99999997
+ 3.26758547e-07 4.99999997 3.26858547e-07 4.99999997 3.26958547e-07 4.99999997 3.27058547e-07 4.99999997 3.27158547e-07 4.99999997 3.27258547e-07 4.99999997 3.27358547e-07 4.99999997 3.27458547e-07 4.99999997
+ 3.27558547e-07 4.99999997 3.27658547e-07 4.99999997 3.27758547e-07 4.99999997 3.27858547e-07 4.99999997 3.27958547e-07 4.99999997 3.28058547e-07 4.99999997 3.28158547e-07 4.99999997 3.28258547e-07 4.99999997
+ 3.28358547e-07 4.99999997 3.28458547e-07 4.99999997 3.28558547e-07 4.99999997 3.28658547e-07 4.99999997 3.28758547e-07 4.99999997 3.28858547e-07 4.99999997 3.28958547e-07 4.99999997 3.29058547e-07 4.99999997
+ 3.29158547e-07 4.99999997 3.29258547e-07 4.99999997 3.29358547e-07 4.99999997 3.29458547e-07 4.99999997 3.29558547e-07 4.99999997 3.29658547e-07 4.99999997 3.29758547e-07 4.99999997 3.29858547e-07 4.99999997
+ 3.29958547e-07 4.99999997 3.30058547e-07 4.99999997 3.30158547e-07 4.99999997 3.30258547e-07 4.99999997 3.30358547e-07 4.99999997 3.30458547e-07 4.99999997 3.30558547e-07 4.99999997 3.30658547e-07 4.99999997
+ 3.30758547e-07 4.99999997 3.30858547e-07 4.99999997 3.30958547e-07 4.99999997 3.31058547e-07 4.99999997 3.31158547e-07 4.99999997 3.31258547e-07 4.99999997 3.31358547e-07 4.99999997 3.31458547e-07 4.99999997
+ 3.31558547e-07 4.99999997 3.31658547e-07 4.99999997 3.31758547e-07 4.99999997 3.31858547e-07 4.99999997 3.31958547e-07 4.99999997 3.32058547e-07 4.99999997 3.32158547e-07 4.99999997 3.32258547e-07 4.99999997
+ 3.32358547e-07 4.99999997 3.32458547e-07 4.99999997 3.32558547e-07 4.99999997 3.32658547e-07 4.99999997 3.32758547e-07 4.99999997 3.32858547e-07 4.99999997 3.32958547e-07 4.99999997 3.33058547e-07 4.99999997
+ 3.33158547e-07 4.99999997 3.33258547e-07 4.99999997 3.33358547e-07 4.99999997 3.33458547e-07 4.99999997 3.33558547e-07 4.99999997 3.33658547e-07 4.99999997 3.33758547e-07 4.99999997 3.33858547e-07 4.99999997
+ 3.33958547e-07 4.99999997 3.34058547e-07 4.99999997 3.34158547e-07 4.99999997 3.34258547e-07 4.99999997 3.34358547e-07 4.99999997 3.34458547e-07 4.99999997 3.34558547e-07 4.99999997 3.34658547e-07 4.99999997
+ 3.34758547e-07 4.99999997 3.34858547e-07 4.99999997 3.34958547e-07 4.99999997 3.35058547e-07 4.99999997 3.35158547e-07 4.99999997 3.35258547e-07 4.99999997 3.35358547e-07 4.99999997 3.35458547e-07 4.99999997
+ 3.35558547e-07 4.99999997 3.35658547e-07 4.99999997 3.35758547e-07 4.99999997 3.35858547e-07 4.99999997 3.35958547e-07 4.99999997 3.36058547e-07 4.99999997 3.36158547e-07 4.99999997 3.36258547e-07 4.99999997
+ 3.36358547e-07 4.99999997 3.36458547e-07 4.99999997 3.36558547e-07 4.99999997 3.36658547e-07 4.99999997 3.36758547e-07 4.99999997 3.36858547e-07 4.99999997 3.36958547e-07 4.99999997 3.37058547e-07 4.99999997
+ 3.37158547e-07 4.99999997 3.37258547e-07 4.99999997 3.37358547e-07 4.99999997 3.37458547e-07 4.99999997 3.37558547e-07 4.99999997 3.37658547e-07 4.99999997 3.37758547e-07 4.99999997 3.37858547e-07 4.99999997
+ 3.37958547e-07 4.99999997 3.38058547e-07 4.99999997 3.38158547e-07 4.99999997 3.38258547e-07 4.99999997 3.38358547e-07 4.99999997 3.38458547e-07 4.99999997 3.38558547e-07 4.99999997 3.38658547e-07 4.99999997
+ 3.38758547e-07 4.99999997 3.38858547e-07 4.99999997 3.38958547e-07 4.99999997 3.39058547e-07 4.99999997 3.39158547e-07 4.99999997 3.39258547e-07 4.99999997 3.39358547e-07 4.99999997 3.39458547e-07 4.99999997
+ 3.39558547e-07 4.99999997 3.39658547e-07 4.99999997 3.39758547e-07 4.99999997 3.39858547e-07 4.99999997 3.39958547e-07 4.99999997 3.40058547e-07 4.99999997 3.40158547e-07 4.99999997 3.40258547e-07 4.99999997
+ 3.40358547e-07 4.99999997 3.40458547e-07 4.99999997 3.40558547e-07 4.99999997 3.40658547e-07 4.99999997 3.40758547e-07 4.99999997 3.40858547e-07 4.99999997 3.40958547e-07 4.99999997 3.41058547e-07 4.99999997
+ 3.41158547e-07 4.99999997 3.41258547e-07 4.99999997 3.41358547e-07 4.99999997 3.41458547e-07 4.99999997 3.41558547e-07 4.99999997 3.41658547e-07 4.99999997 3.41758547e-07 4.99999997 3.41858547e-07 4.99999997
+ 3.41958547e-07 4.99999997 3.42058547e-07 4.99999997 3.42158547e-07 4.99999997 3.42258547e-07 4.99999997 3.42358547e-07 4.99999997 3.42458547e-07 4.99999997 3.42558547e-07 4.99999997 3.42658547e-07 4.99999997
+ 3.42758547e-07 4.99999997 3.42858547e-07 4.99999997 3.42958547e-07 4.99999997 3.43058547e-07 4.99999997 3.43158547e-07 4.99999997 3.43258547e-07 4.99999997 3.43358547e-07 4.99999997 3.43458547e-07 4.99999997
+ 3.43558547e-07 4.99999997 3.43658547e-07 4.99999997 3.43758547e-07 4.99999997 3.43858547e-07 4.99999997 3.43958547e-07 4.99999997 3.44058547e-07 4.99999997 3.44158547e-07 4.99999997 3.44258547e-07 4.99999997
+ 3.44358547e-07 4.99999997 3.44458547e-07 4.99999997 3.44558547e-07 4.99999997 3.44658547e-07 4.99999997 3.44758547e-07 4.99999997 3.44858547e-07 4.99999997 3.44958547e-07 4.99999997 3.45058547e-07 4.99999997
+ 3.45158547e-07 4.99999997 3.45258547e-07 4.99999997 3.45358547e-07 4.99999997 3.45458547e-07 4.99999997 3.45558547e-07 4.99999997 3.45658547e-07 4.99999997 3.45758547e-07 4.99999997 3.45858547e-07 4.99999997
+ 3.45958547e-07 4.99999997 3.46058547e-07 4.99999997 3.46158547e-07 4.99999997 3.46258547e-07 4.99999997 3.46358547e-07 4.99999997 3.46458547e-07 4.99999997 3.46558547e-07 4.99999997 3.46658547e-07 4.99999997
+ 3.46758547e-07 4.99999997 3.46858547e-07 4.99999997 3.46958547e-07 4.99999997 3.47058547e-07 4.99999997 3.47158547e-07 4.99999997 3.47258547e-07 4.99999997 3.47358547e-07 4.99999997 3.47458547e-07 4.99999997
+ 3.47558547e-07 4.99999997 3.47658547e-07 4.99999997 3.47758547e-07 4.99999997 3.47858547e-07 4.99999997 3.47958547e-07 4.99999997 3.48058547e-07 4.99999997 3.48158547e-07 4.99999997 3.48258547e-07 4.99999997
+ 3.48358547e-07 4.99999997 3.48458547e-07 4.99999997 3.48558547e-07 4.99999997 3.48658547e-07 4.99999997 3.48758547e-07 4.99999997 3.48858547e-07 4.99999997 3.48958547e-07 4.99999997 3.49058547e-07 4.99999997
+ 3.49158547e-07 4.99999997 3.49258547e-07 4.99999997 3.49358547e-07 4.99999997 3.49458547e-07 4.99999997 3.49558547e-07 4.99999997 3.49658547e-07 4.99999997 3.49758547e-07 4.99999997 3.49858547e-07 4.99999997
+ 3.49958547e-07 4.99999997 3.50058547e-07 4.99999997 3.50158547e-07 4.99999997 3.50258547e-07 4.99999997 3.50358547e-07 4.99999997 3.50458547e-07 4.99999997 3.50558547e-07 4.99999997 3.50658547e-07 4.99999997
+ 3.50758547e-07 4.99999997 3.50858547e-07 4.99999997 3.50958547e-07 4.99999997 3.51e-07 4.99999997 3.5101e-07 4.99999997 3.5103e-07 4.99999997 3.5107e-07 4.99999997 3.5115e-07 4.99999997
+ 3.5125e-07 4.99999997 3.5135e-07 4.99999997 3.5145e-07 4.99999997 3.5155e-07 4.99999997 3.5165e-07 4.99999997 3.5175e-07 4.99999997 3.5185e-07 4.99999997 3.51930828e-07 5.00000123
+ 3.52e-07 5.00000148 3.52008608e-07 4.99998858 3.52025825e-07 4.99996426 3.52060258e-07 5.00000424 3.52106188e-07 5.00004614 3.52150118e-07 4.99998884 3.5219811e-07 4.99996906 3.522555e-07 5.0000164
+ 3.52312176e-07 4.99999727 3.52404431e-07 5.00000287 3.52490759e-07 4.99999775 3.52590759e-07 5.0000011 3.52690759e-07 4.99999973 3.52790759e-07 4.99999956 3.52890759e-07 5.00000078 3.52990759e-07 4.99999897
+ 3.53090759e-07 5.00000104 3.53190759e-07 4.99999892 3.53290759e-07 5.00000096 3.53390759e-07 4.99999906 3.53490759e-07 5.00000079 3.53590759e-07 4.99999924 3.53690759e-07 5.00000062 3.53790759e-07 4.99999939
+ 3.53890759e-07 5.00000049 3.53990759e-07 4.99999951 3.54090759e-07 5.00000038 3.54190759e-07 4.9999996 3.54290759e-07 5.00000031 3.54390759e-07 4.99999966 3.54490759e-07 5.00000025 3.54590759e-07 4.99999971
+ 3.54690759e-07 5.00000021 3.54790759e-07 4.99999975 3.54890759e-07 5.00000018 3.54990759e-07 4.99999978 3.55090759e-07 5.00000015 3.55190759e-07 4.9999998 3.55290759e-07 5.00000013 3.55390759e-07 4.99999983
+ 3.55490759e-07 5.00000011 3.55590759e-07 4.99999984 3.55690759e-07 5.00000009 3.55790759e-07 4.99999986 3.55890759e-07 5.00000008 3.55990759e-07 4.99999987 3.56090759e-07 5.00000007 3.56190759e-07 4.99999988
+ 3.56290759e-07 5.00000006 3.56390759e-07 4.99999989 3.56490759e-07 5.00000005 3.56590759e-07 4.9999999 3.56690759e-07 5.00000004 3.56790759e-07 4.99999991 3.56890759e-07 5.00000003 3.56990759e-07 4.99999992
+ 3.57090759e-07 5.00000002 3.57190759e-07 4.99999992 3.57290759e-07 5.00000001 3.57390759e-07 4.99999993 3.57490759e-07 5.00000001 3.57590759e-07 4.99999994 3.57690759e-07 5.00000001 3.57790759e-07 4.99999994
+ 3.57890759e-07 5.0 3.57990759e-07 4.99999994 3.58090759e-07 5.0 3.58190759e-07 4.99999995 3.58290759e-07 4.99999999 3.58390759e-07 4.99999995 3.58490759e-07 4.99999999 3.58590759e-07 4.99999995
+ 3.58690759e-07 4.99999999 3.58790759e-07 4.99999996 3.58890759e-07 4.99999999 3.58990759e-07 4.99999996 3.59090759e-07 4.99999999 3.59190759e-07 4.99999996 3.59290759e-07 4.99999998 3.59390759e-07 4.99999996
+ 3.59490759e-07 4.99999998 3.59590759e-07 4.99999996 3.59690759e-07 4.99999998 3.59790759e-07 4.99999996 3.59890759e-07 4.99999998 3.59990759e-07 4.99999996 3.60090759e-07 4.99999998 3.60190759e-07 4.99999997
+ 3.60290759e-07 4.99999998 3.60390759e-07 4.99999997 3.60490759e-07 4.99999998 3.60590759e-07 4.99999997 3.60690759e-07 4.99999998 3.60790759e-07 4.99999997 3.60890759e-07 4.99999998 3.60990759e-07 4.99999997
+ 3.61090759e-07 4.99999998 3.61190759e-07 4.99999997 3.61290759e-07 4.99999998 3.61390759e-07 4.99999997 3.61490759e-07 4.99999997 3.61590759e-07 4.99999997 3.61690759e-07 4.99999997 3.61790759e-07 4.99999997
+ 3.61890759e-07 4.99999997 3.61990759e-07 4.99999997 3.62090759e-07 4.99999997 3.62190759e-07 4.99999997 3.62290759e-07 4.99999997 3.62390759e-07 4.99999997 3.62490759e-07 4.99999997 3.62590759e-07 4.99999997
+ 3.62690759e-07 4.99999997 3.62790759e-07 4.99999997 3.62890759e-07 4.99999997 3.62990759e-07 4.99999997 3.63090759e-07 4.99999997 3.63190759e-07 4.99999997 3.63290759e-07 4.99999997 3.63390759e-07 4.99999997
+ 3.63490759e-07 4.99999997 3.63590759e-07 4.99999997 3.63690759e-07 4.99999997 3.63790759e-07 4.99999997 3.63890759e-07 4.99999997 3.63990759e-07 4.99999997 3.64090759e-07 4.99999997 3.64190759e-07 4.99999997
+ 3.64290759e-07 4.99999997 3.64390759e-07 4.99999997 3.64490759e-07 4.99999997 3.64590759e-07 4.99999997 3.64690759e-07 4.99999997 3.64790759e-07 4.99999997 3.64890759e-07 4.99999997 3.64990759e-07 4.99999997
+ 3.65090759e-07 4.99999997 3.65190759e-07 4.99999997 3.65290759e-07 4.99999997 3.65390759e-07 4.99999997 3.65490759e-07 4.99999997 3.65590759e-07 4.99999997 3.65690759e-07 4.99999997 3.65790759e-07 4.99999997
+ 3.65890759e-07 4.99999997 3.65990759e-07 4.99999997 3.66090759e-07 4.99999997 3.66190759e-07 4.99999997 3.66290759e-07 4.99999997 3.66390759e-07 4.99999997 3.66490759e-07 4.99999997 3.66590759e-07 4.99999997
+ 3.66690759e-07 4.99999997 3.66790759e-07 4.99999997 3.66890759e-07 4.99999997 3.66990759e-07 4.99999997 3.67090759e-07 4.99999997 3.67190759e-07 4.99999997 3.67290759e-07 4.99999997 3.67390759e-07 4.99999997
+ 3.67490759e-07 4.99999997 3.67590759e-07 4.99999997 3.67690759e-07 4.99999997 3.67790759e-07 4.99999997 3.67890759e-07 4.99999997 3.67990759e-07 4.99999997 3.68090759e-07 4.99999997 3.68190759e-07 4.99999997
+ 3.68290759e-07 4.99999997 3.68390759e-07 4.99999997 3.68490759e-07 4.99999997 3.68590759e-07 4.99999997 3.68690759e-07 4.99999997 3.68790759e-07 4.99999997 3.68890759e-07 4.99999997 3.68990759e-07 4.99999997
+ 3.69090759e-07 4.99999997 3.69190759e-07 4.99999997 3.69290759e-07 4.99999997 3.69390759e-07 4.99999997 3.69490759e-07 4.99999997 3.69590759e-07 4.99999997 3.69690759e-07 4.99999997 3.69790759e-07 4.99999997
+ 3.69890759e-07 4.99999997 3.69990759e-07 4.99999997 3.70090759e-07 4.99999997 3.70190759e-07 4.99999997 3.70290759e-07 4.99999997 3.70390759e-07 4.99999997 3.70490759e-07 4.99999997 3.70590759e-07 4.99999997
+ 3.70690759e-07 4.99999997 3.70790759e-07 4.99999997 3.70890759e-07 4.99999997 3.70990759e-07 4.99999997 3.71090759e-07 4.99999997 3.71190759e-07 4.99999997 3.71290759e-07 4.99999997 3.71390759e-07 4.99999997
+ 3.71490759e-07 4.99999997 3.71590759e-07 4.99999997 3.71690759e-07 4.99999997 3.71790759e-07 4.99999997 3.71890759e-07 4.99999997 3.71990759e-07 4.99999997 3.72090759e-07 4.99999997 3.72190759e-07 4.99999997
+ 3.72290759e-07 4.99999997 3.72390759e-07 4.99999997 3.72490759e-07 4.99999997 3.72590759e-07 4.99999997 3.72690759e-07 4.99999997 3.72790759e-07 4.99999997 3.72890759e-07 4.99999997 3.72990759e-07 4.99999997
+ 3.73090759e-07 4.99999997 3.73190759e-07 4.99999997 3.73290759e-07 4.99999997 3.73390759e-07 4.99999997 3.73490759e-07 4.99999997 3.73590759e-07 4.99999997 3.73690759e-07 4.99999997 3.73790759e-07 4.99999997
+ 3.73890759e-07 4.99999997 3.73990759e-07 4.99999997 3.74090759e-07 4.99999997 3.74190759e-07 4.99999997 3.74290759e-07 4.99999997 3.74390759e-07 4.99999997 3.74490759e-07 4.99999997 3.74590759e-07 4.99999997
+ 3.74690759e-07 4.99999997 3.74790759e-07 4.99999997 3.74890759e-07 4.99999997 3.74990759e-07 4.99999997 3.75090759e-07 4.99999997 3.75190759e-07 4.99999997 3.75290759e-07 4.99999997 3.75390759e-07 4.99999997
+ 3.75490759e-07 4.99999997 3.75590759e-07 4.99999997 3.75690759e-07 4.99999997 3.75790759e-07 4.99999997 3.75890759e-07 4.99999997 3.75990759e-07 4.99999997 3.76090759e-07 4.99999997 3.76190759e-07 4.99999997
+ 3.76290759e-07 4.99999997 3.76390759e-07 4.99999997 3.76490759e-07 4.99999997 3.76590759e-07 4.99999997 3.76690759e-07 4.99999997 3.76790759e-07 4.99999997 3.76890759e-07 4.99999997 3.76990759e-07 4.99999997
+ 3.77090759e-07 4.99999997 3.77190759e-07 4.99999997 3.77290759e-07 4.99999997 3.77390759e-07 4.99999997 3.77490759e-07 4.99999997 3.77590759e-07 4.99999997 3.77690759e-07 4.99999997 3.77790759e-07 4.99999997
+ 3.77890759e-07 4.99999997 3.77990759e-07 4.99999997 3.78090759e-07 4.99999997 3.78190759e-07 4.99999997 3.78290759e-07 4.99999997 3.78390759e-07 4.99999997 3.78490759e-07 4.99999997 3.78590759e-07 4.99999997
+ 3.78690759e-07 4.99999997 3.78790759e-07 4.99999997 3.78890759e-07 4.99999997 3.78990759e-07 4.99999997 3.79090759e-07 4.99999997 3.79190759e-07 4.99999997 3.79290759e-07 4.99999997 3.79390759e-07 4.99999997
+ 3.79490759e-07 4.99999997 3.79590759e-07 4.99999997 3.79690759e-07 4.99999997 3.79790759e-07 4.99999997 3.79890759e-07 4.99999997 3.79990759e-07 4.99999997 3.80090759e-07 4.99999997 3.80190759e-07 4.99999997
+ 3.80290759e-07 4.99999997 3.80390759e-07 4.99999997 3.80490759e-07 4.99999997 3.80590759e-07 4.99999997 3.80690759e-07 4.99999997 3.80790759e-07 4.99999997 3.80890759e-07 4.99999997 3.80990759e-07 4.99999997
+ 3.81090759e-07 4.99999997 3.81190759e-07 4.99999997 3.81290759e-07 4.99999997 3.81390759e-07 4.99999997 3.81490759e-07 4.99999997 3.81590759e-07 4.99999997 3.81690759e-07 4.99999997 3.81790759e-07 4.99999997
+ 3.81890759e-07 4.99999997 3.81990759e-07 4.99999997 3.82090759e-07 4.99999997 3.82190759e-07 4.99999997 3.82290759e-07 4.99999997 3.82390759e-07 4.99999997 3.82490759e-07 4.99999997 3.82590759e-07 4.99999997
+ 3.82690759e-07 4.99999997 3.82790759e-07 4.99999997 3.82890759e-07 4.99999997 3.82990759e-07 4.99999997 3.83090759e-07 4.99999997 3.83190759e-07 4.99999997 3.83290759e-07 4.99999997 3.83390759e-07 4.99999997
+ 3.83490759e-07 4.99999997 3.83590759e-07 4.99999997 3.83690759e-07 4.99999997 3.83790759e-07 4.99999997 3.83890759e-07 4.99999997 3.83990759e-07 4.99999997 3.84090759e-07 4.99999997 3.84190759e-07 4.99999997
+ 3.84290759e-07 4.99999997 3.84390759e-07 4.99999997 3.84490759e-07 4.99999997 3.84590759e-07 4.99999997 3.84690759e-07 4.99999997 3.84790759e-07 4.99999997 3.84890759e-07 4.99999997 3.84990759e-07 4.99999997
+ 3.85090759e-07 4.99999997 3.85190759e-07 4.99999997 3.85290759e-07 4.99999997 3.85390759e-07 4.99999997 3.85490759e-07 4.99999997 3.85590759e-07 4.99999997 3.85690759e-07 4.99999997 3.85790759e-07 4.99999997
+ 3.85890759e-07 4.99999997 3.85990759e-07 4.99999997 3.86090759e-07 4.99999997 3.86190759e-07 4.99999997 3.86290759e-07 4.99999997 3.86390759e-07 4.99999997 3.86490759e-07 4.99999997 3.86590759e-07 4.99999997
+ 3.86690759e-07 4.99999997 3.86790759e-07 4.99999997 3.86890759e-07 4.99999997 3.86990759e-07 4.99999997 3.87090759e-07 4.99999997 3.87190759e-07 4.99999997 3.87290759e-07 4.99999997 3.87390759e-07 4.99999997
+ 3.87490759e-07 4.99999997 3.87590759e-07 4.99999997 3.87690759e-07 4.99999997 3.87790759e-07 4.99999997 3.87890759e-07 4.99999997 3.87990759e-07 4.99999997 3.88090759e-07 4.99999997 3.88190759e-07 4.99999997
+ 3.88290759e-07 4.99999997 3.88390759e-07 4.99999997 3.88490759e-07 4.99999997 3.88590759e-07 4.99999997 3.88690759e-07 4.99999997 3.88790759e-07 4.99999997 3.88890759e-07 4.99999997 3.88990759e-07 4.99999997
+ 3.89090759e-07 4.99999997 3.89190759e-07 4.99999997 3.89290759e-07 4.99999997 3.89390759e-07 4.99999997 3.89490759e-07 4.99999997 3.89590759e-07 4.99999997 3.89690759e-07 4.99999997 3.89790759e-07 4.99999997
+ 3.89890759e-07 4.99999997 3.89990759e-07 4.99999997 3.90090759e-07 4.99999997 3.90190759e-07 4.99999997 3.90290759e-07 4.99999997 3.90390759e-07 4.99999997 3.90490759e-07 4.99999997 3.90590759e-07 4.99999997
+ 3.90690759e-07 4.99999997 3.90790759e-07 4.99999997 3.90890759e-07 4.99999997 3.90990759e-07 4.99999997 3.91090759e-07 4.99999997 3.91190759e-07 4.99999997 3.91290759e-07 4.99999997 3.91390759e-07 4.99999997
+ 3.91490759e-07 4.99999997 3.91590759e-07 4.99999997 3.91690759e-07 4.99999997 3.91790759e-07 4.99999997 3.91890759e-07 4.99999997 3.91990759e-07 4.99999997 3.92090759e-07 4.99999997 3.92190759e-07 4.99999997
+ 3.92290759e-07 4.99999997 3.92390759e-07 4.99999997 3.92490759e-07 4.99999997 3.92590759e-07 4.99999997 3.92690759e-07 4.99999997 3.92790759e-07 4.99999997 3.92890759e-07 4.99999997 3.92990759e-07 4.99999997
+ 3.93090759e-07 4.99999997 3.93190759e-07 4.99999997 3.93290759e-07 4.99999997 3.93390759e-07 4.99999997 3.93490759e-07 4.99999997 3.93590759e-07 4.99999997 3.93690759e-07 4.99999997 3.93790759e-07 4.99999997
+ 3.93890759e-07 4.99999997 3.93990759e-07 4.99999997 3.94090759e-07 4.99999997 3.94190759e-07 4.99999997 3.94290759e-07 4.99999997 3.94390759e-07 4.99999997 3.94490759e-07 4.99999997 3.94590759e-07 4.99999997
+ 3.94690759e-07 4.99999997 3.94790759e-07 4.99999997 3.94890759e-07 4.99999997 3.94990759e-07 4.99999997 3.95090759e-07 4.99999997 3.95190759e-07 4.99999997 3.95290759e-07 4.99999997 3.95390759e-07 4.99999997
+ 3.95490759e-07 4.99999997 3.95590759e-07 4.99999997 3.95690759e-07 4.99999997 3.95790759e-07 4.99999997 3.95890759e-07 4.99999997 3.95990759e-07 4.99999997 3.96090759e-07 4.99999997 3.96190759e-07 4.99999997
+ 3.96290759e-07 4.99999997 3.96390759e-07 4.99999997 3.96490759e-07 4.99999997 3.96590759e-07 4.99999997 3.96690759e-07 4.99999997 3.96790759e-07 4.99999997 3.96890759e-07 4.99999997 3.96990759e-07 4.99999997
+ 3.97090759e-07 4.99999997 3.97190759e-07 4.99999997 3.97290759e-07 4.99999997 3.97390759e-07 4.99999997 3.97490759e-07 4.99999997 3.97590759e-07 4.99999997 3.97690759e-07 4.99999997 3.97790759e-07 4.99999997
+ 3.97890759e-07 4.99999997 3.97990759e-07 4.99999997 3.98090759e-07 4.99999997 3.98190759e-07 4.99999997 3.98290759e-07 4.99999997 3.98390759e-07 4.99999997 3.98490759e-07 4.99999997 3.98590759e-07 4.99999997
+ 3.98690759e-07 4.99999997 3.98790759e-07 4.99999997 3.98890759e-07 4.99999997 3.98990759e-07 4.99999997 3.99090759e-07 4.99999997 3.99190759e-07 4.99999997 3.99290759e-07 4.99999997 3.99390759e-07 4.99999997
+ 3.99490759e-07 4.99999997 3.99590759e-07 4.99999997 3.99690759e-07 4.99999997 3.99790759e-07 4.99999997 3.99890759e-07 4.99999997 3.99990759e-07 4.99999997 4e-07 4.99999997 4.0001e-07 4.99999997
+ 4.0003e-07 4.99999997 4.0007e-07 4.99999997 4.0015e-07 4.99999997 4.0025e-07 4.99999997 4.0035e-07 4.99999997 4.0045e-07 4.99999997 4.0055e-07 4.99999997 4.0065e-07 4.99999997
+ 4.0075e-07 5.00000001 4.0085e-07 4.99999686 4.00931913e-07 5.00000385 4.01e-07 5.00010633 4.01008477e-07 5.00014453 4.01025432e-07 5.00027393 4.01059342e-07 4.99937073 4.01090545e-07 4.99743534
+ 4.01143412e-07 4.99875515 4.01199108e-07 5.05834962 4.01266691e-07 4.82390127 4.01329415e-07 1.08191107 4.01394829e-07 -0.0834648083 4.01464618e-07 0.122803197 4.01533535e-07 -0.0865031891 4.01610366e-07 0.0799022498
+ 4.01709241e-07 -0.071357353 4.01809241e-07 0.0656628381 4.01909241e-07 -0.0593137472 4.02009241e-07 0.0545273436 4.02109241e-07 -0.0493042956 4.02209241e-07 0.0453245048 4.02309241e-07 -0.0410570554 4.02409241e-07 0.037700894
+ 4.02509241e-07 -0.0342011994 4.02609241e-07 0.0313787965 4.02709241e-07 -0.0285001312 4.02809241e-07 0.0261309755 4.02909241e-07 -0.0237572942 4.03009241e-07 0.0217710974 4.03109241e-07 -0.0198097687 4.03209241e-07 0.0181460851
+ 4.03309241e-07 -0.0165226519 4.03409241e-07 0.0151299819 4.03509241e-07 -0.0137842547 4.03609241e-07 0.0126189805 4.03709241e-07 -0.0115020691 4.03809241e-07 0.0105273918 4.03909241e-07 -0.00959941956 4.04009241e-07 0.00878437449
+ 4.04109241e-07 -0.0080127004 4.04209241e-07 0.00733127901 4.04309241e-07 -0.00668910201 4.04409241e-07 0.00611948647 4.04509241e-07 -0.00558474235 4.04609241e-07 0.00510864727 4.04709241e-07 -0.00466313017 4.04809241e-07 0.00426524119
+ 4.04909241e-07 -0.00389389982 4.05009241e-07 0.00356139756 4.05109241e-07 -0.00325176812 4.05209241e-07 0.00297392599 4.05309241e-07 -0.00271567297 4.05409241e-07 0.00248351831 4.05509241e-07 -0.00226806096 4.05609241e-07 0.00207409017
+ 4.05709241e-07 -0.00189429747 4.05809241e-07 0.00173223667 4.05909241e-07 -0.00158217745 4.06009241e-07 0.00144678179 4.06109241e-07 -0.00132151935 4.06209241e-07 0.00120840479 4.06309241e-07 -0.00110382775 4.06409241e-07 0.0010093302
+ 4.06509241e-07 -0.000922012818 4.06609241e-07 0.000843070142 4.06709241e-07 -0.00077015679 4.06809241e-07 0.000704210127 4.06909241e-07 -0.000641698121 4.07009241e-07 0.000588620508 4.07109241e-07 -0.000537460404 4.07209241e-07 0.00049143601
+ 4.07309241e-07 -0.000448954494 4.07409241e-07 0.000410509151 4.07509241e-07 -0.00037502548 4.07609241e-07 0.000342912489 4.07709241e-07 -0.000313272133 4.07809241e-07 0.000286449239 4.07909241e-07 -0.000260434291 4.08009241e-07 0.000239494613
+ 4.08109241e-07 -0.000217572043 4.08209241e-07 0.000200138431 4.08309241e-07 -0.000181776513 4.08409241e-07 0.000168412028 4.08509241e-07 -0.000151700166 4.08609241e-07 0.000140636669 4.08709241e-07 -0.000126668718 4.08809241e-07 0.000117445566
+ 4.08909241e-07 -0.00010577273 4.09009241e-07 9.80823968e-05 4.09109241e-07 -8.83271665e-05 4.09209241e-07 8.19142604e-05 4.09309241e-07 -7.37611653e-05 4.09409241e-07 6.84132514e-05 4.09509241e-07 -6.15986662e-05 4.09609241e-07 5.71389142e-05
+ 4.09709241e-07 -5.14425502e-05 4.09809241e-07 4.77236794e-05 4.09909241e-07 -4.29614712e-05 4.10009241e-07 3.98607554e-05 4.10109241e-07 -3.5878914e-05 4.10209241e-07 3.32940479e-05 4.10309241e-07 -2.99640861e-05 4.10409241e-07 2.78097581e-05
+ 4.10509241e-07 -2.50243268e-05 4.10609241e-07 2.32293653e-05 4.10709241e-07 -2.08987797e-05 4.10809241e-07 1.94038161e-05 4.10909241e-07 -1.7453167e-05 4.11009241e-07 1.62086675e-05 4.11109241e-07 -1.45753822e-05 4.11209241e-07 1.35400087e-05
+ 4.11309241e-07 -1.21718182e-05 4.11409241e-07 1.13110661e-05 4.11509241e-07 -1.01643087e-05 4.11609241e-07 9.44937439e-06 4.11709241e-07 -8.48757837e-06 4.11809241e-07 7.89441434e-06 4.11909241e-07 -7.08713851e-06 4.12009241e-07 6.59570205e-06
+ 4.12109241e-07 -5.91746374e-06 4.12209241e-07 5.51092447e-06 4.12309241e-07 -4.94046151e-06 4.12409241e-07 4.60484172e-06 4.12509241e-07 -4.12441064e-06 4.12609241e-07 3.84802635e-06 4.12709241e-07 -3.44279985e-06 4.12809241e-07 3.21589029e-06
+ 4.12909241e-07 -2.8734813e-06 4.13009241e-07 2.68789385e-06 4.13109241e-07 -2.39795499e-06 4.13209241e-07 2.2468806e-06 4.13309241e-07 -2.00076871e-06 4.13409241e-07 1.87852049e-06 4.13509241e-07 -1.66901602e-06 4.13609241e-07 1.57084431e-06
+ 4.13709241e-07 -1.39191691e-06 4.13809241e-07 1.31385476e-06 4.13909241e-07 -1.16046737e-06 4.14009241e-07 1.09920149e-06 4.14109241e-07 -9.67146834e-07 4.14209241e-07 9.19909936e-07 4.14309241e-07 -8.05673783e-07 4.14409241e-07 7.70154473e-07
+ 4.14509241e-07 -6.7080149e-07 4.14609241e-07 6.45069406e-07 4.14709241e-07 -5.58147936e-07 4.14809241e-07 5.40590661e-07 4.14909241e-07 -4.64052764e-07 4.15009241e-07 4.53323507e-07 4.15109241e-07 -3.8545863e-07 4.15209241e-07 3.80432504e-07
+ 4.15309241e-07 -3.19811888e-07 4.15409241e-07 3.1954934e-07 4.15509241e-07 -2.64979597e-07 4.15609241e-07 2.68695866e-07 4.15709241e-07 -2.19180201e-07 4.15809241e-07 2.26219815e-07 4.15909241e-07 -1.8092564e-07 4.16009241e-07 1.90741111e-07
+ 4.16109241e-07 -1.48972995e-07 4.16209241e-07 1.6110703e-07 4.16309241e-07 -1.22284104e-07 4.16409241e-07 1.36354747e-07 4.16509241e-07 -9.99918295e-08 4.16609241e-07 1.15680046e-07 4.16709241e-07 -8.13718871e-08 4.16809241e-07 9.84112047e-08
+ 4.16909241e-07 -6.58223732e-08 4.17009241e-07 8.39929854e-08 4.17109241e-07 -5.28400399e-08 4.17209241e-07 7.19556154e-08 4.17309241e-07 -4.2001428e-08 4.17409241e-07 6.19059216e-08 4.17509241e-07 -3.29525414e-08 4.17609241e-07 5.35156811e-08
+ 4.17709241e-07 -2.53978478e-08 4.17809241e-07 4.65108741e-08 4.17909241e-07 -1.90906165e-08 4.18009241e-07 4.06627305e-08 4.18109241e-07 -1.38111838e-08 4.18209241e-07 3.57678315e-08 4.18309241e-07 -9.41798334e-09 4.18409241e-07 3.1694159e-08
+ 4.18509241e-07 -5.74987452e-09 4.18609241e-07 2.82930291e-08 4.18709241e-07 -2.68736189e-09 4.18809241e-07 2.54534267e-08 4.18909241e-07 -1.30474076e-10 4.19009241e-07 2.30826487e-08 4.19109241e-07 2.0042642e-09 4.19209241e-07 2.11293847e-08
+ 4.19309241e-07 3.76433662e-09 4.19409241e-07 1.95203311e-08 4.19509241e-07 5.21432739e-09 4.19609241e-07 1.81947455e-08 4.19709241e-07 6.40887912e-09 4.19809241e-07 1.71026803e-08 4.19909241e-07 7.39299616e-09 4.20009241e-07 1.62029944e-08
+ 4.20109241e-07 8.20375165e-09 4.20209241e-07 1.53618153e-08 4.20309241e-07 8.8574762e-09 4.20409241e-07 1.47630591e-08 4.20509241e-07 9.40108799e-09 4.20609241e-07 1.42694719e-08 4.20709241e-07 9.84925339e-09 4.20809241e-07 1.38625606e-08
+ 4.20909241e-07 1.02187129e-08 4.21009241e-07 1.35271143e-08 4.21109241e-07 1.05232837e-08 4.21209241e-07 1.3250585e-08 4.21309241e-07 1.07743598e-08 4.21409241e-07 1.30226261e-08 4.21509241e-07 1.09813363e-08 4.21609241e-07 1.28347068e-08
+ 4.21709241e-07 1.11519594e-08 4.21809241e-07 1.26797947e-08 4.21909241e-07 1.12926134e-08 4.22009241e-07 1.25520922e-08 4.22109241e-07 1.14085626e-08 4.22209241e-07 1.24468206e-08 4.22309241e-07 1.1504146e-08 4.22409241e-07 1.2360039e-08
+ 4.22509241e-07 1.1582941e-08 4.22609241e-07 1.22885009e-08 4.22709241e-07 1.1647896e-08 4.22809241e-07 1.22295282e-08 4.22909241e-07 1.17014423e-08 4.23009241e-07 1.21809137e-08 4.23109241e-07 1.17455835e-08 4.23209241e-07 1.21408383e-08
+ 4.23309241e-07 1.1781972e-08 4.23409241e-07 1.21078022e-08 4.23509241e-07 1.18119692e-08 4.23609241e-07 1.20805691e-08 4.23709241e-07 1.18366976e-08 4.23809241e-07 1.20581191e-08 4.23909241e-07 1.18570829e-08 4.24009241e-07 1.2039613e-08
+ 4.24109241e-07 1.18738874e-08 4.24209241e-07 1.20243573e-08 4.24309241e-07 1.18877405e-08 4.24409241e-07 1.20117812e-08 4.24509241e-07 1.18991607e-08 4.24609241e-07 1.20014142e-08 4.24709241e-07 1.19085752e-08 4.24809241e-07 1.19928685e-08
+ 4.24909241e-07 1.1916336e-08 4.25009241e-07 1.19858237e-08 4.25109241e-07 1.19227338e-08 4.25209241e-07 1.19800167e-08 4.25309241e-07 1.1928008e-08 4.25409241e-07 1.19752293e-08 4.25509241e-07 1.1932356e-08 4.25609241e-07 1.19712831e-08
+ 4.25709241e-07 1.19359405e-08 4.25809241e-07 1.19680301e-08 4.25909241e-07 1.19388954e-08 4.26009241e-07 1.19653485e-08 4.26109241e-07 1.19413317e-08 4.26209241e-07 1.19631381e-08 4.26309241e-07 1.19433398e-08 4.26409241e-07 1.19613163e-08
+ 4.26509241e-07 1.19449952e-08 4.26609241e-07 1.19598143e-08 4.26709241e-07 1.19463603e-08 4.26809241e-07 1.19585764e-08 4.26909241e-07 1.19474858e-08 4.27009241e-07 1.19575561e-08 4.27109241e-07 1.19484131e-08 4.27209241e-07 1.19567147e-08
+ 4.27309241e-07 1.19491778e-08 4.27409241e-07 1.19560216e-08 4.27509241e-07 1.19498085e-08 4.27609241e-07 1.19554502e-08 4.27709241e-07 1.19503281e-08 4.27809241e-07 1.19549796e-08 4.27909241e-07 1.19507571e-08 4.28009241e-07 1.1954591e-08
+ 4.28109241e-07 1.19511105e-08 4.28209241e-07 1.19542709e-08 4.28309241e-07 1.19514019e-08 4.28409241e-07 1.19540074e-08 4.28509241e-07 1.19516422e-08 4.28609241e-07 1.19537901e-08 4.28709241e-07 1.19518406e-08 4.28809241e-07 1.19536112e-08
+ 4.28909241e-07 1.19520038e-08 4.29009241e-07 1.19534636e-08 4.29109241e-07 1.19521388e-08 4.29209241e-07 1.19533421e-08 4.29309241e-07 1.19522498e-08 4.29409241e-07 1.19532421e-08 4.29509241e-07 1.19523416e-08 4.29609241e-07 1.19531595e-08
+ 4.29709241e-07 1.19524172e-08 4.29809241e-07 1.19530916e-08 4.29909241e-07 1.19524796e-08 4.30009241e-07 1.19530356e-08 4.30109241e-07 1.19525312e-08 4.30209241e-07 1.19529896e-08 4.30309241e-07 1.19525737e-08 4.30409241e-07 1.19529517e-08
+ 4.30509241e-07 1.19526087e-08 4.30609241e-07 1.19529205e-08 4.30709241e-07 1.19526376e-08 4.30809241e-07 1.1952895e-08 4.30909241e-07 1.19526615e-08 4.31009241e-07 1.19528739e-08 4.31109241e-07 1.19526815e-08 4.31209241e-07 1.19528563e-08
+ 4.31309241e-07 1.19526979e-08 4.31409241e-07 1.19528421e-08 4.31509241e-07 1.19527114e-08 4.31609241e-07 1.19528302e-08 4.31709241e-07 1.19527227e-08 4.31809241e-07 1.19528207e-08 4.31909241e-07 1.19527321e-08 4.32009241e-07 1.19528129e-08
+ 4.32109241e-07 1.195274e-08 4.32209241e-07 1.19528062e-08 4.32309241e-07 1.19527462e-08 4.32409241e-07 1.19528013e-08 4.32509241e-07 1.19527515e-08 4.32609241e-07 1.1952797e-08 4.32709241e-07 1.19527562e-08 4.32809241e-07 1.19527933e-08
+ 4.32909241e-07 1.19527596e-08 4.33009241e-07 1.19527905e-08 4.33109241e-07 1.19527629e-08 4.33209241e-07 1.19527881e-08 4.33309241e-07 1.19527652e-08 4.33409241e-07 1.19527862e-08 4.33509241e-07 1.19527677e-08 4.33609241e-07 1.19527844e-08
+ 4.33709241e-07 1.19527695e-08 4.33809241e-07 1.19527831e-08 4.33909241e-07 1.19527709e-08 4.34009241e-07 1.19527825e-08 4.34109241e-07 1.19527723e-08 4.34209241e-07 1.19527816e-08 4.34309241e-07 1.1952773e-08 4.34409241e-07 1.19527811e-08
+ 4.34509241e-07 1.19527742e-08 4.34609241e-07 1.19527806e-08 4.34709241e-07 1.1952775e-08 4.34809241e-07 1.19527803e-08 4.34909241e-07 1.19527755e-08 4.35009241e-07 1.19527798e-08 4.35109241e-07 1.19527765e-08 4.35209241e-07 1.19527798e-08
+ 4.35309241e-07 1.19527769e-08 4.35409241e-07 1.19527795e-08 4.35509241e-07 1.19527774e-08 4.35609241e-07 1.195278e-08 4.35709241e-07 1.19527777e-08 4.35809241e-07 1.19527796e-08 4.35909241e-07 1.19527777e-08 4.36009241e-07 1.19527797e-08
+ 4.36109241e-07 1.19527781e-08 4.36209241e-07 1.195278e-08 4.36309241e-07 1.19527783e-08 4.36409241e-07 1.19527801e-08 4.36509241e-07 1.19527786e-08 4.36609241e-07 1.19527798e-08 4.36709241e-07 1.1952779e-08 4.36809241e-07 1.19527798e-08
+ 4.36909241e-07 1.19527794e-08 4.37009241e-07 1.195278e-08 4.37109241e-07 1.19527793e-08 4.37209241e-07 1.19527801e-08 4.37309241e-07 1.19527796e-08 4.37409241e-07 1.19527802e-08 4.37509241e-07 1.19527801e-08 4.37609241e-07 1.19527805e-08
+ 4.37709241e-07 1.19527803e-08 4.37809241e-07 1.19527805e-08 4.37909241e-07 1.19527802e-08 4.38009241e-07 1.19527807e-08 4.38109241e-07 1.19527803e-08 4.38209241e-07 1.19527808e-08 4.38309241e-07 1.19527805e-08 4.38409241e-07 1.19527805e-08
+ 4.38509241e-07 1.19527805e-08 4.38609241e-07 1.19527808e-08 4.38709241e-07 1.1952781e-08 4.38809241e-07 1.1952781e-08 4.38909241e-07 1.19527809e-08 4.39009241e-07 1.19527809e-08 4.39109241e-07 1.19527812e-08 4.39209241e-07 1.19527812e-08
+ 4.39309241e-07 1.19527815e-08 4.39409241e-07 1.19527815e-08 4.39509241e-07 1.19527812e-08 4.39609241e-07 1.19527817e-08 4.39709241e-07 1.19527816e-08 4.39809241e-07 1.19527814e-08 4.39909241e-07 1.19527816e-08 4.40009241e-07 1.19527817e-08
+ 4.40109241e-07 1.19527818e-08 4.40209241e-07 1.1952782e-08 4.40309241e-07 1.19527818e-08 4.40409241e-07 1.19527819e-08 4.40509241e-07 1.19527818e-08 4.40609241e-07 1.19527822e-08 4.40709241e-07 1.1952782e-08 4.40809241e-07 1.19527822e-08
+ 4.40909241e-07 1.19527818e-08 4.41009241e-07 1.19527822e-08 4.41109241e-07 1.19527819e-08 4.41209241e-07 1.19527825e-08 4.41309241e-07 1.19527821e-08 4.41409241e-07 1.19527822e-08 4.41509241e-07 1.19527822e-08 4.41609241e-07 1.19527826e-08
+ 4.41709241e-07 1.19527824e-08 4.41809241e-07 1.19527828e-08 4.41909241e-07 1.19527824e-08 4.42009241e-07 1.19527829e-08 4.42109241e-07 1.19527827e-08 4.42209241e-07 1.19527826e-08 4.42309241e-07 1.19527826e-08 4.42409241e-07 1.19527828e-08
+ 4.42509241e-07 1.19527827e-08 4.42609241e-07 1.19527831e-08 4.42709241e-07 1.19527827e-08 4.42809241e-07 1.19527828e-08 4.42909241e-07 1.19527827e-08 4.43009241e-07 1.19527834e-08 4.43109241e-07 1.19527828e-08 4.43209241e-07 1.19527832e-08
+ 4.43309241e-07 1.19527831e-08 4.43409241e-07 1.19527834e-08 4.43509241e-07 1.19527833e-08 4.43609241e-07 1.19527833e-08 4.43709241e-07 1.19527832e-08 4.43809241e-07 1.19527834e-08 4.43909241e-07 1.19527835e-08 4.44009241e-07 1.19527832e-08
+ 4.44109241e-07 1.19527834e-08 4.44209241e-07 1.19527835e-08 4.44309241e-07 1.19527837e-08 4.44409241e-07 1.19527833e-08 4.44509241e-07 1.19527838e-08 4.44609241e-07 1.19527834e-08 4.44709241e-07 1.19527835e-08 4.44809241e-07 1.19527838e-08
+ 4.44909241e-07 1.19527838e-08 4.45009241e-07 1.1952784e-08 4.45109241e-07 1.19527838e-08 4.45209241e-07 1.19527837e-08 4.45309241e-07 1.19527837e-08 4.45409241e-07 1.19527837e-08 4.45509241e-07 1.1952784e-08 4.45609241e-07 1.19527841e-08
+ 4.45709241e-07 1.1952784e-08 4.45809241e-07 1.1952784e-08 4.45909241e-07 1.19527841e-08 4.46009241e-07 1.19527841e-08 4.46109241e-07 1.19527842e-08 4.46209241e-07 1.19527842e-08 4.46309241e-07 1.1952784e-08 4.46409241e-07 1.19527842e-08
+ 4.46509241e-07 1.19527844e-08 4.46609241e-07 1.19527843e-08 4.46709241e-07 1.19527841e-08 4.46809241e-07 1.19527842e-08 4.46909241e-07 1.19527846e-08 4.47009241e-07 1.19527842e-08 4.47109241e-07 1.19527845e-08 4.47209241e-07 1.19527841e-08
+ 4.47309241e-07 1.19527847e-08 4.47409241e-07 1.19527844e-08 4.47509241e-07 1.19527847e-08 4.47609241e-07 1.19527845e-08 4.47709241e-07 1.19527847e-08 4.47809241e-07 1.19527843e-08 4.47909241e-07 1.19527847e-08 4.48009241e-07 1.19527843e-08
+ 4.48109241e-07 1.19527848e-08 4.48209241e-07 1.19527844e-08 4.48309241e-07 1.19527851e-08 4.48409241e-07 1.19527847e-08 4.48509241e-07 1.1952785e-08 4.48609241e-07 1.19527843e-08 4.48709241e-07 1.19527852e-08 4.48809241e-07 1.19527844e-08
+ 4.48909241e-07 1.19527852e-08 4.49009241e-07 1.19527845e-08 4.49109241e-07 1.19527853e-08 4.49209241e-07 1.19527845e-08 4.49309241e-07 1.19527853e-08 4.49409241e-07 1.19527847e-08 4.49509241e-07 1.1952785e-08 4.49609241e-07 1.19527849e-08
+ 4.49709241e-07 1.19527851e-08 4.49809241e-07 1.19527848e-08 4.49909241e-07 1.19527852e-08 4.50009241e-07 1.19527849e-08 4.50109241e-07 1.19527849e-08 4.50209241e-07 1.1952785e-08 4.50309241e-07 1.19527853e-08 4.50409241e-07 1.19527853e-08
+ 4.50509241e-07 1.1952785e-08 4.50609241e-07 1.19527854e-08 4.50709241e-07 1.19527851e-08 4.50809241e-07 1.19527855e-08 4.50909241e-07 1.19527853e-08 4.51e-07 1.19527852e-08 4.5101e-07 1.19390964e-08 4.5103e-07 1.20196141e-08
+ 4.5107e-07 1.18477351e-08 4.5115e-07 1.20721808e-08 4.5125e-07 1.18298605e-08 4.5135e-07 1.2069468e-08 4.5145e-07 1.1851929e-08 4.5155e-07 1.20304653e-08 4.5165e-07 1.19012718e-08 4.5175e-07 1.19750949e-08
+ 4.5185e-07 1.19638076e-08 4.51930828e-07 1.89264353e-07 4.52e-07 2.6011952e-07 4.52008608e-07 -7.14340553e-06 4.52025825e-07 -6.92152579e-06 4.52060258e-07 1.22318635e-05 4.52106181e-07 -2.07308553e-07 4.52150081e-07 -6.86147133e-06
+ 4.52198026e-07 -7.40021862e-07 4.5225538e-07 5.62676254e-06 4.52312019e-07 -4.8081976e-06 4.52404232e-07 3.76387955e-06 4.52504232e-07 -3.03362411e-06 4.52604232e-07 2.49152677e-06 4.52704232e-07 -2.0066143e-06 4.52804232e-07 1.66419859e-06
+ 4.52904232e-07 -1.34587456e-06 4.53004232e-07 1.13667787e-06 4.53104232e-07 -9.25169787e-07 4.53204232e-07 7.99904053e-07 4.53304232e-07 -6.55185529e-07 4.53404232e-07 5.82278078e-07 4.53504232e-07 -4.79264614e-07 4.53604232e-07 4.39148788e-07
+ 4.53704232e-07 -3.62367893e-07 4.53804232e-07 3.42983277e-07 4.53904232e-07 -2.82863542e-07 4.54004232e-07 2.7670735e-07 4.54104232e-07 -2.27290235e-07 4.54204232e-07 2.29706838e-07 4.54304232e-07 -1.87298528e-07 4.54404232e-07 1.95374429e-07
+ 4.54504232e-07 -1.5762143e-07 4.54604232e-07 1.69487684e-07 4.54704232e-07 -1.34878215e-07 4.54804232e-07 1.49328817e-07 4.54904232e-07 -1.16888777e-07 4.55004232e-07 1.33147156e-07 4.55104232e-07 -1.02245866e-07 4.55204232e-07 1.19804709e-07
+ 4.55304232e-07 -9.0026523e-08 4.55404232e-07 1.08549071e-07 4.55504232e-07 -7.96164004e-08 4.55604232e-07 9.88760457e-08 4.55704232e-07 -7.05996948e-08 4.55804232e-07 9.04391846e-08 4.55904232e-07 -6.2686541e-08 4.56004232e-07 8.29959183e-08
+ 4.56104232e-07 -5.56733952e-08 4.56204232e-07 7.63728478e-08 4.56304232e-07 -4.94109317e-08 4.56404232e-07 7.04403304e-08 4.56504232e-07 -4.37857097e-08 4.56604232e-07 6.50985338e-08 4.56704232e-07 -3.87103507e-08 4.56804232e-07 6.0270823e-08
+ 4.56904232e-07 -3.41165906e-08 4.57004232e-07 5.58953144e-08 4.57104232e-07 -2.9947954e-08 4.57204232e-07 5.19203753e-08 4.57304232e-07 -2.61574244e-08 4.57404232e-07 4.83032381e-08 4.57504232e-07 -2.27059202e-08 4.57604232e-07 4.50079067e-08
+ 4.57704232e-07 -1.95601254e-08 4.57804232e-07 4.20039858e-08 4.57904232e-07 -1.66928494e-08 4.58004232e-07 3.92662433e-08 4.58104232e-07 -1.40797467e-08 4.58204232e-07 3.67710487e-08 4.58304232e-07 -1.1697754e-08 4.58404232e-07 3.44962388e-08
+ 4.58504232e-07 -9.52592197e-09 4.58604232e-07 3.24219686e-08 4.58704232e-07 -7.54543122e-09 4.58804232e-07 3.05303505e-08 4.58904232e-07 -5.739243e-09 4.59004232e-07 2.88051115e-08 4.59104232e-07 -4.091814e-09 4.59204232e-07 2.72314284e-08
+ 4.59304232e-07 -2.58905e-09 4.59404232e-07 2.57959148e-08 4.59504232e-07 -1.21823585e-09 4.59604232e-07 2.44864712e-08 4.59704232e-07 3.19395066e-11 4.59804232e-07 2.32925136e-08 4.59904232e-07 1.16462459e-09 4.60004232e-07 2.22173191e-08
+ 4.60104232e-07 2.18546942e-09 4.60204232e-07 2.12478757e-08 4.60304232e-07 3.10627826e-09 4.60404232e-07 2.03731002e-08 4.60504232e-07 3.9374668e-09 4.60604232e-07 1.9583196e-08 4.60704232e-07 4.68825634e-09 4.60804232e-07 1.88694753e-08
+ 4.60904232e-07 5.366838e-09 4.61004232e-07 1.82242125e-08 4.61104232e-07 5.98050093e-09 4.61204232e-07 1.76405257e-08 4.61304232e-07 6.53574531e-09 4.61404232e-07 1.71122738e-08 4.61504232e-07 7.0383761e-09 4.61604232e-07 1.66339683e-08
+ 4.61704232e-07 7.49358262e-09 4.61804232e-07 1.62007002e-08 4.61904232e-07 7.90601137e-09 4.62004232e-07 1.58080699e-08 4.62104232e-07 8.27982835e-09 4.62204232e-07 1.54521331e-08 4.62304232e-07 8.61876867e-09 4.62404232e-07 1.51293527e-08
+ 4.62504232e-07 8.92618207e-09 4.62604232e-07 1.48365573e-08 4.62704232e-07 9.20506357e-09 4.62804232e-07 1.4570932e-08 4.62904232e-07 9.45804934e-09 4.63004232e-07 1.43299976e-08 4.63104232e-07 9.68749864e-09 4.63204232e-07 1.41114866e-08
+ 4.63304232e-07 9.89559759e-09 4.63404232e-07 1.39132949e-08 4.63504232e-07 1.00843645e-08 4.63604232e-07 1.37334932e-08 4.63704232e-07 1.02556396e-08 4.63804232e-07 1.35703296e-08 4.63904232e-07 1.04110868e-08 4.64004232e-07 1.34221844e-08
+ 4.64104232e-07 1.05522192e-08 4.64204232e-07 1.32880898e-08 4.64304232e-07 1.06794395e-08 4.64404232e-07 1.3166998e-08 4.64504232e-07 1.0795133e-08 4.64604232e-07 1.30563922e-08 4.64704232e-07 1.09007875e-08 4.64804232e-07 1.29555432e-08
+ 4.64904232e-07 1.09969992e-08 4.65004232e-07 1.28637764e-08 4.65104232e-07 1.10845362e-08 4.65204232e-07 1.27802766e-08 4.65304232e-07 1.11641361e-08 4.65404232e-07 1.27044499e-08 4.65504232e-07 1.12363761e-08 4.65604232e-07 1.26355459e-08
+ 4.65704232e-07 1.13021394e-08 4.65804232e-07 1.25728633e-08 4.65904232e-07 1.13617871e-08 4.66004232e-07 1.25161193e-08 4.66104232e-07 1.14157949e-08 4.66204232e-07 1.24646916e-08 4.66304232e-07 1.14647826e-08 4.66404232e-07 1.24180176e-08
+ 4.66504232e-07 1.15092594e-08 4.66604232e-07 1.237563e-08 4.66704232e-07 1.15496589e-08 4.66804232e-07 1.23371224e-08 4.66904232e-07 1.15863662e-08 4.67004232e-07 1.23021307e-08 4.67104232e-07 1.1619721e-08 4.67204232e-07 1.22703341e-08
+ 4.67304232e-07 1.16500729e-08 4.67404232e-07 1.22412999e-08 4.67504232e-07 1.16778119e-08 4.67604232e-07 1.22148984e-08 4.67704232e-07 1.17029105e-08 4.67804232e-07 1.21910167e-08 4.67904232e-07 1.17256513e-08 4.68004232e-07 1.21693516e-08
+ 4.68104232e-07 1.17462983e-08 4.68204232e-07 1.21496707e-08 4.68304232e-07 1.17650612e-08 4.68404232e-07 1.21317817e-08 4.68504232e-07 1.17821174e-08 4.68604232e-07 1.21155185e-08 4.68704232e-07 1.17976252e-08 4.68804232e-07 1.21007312e-08
+ 4.68904232e-07 1.18117253e-08 4.69004232e-07 1.20872868e-08 4.69104232e-07 1.18245444e-08 4.69204232e-07 1.20750639e-08 4.69304232e-07 1.18361993e-08 4.69404232e-07 1.20639507e-08 4.69504232e-07 1.1846796e-08 4.69604232e-07 1.20538464e-08
+ 4.69704232e-07 1.18564305e-08 4.69804232e-07 1.20446598e-08 4.69904232e-07 1.18651899e-08 4.70004232e-07 1.20363082e-08 4.70104232e-07 1.18731531e-08 4.70204232e-07 1.20287149e-08 4.70304232e-07 1.18803934e-08 4.70404232e-07 1.20218113e-08
+ 4.70504232e-07 1.1886976e-08 4.70604232e-07 1.20155352e-08 4.70704232e-07 1.18929603e-08 4.70804232e-07 1.20098294e-08 4.70904232e-07 1.18984008e-08 4.71004232e-07 1.20046417e-08 4.71104232e-07 1.19033474e-08 4.71204232e-07 1.19999252e-08
+ 4.71304232e-07 1.19078446e-08 4.71404232e-07 1.19956366e-08 4.71504232e-07 1.19119332e-08 4.71604232e-07 1.19917385e-08 4.71704232e-07 1.191565e-08 4.71804232e-07 1.1988195e-08 4.71904232e-07 1.19190288e-08 4.72004232e-07 1.19849733e-08
+ 4.72104232e-07 1.19221004e-08 4.72204232e-07 1.19820448e-08 4.72304232e-07 1.19248928e-08 4.72404232e-07 1.19793827e-08 4.72504232e-07 1.1927431e-08 4.72604232e-07 1.19769624e-08 4.72704232e-07 1.19297386e-08 4.72804232e-07 1.19747622e-08
+ 4.72904232e-07 1.19318362e-08 4.73004232e-07 1.19727623e-08 4.73104232e-07 1.19337437e-08 4.73204232e-07 1.1970944e-08 4.73304232e-07 1.1935477e-08 4.73404232e-07 1.1969291e-08 4.73504232e-07 1.19370532e-08 4.73604232e-07 1.19677883e-08
+ 4.73704232e-07 1.19384858e-08 4.73804232e-07 1.19664222e-08 4.73904232e-07 1.19397882e-08 4.74004232e-07 1.19651805e-08 4.74104232e-07 1.19409721e-08 4.74204232e-07 1.19640516e-08 4.74304232e-07 1.19420486e-08 4.74404232e-07 1.19630252e-08
+ 4.74504232e-07 1.19430271e-08 4.74604232e-07 1.19620926e-08 4.74704232e-07 1.19439165e-08 4.74804232e-07 1.19612444e-08 4.74904232e-07 1.19447251e-08 4.75004232e-07 1.19604736e-08 4.75104232e-07 1.194546e-08 4.75204232e-07 1.19597726e-08
+ 4.75304232e-07 1.19461283e-08 4.75404232e-07 1.19591356e-08 4.75504232e-07 1.19467359e-08 4.75604232e-07 1.19585564e-08 4.75704232e-07 1.19472881e-08 4.75804232e-07 1.19580298e-08 4.75904232e-07 1.19477901e-08 4.76004232e-07 1.19575511e-08
+ 4.76104232e-07 1.19482464e-08 4.76204232e-07 1.19571159e-08 4.76304232e-07 1.19486616e-08 4.76404232e-07 1.19567204e-08 4.76504232e-07 1.19490386e-08 4.76604232e-07 1.19563607e-08 4.76704232e-07 1.19493814e-08 4.76804232e-07 1.1956034e-08
+ 4.76904232e-07 1.19496932e-08 4.77004232e-07 1.19557368e-08 4.77104232e-07 1.19499765e-08 4.77204232e-07 1.19554666e-08 4.77304232e-07 1.19502341e-08 4.77404232e-07 1.19552209e-08 4.77504232e-07 1.1950468e-08 4.77604232e-07 1.19549981e-08
+ 4.77704232e-07 1.19506811e-08 4.77804232e-07 1.19547948e-08 4.77904232e-07 1.19508742e-08 4.78004232e-07 1.19546106e-08 4.78104232e-07 1.19510502e-08 4.78204232e-07 1.19544431e-08 4.78304232e-07 1.19512097e-08 4.78404232e-07 1.19542909e-08
+ 4.78504232e-07 1.1951355e-08 4.78604232e-07 1.19541526e-08 4.78704232e-07 1.19514868e-08 4.78804232e-07 1.19540269e-08 4.78904232e-07 1.19516066e-08 4.79004232e-07 1.1953913e-08 4.79104232e-07 1.19517152e-08 4.79204232e-07 1.19538094e-08
+ 4.79304232e-07 1.1951814e-08 4.79404232e-07 1.19537151e-08 4.79504232e-07 1.19519038e-08 4.79604232e-07 1.195363e-08 4.79704232e-07 1.19519848e-08 4.79804232e-07 1.19535523e-08 4.79904232e-07 1.19520586e-08 4.80004232e-07 1.19534823e-08
+ 4.80104232e-07 1.19521255e-08 4.80204232e-07 1.19534183e-08 4.80304232e-07 1.19521866e-08 4.80404232e-07 1.19533604e-08 4.80504232e-07 1.19522416e-08 4.80604232e-07 1.19533078e-08 4.80704232e-07 1.19522918e-08 4.80804232e-07 1.19532599e-08
+ 4.80904232e-07 1.19523373e-08 4.81004232e-07 1.19532166e-08 4.81104232e-07 1.19523784e-08 4.81204232e-07 1.19531776e-08 4.81304232e-07 1.1952416e-08 4.81404232e-07 1.19531418e-08 4.81504232e-07 1.19524499e-08 4.81604232e-07 1.19531095e-08
+ 4.81704232e-07 1.19524808e-08 4.81804232e-07 1.195308e-08 4.81904232e-07 1.19525088e-08 4.82004232e-07 1.19530532e-08 4.82104232e-07 1.19525343e-08 4.82204232e-07 1.19530289e-08 4.82304232e-07 1.19525575e-08 4.82404232e-07 1.19530069e-08
+ 4.82504232e-07 1.19525784e-08 4.82604232e-07 1.1952987e-08 4.82704232e-07 1.19525975e-08 4.82804232e-07 1.19529686e-08 4.82904232e-07 1.1952615e-08 4.83004232e-07 1.19529521e-08 4.83104232e-07 1.19526309e-08 4.83204232e-07 1.19529372e-08
+ 4.83304232e-07 1.19526453e-08 4.83404232e-07 1.19529233e-08 4.83504232e-07 1.19526581e-08 4.83604232e-07 1.19529112e-08 4.83704232e-07 1.195267e-08 4.83804232e-07 1.19529e-08 4.83904232e-07 1.19526806e-08 4.84004232e-07 1.19528896e-08
+ 4.84104232e-07 1.19526905e-08 4.84204232e-07 1.19528807e-08 4.84304232e-07 1.19526992e-08 4.84404232e-07 1.19528719e-08 4.84504232e-07 1.19527074e-08 4.84604232e-07 1.19528643e-08 4.84704232e-07 1.19527149e-08 4.84804232e-07 1.19528573e-08
+ 4.84904232e-07 1.19527213e-08 4.85004232e-07 1.19528511e-08 4.85104232e-07 1.19527272e-08 4.85204232e-07 1.19528455e-08 4.85304232e-07 1.19527329e-08 4.85404232e-07 1.19528401e-08 4.85504232e-07 1.19527377e-08 4.85604232e-07 1.19528353e-08
+ 4.85704232e-07 1.19527426e-08 4.85804232e-07 1.19528309e-08 4.85904232e-07 1.19527464e-08 4.86004232e-07 1.1952827e-08 4.86104232e-07 1.19527504e-08 4.86204232e-07 1.19528234e-08 4.86304232e-07 1.19527537e-08 4.86404232e-07 1.19528201e-08
+ 4.86504232e-07 1.19527571e-08 4.86604232e-07 1.19528171e-08 4.86704232e-07 1.19527596e-08 4.86804232e-07 1.19528143e-08 4.86904232e-07 1.19527623e-08 4.87004232e-07 1.1952812e-08 4.87104232e-07 1.19527647e-08 4.87204232e-07 1.19528097e-08
+ 4.87304232e-07 1.1952767e-08 4.87404232e-07 1.19528077e-08 4.87504232e-07 1.19527686e-08 4.87604232e-07 1.19528058e-08 4.87704232e-07 1.19527704e-08 4.87804232e-07 1.19528041e-08 4.87904232e-07 1.19527722e-08 4.88004232e-07 1.19528026e-08
+ 4.88104232e-07 1.19527737e-08 4.88204232e-07 1.19528012e-08 4.88304232e-07 1.19527749e-08 4.88404232e-07 1.19528e-08 4.88504232e-07 1.19527761e-08 4.88604232e-07 1.19527989e-08 4.88704232e-07 1.19527772e-08 4.88804232e-07 1.19527978e-08
+ 4.88904232e-07 1.1952778e-08 4.89004232e-07 1.19527973e-08 4.89104232e-07 1.19527788e-08 4.89204232e-07 1.19527963e-08 4.89304232e-07 1.19527795e-08 4.89404232e-07 1.19527953e-08 4.89504232e-07 1.19527807e-08 4.89604232e-07 1.19527945e-08
+ 4.89704232e-07 1.19527813e-08 4.89804232e-07 1.19527938e-08 4.89904232e-07 1.19527818e-08 4.90004232e-07 1.19527935e-08 4.90104232e-07 1.19527823e-08 4.90204232e-07 1.19527933e-08 4.90304232e-07 1.19527828e-08 4.90404232e-07 1.19527925e-08
+ 4.90504232e-07 1.19527832e-08 4.90604232e-07 1.1952792e-08 4.90704232e-07 1.19527837e-08 4.90804232e-07 1.19527918e-08 4.90904232e-07 1.19527841e-08 4.91004232e-07 1.19527912e-08 4.91104232e-07 1.19527845e-08 4.91204232e-07 1.19527911e-08
+ 4.91304232e-07 1.19527848e-08 4.91404232e-07 1.19527905e-08 4.91504232e-07 1.19527849e-08 4.91604232e-07 1.19527903e-08 4.91704232e-07 1.19527855e-08 4.91804232e-07 1.19527899e-08 4.91904232e-07 1.19527856e-08 4.92004232e-07 1.19527898e-08
+ 4.92104232e-07 1.19527858e-08 4.92204232e-07 1.195279e-08 4.92304232e-07 1.19527859e-08 4.92404232e-07 1.19527898e-08 4.92504232e-07 1.19527861e-08 4.92604232e-07 1.19527893e-08 4.92704232e-07 1.19527862e-08 4.92804232e-07 1.19527895e-08
+ 4.92904232e-07 1.19527864e-08 4.93004232e-07 1.19527893e-08 4.93104232e-07 1.19527865e-08 4.93204232e-07 1.19527891e-08 4.93304232e-07 1.19527868e-08 4.93404232e-07 1.1952789e-08 4.93504232e-07 1.19527868e-08 4.93604232e-07 1.19527888e-08
+ 4.93704232e-07 1.19527868e-08 4.93804232e-07 1.19527888e-08 4.93904232e-07 1.19527869e-08 4.94004232e-07 1.19527887e-08 4.94104232e-07 1.1952787e-08 4.94204232e-07 1.19527889e-08 4.94304232e-07 1.19527868e-08 4.94404232e-07 1.19527888e-08
+ 4.94504232e-07 1.19527872e-08 4.94604232e-07 1.19527885e-08 4.94704232e-07 1.19527871e-08 4.94804232e-07 1.19527882e-08 4.94904232e-07 1.19527875e-08 4.95004232e-07 1.19527881e-08 4.95104232e-07 1.19527873e-08 4.95204232e-07 1.19527883e-08
+ 4.95304232e-07 1.19527876e-08 4.95404232e-07 1.19527881e-08 4.95504232e-07 1.19527877e-08 4.95604232e-07 1.1952788e-08 4.95704232e-07 1.19527876e-08 4.95804232e-07 1.19527881e-08 4.95904232e-07 1.19527876e-08 4.96004232e-07 1.1952788e-08
+ 4.96104232e-07 1.1952788e-08 4.96204232e-07 1.19527879e-08 4.96304232e-07 1.19527877e-08 4.96404232e-07 1.1952788e-08 4.96504232e-07 1.19527878e-08 4.96604232e-07 1.19527879e-08 4.96704232e-07 1.19527877e-08 4.96804232e-07 1.1952788e-08
+ 4.96904232e-07 1.19527879e-08 4.97004232e-07 1.19527881e-08 4.97104232e-07 1.19527881e-08 4.97204232e-07 1.19527877e-08 4.97304232e-07 1.1952788e-08 4.97404232e-07 1.19527881e-08 4.97504232e-07 1.19527878e-08 4.97604232e-07 1.1952788e-08
+ 4.97704232e-07 1.1952788e-08 4.97804232e-07 1.19527878e-08 4.97904232e-07 1.1952788e-08 4.98004232e-07 1.19527879e-08 4.98104232e-07 1.19527878e-08 4.98204232e-07 1.19527877e-08 4.98304232e-07 1.1952788e-08 4.98404232e-07 1.1952788e-08
+ 4.98504232e-07 1.19527878e-08 4.98604232e-07 1.19527882e-08 4.98704232e-07 1.19527879e-08 4.98804232e-07 1.1952788e-08 4.98904232e-07 1.19527879e-08 4.99004232e-07 1.19527882e-08 4.99104232e-07 1.19527878e-08 4.99204232e-07 1.19527882e-08
+ 4.99304232e-07 1.19527878e-08 4.99404232e-07 1.19527879e-08 4.99504232e-07 1.19527878e-08 4.99604232e-07 1.19527881e-08 4.99704232e-07 1.19527879e-08 4.99804232e-07 1.19527878e-08 4.99904232e-07 1.19527879e-08 5e-07 1.19527881e-08
+ 5.0001e-07 1.19847862e-08 5.0003e-07 1.17957473e-08 5.0007e-07 1.21960663e-08 5.0015e-07 1.16790212e-08 5.0025e-07 1.22357527e-08 5.0035e-07 1.16768705e-08 5.0045e-07 1.22053472e-08 5.0055e-07 1.17434326e-08
+ 5.0065e-07 1.18632203e-08 5.0075e-07 2.60700187e-08 5.0085e-07 -6.67652971e-07 5.00932051e-07 4.41565399e-06 5.01e-07 -1.00425785e-05 5.01008488e-07 -1.02352439e-05 5.01025463e-07 4.62438714e-06 5.01059414e-07 6.10068297e-06
+ 5.0109062e-07 2.93430931e-06 5.0114347e-07 -1.23168868e-07 5.01199151e-07 8.33058792e-06 5.01299151e-07 -3.00514879e-05 5.01399151e-07 0.000133952605 5.01499151e-07 -0.000207264225 5.01599151e-07 0.000192426471 5.01699151e-07 -0.000285523601
+ 5.01799151e-07 0.000366852825 5.01893327e-07 -0.00036846974 5.01993327e-07 0.000376973588 5.02093327e-07 -0.000371315116 5.02193327e-07 0.000359140809 5.02293327e-07 -0.000341874797 5.02393327e-07 0.000321770317 5.02493327e-07 -0.000299895372
+ 5.02593327e-07 0.000277811836 5.02693327e-07 -0.000255845433 5.02793327e-07 0.000234952298 5.02893327e-07 -0.000215003446 5.02993327e-07 0.000196566982 5.03093327e-07 -0.000179310692 5.03193327e-07 0.000163591693 5.03293327e-07 -0.000149019485
+ 5.03393327e-07 0.0001358423 5.03493327e-07 -0.00012367801 5.03593327e-07 0.000112719887 5.03693327e-07 -0.000102618211 5.03793327e-07 9.35370426e-05 5.03893327e-07 -8.51645593e-05 5.03993327e-07 7.76479395e-05 5.04093327e-07 -7.07110531e-05
+ 5.04193327e-07 6.44902504e-05 5.04293327e-07 -5.87404539e-05 5.04393327e-07 5.35903595e-05 5.04493327e-07 -4.88209881e-05 5.04593327e-07 4.45552201e-05 5.04693327e-07 -4.05956834e-05 5.04793327e-07 3.70606357e-05 5.04893327e-07 -3.37704863e-05
+ 5.04993327e-07 3.08397242e-05 5.05093327e-07 -2.81033671e-05 5.05193327e-07 2.56727906e-05 5.05293327e-07 -2.33950168e-05 5.05393327e-07 2.13788324e-05 5.05493327e-07 -1.94811354e-05 5.05593327e-07 1.78085526e-05 5.05693327e-07 -1.62261184e-05
+ 5.05793327e-07 1.48386552e-05 5.05893327e-07 -1.35179108e-05 5.05993327e-07 1.23671987e-05 5.06093327e-07 -1.12638134e-05 5.06193327e-07 1.03098066e-05 5.06293327e-07 -9.38706102e-06 5.06393327e-07 8.59657348e-06 5.06493327e-07 -7.824026e-06
+ 5.06593327e-07 7.16953335e-06 5.06693327e-07 -6.48075399e-06 5.06793327e-07 5.98664906e-06 5.06893327e-07 -5.40521902e-06 5.06993327e-07 4.9972539e-06 5.07093327e-07 -4.50840114e-06 5.07193327e-07 4.17217679e-06 5.07293327e-07 -3.76047466e-06
+ 5.07393327e-07 3.48401778e-06 5.07493327e-07 -3.13661854e-06 5.07593327e-07 2.90996505e-06 5.07693327e-07 -2.61617076e-06 5.07793327e-07 2.43102733e-06 5.07893327e-07 -2.18192815e-06 5.07993327e-07 2.04442042e-06 5.08093327e-07 -1.81749786e-06
+ 5.08193327e-07 1.70770947e-06 5.08293327e-07 -1.51444849e-06 5.08393327e-07 1.42684781e-06 5.08493327e-07 -1.26166668e-06 5.08593327e-07 1.1925578e-06 5.08693327e-07 -1.05078906e-06 5.08793327e-07 9.97096861e-07 5.08893327e-07 -8.74852071e-07
+ 5.08993327e-07 8.34014161e-07 5.09093327e-07 -7.28053117e-07 5.09193327e-07 6.97935565e-07 5.09293327e-07 -6.05557653e-07 5.09393327e-07 5.84381408e-07 5.09493327e-07 -5.03334641e-07 5.09593327e-07 4.89616695e-07 5.09693327e-07 -4.18023602e-07
+ 5.09793327e-07 4.10527791e-07 5.09893327e-07 -3.46822422e-07 5.09993327e-07 3.44517445e-07 5.10093327e-07 -2.87393597e-07 5.10193327e-07 2.89419646e-07 5.10293327e-07 -2.37788026e-07 5.10393327e-07 2.4342808e-07 5.10493327e-07 -1.96380018e-07
+ 5.10593327e-07 2.05035977e-07 5.10693327e-07 -1.61813343e-07 5.10793327e-07 1.72986222e-07 5.10893327e-07 -1.32956444e-07 5.10993327e-07 1.4622993e-07 5.11093327e-07 -1.08865152e-07 5.11193327e-07 1.23891857e-07 5.11293327e-07 -8.87516066e-08
+ 5.11393327e-07 1.05241666e-07 5.11493327e-07 -7.19604537e-08 5.11593327e-07 8.96740329e-08 5.11693327e-07 -5.7945955e-08 5.11793327e-07 7.66819097e-08 5.11893327e-07 -4.62495986e-08 5.11993327e-07 6.58388037e-08 5.12093327e-07 -3.64880341e-08
+ 5.12193327e-07 5.67891468e-08 5.12293327e-07 -2.83407877e-08 5.12393327e-07 4.9235939e-08 5.12493327e-07 -2.15406662e-08 5.12593327e-07 4.29315531e-08 5.12693327e-07 -1.58507319e-08 5.12793327e-07 3.76566188e-08 5.12893327e-07 -1.11162827e-08
+ 5.12993327e-07 3.32669801e-08 5.13093327e-07 -7.16407417e-09 5.13193327e-07 2.96027727e-08 5.13293327e-07 -3.86498902e-09 5.13393327e-07 2.65440783e-08 5.13493327e-07 -1.11106202e-09 5.13593327e-07 2.39907996e-08 5.13693327e-07 1.18782961e-09
+ 5.13793327e-07 2.18748402e-08 5.13893327e-07 3.09374742e-09 5.13993327e-07 2.01325724e-08 5.14093327e-07 4.66365543e-09 5.14193327e-07 1.86974615e-08 5.14293327e-07 5.95680469e-09 5.14393327e-07 1.75153374e-08 5.14493327e-07 7.02199834e-09
+ 5.14593327e-07 1.65415938e-08 5.14693327e-07 7.89942534e-09 5.14793327e-07 1.57394952e-08 5.14893327e-07 8.62218719e-09 5.14993327e-07 1.49812767e-08 5.15093327e-07 9.20369131e-09 5.15193327e-07 1.44482747e-08 5.15293327e-07 9.68756086e-09
+ 5.15393327e-07 1.40089632e-08 5.15493327e-07 1.00864088e-08 5.15593327e-07 1.36468572e-08 5.15693327e-07 1.04151538e-08 5.15793327e-07 1.33484019e-08 5.15893327e-07 1.06861085e-08 5.15993327e-07 1.31024163e-08 5.16093327e-07 1.09094248e-08
+ 5.16193327e-07 1.2899682e-08 5.16293327e-07 1.10934721e-08 5.16393327e-07 1.27326001e-08 5.16493327e-07 1.12451506e-08 5.16593327e-07 1.25949073e-08 5.16693327e-07 1.13701464e-08 5.16793327e-07 1.24814388e-08 5.16893327e-07 1.1473149e-08
+ 5.16993327e-07 1.23879382e-08 5.17093327e-07 1.15580225e-08 5.17193327e-07 1.23108973e-08 5.17293327e-07 1.16279524e-08 5.17393327e-07 1.22474232e-08 5.17493327e-07 1.1685565e-08 5.17593327e-07 1.21951318e-08 5.17693327e-07 1.17330256e-08
+ 5.17793327e-07 1.21520569e-08 5.17893327e-07 1.17721191e-08 5.17993327e-07 1.2116578e-08 5.18093327e-07 1.18043163e-08 5.18193327e-07 1.20873599e-08 5.18293327e-07 1.18308301e-08 5.18393327e-07 1.20633014e-08 5.18493327e-07 1.18526595e-08
+ 5.18593327e-07 1.20434955e-08 5.18693327e-07 1.18706287e-08 5.18793327e-07 1.20271936e-08 5.18893327e-07 1.18854168e-08 5.18993327e-07 1.20137794e-08 5.19093327e-07 1.18975839e-08 5.19193327e-07 1.20027446e-08 5.19293327e-07 1.19075908e-08
+ 5.19393327e-07 1.1993671e-08 5.19493327e-07 1.19158181e-08 5.19593327e-07 1.1986211e-08 5.19693327e-07 1.19225814e-08 5.19793327e-07 1.19800806e-08 5.19893327e-07 1.19281375e-08 5.19993327e-07 1.19750459e-08 5.20093327e-07 1.19326989e-08
+ 5.20193327e-07 1.19709139e-08 5.20293327e-07 1.19364417e-08 5.20393327e-07 1.19675244e-08 5.20493327e-07 1.19395104e-08 5.20593327e-07 1.19647463e-08 5.20693327e-07 1.1942025e-08 5.20793327e-07 1.19624706e-08 5.20893327e-07 1.19440839e-08
+ 5.20993327e-07 1.19606085e-08 5.21093327e-07 1.19457677e-08 5.21193327e-07 1.19590861e-08 5.21293327e-07 1.19471437e-08 5.21393327e-07 1.19578434e-08 5.21493327e-07 1.19482659e-08 5.21593327e-07 1.19568302e-08 5.21693327e-07 1.19491801e-08
+ 5.21793327e-07 1.19560054e-08 5.21893327e-07 1.19499238e-08 5.21993327e-07 1.19553349e-08 5.22093327e-07 1.19505278e-08 5.22193327e-07 1.19547912e-08 5.22293327e-07 1.19510175e-08 5.22393327e-07 1.19543507e-08 5.22493327e-07 1.19514133e-08
+ 5.22593327e-07 1.19539955e-08 5.22693327e-07 1.19517322e-08 5.22793327e-07 1.19537093e-08 5.22893327e-07 1.19519887e-08 5.22993327e-07 1.19534793e-08 5.23093327e-07 1.19521941e-08 5.23193327e-07 1.19532957e-08 5.23293327e-07 1.19523583e-08
+ 5.23393327e-07 1.19531496e-08 5.23493327e-07 1.19524882e-08 5.23593327e-07 1.1953034e-08 5.23693327e-07 1.19525908e-08 5.23793327e-07 1.19529433e-08 5.23893327e-07 1.19526709e-08 5.23993327e-07 1.19528726e-08 5.24093327e-07 1.19527333e-08
+ 5.24193327e-07 1.19528182e-08 5.24293327e-07 1.19527805e-08 5.24393327e-07 1.19527765e-08 5.24493327e-07 1.19528169e-08 5.24593327e-07 1.19527452e-08 5.24693327e-07 1.19528438e-08 5.24793327e-07 1.19527223e-08 5.24893327e-07 1.19528631e-08
+ 5.24993327e-07 1.19527059e-08 5.25093327e-07 1.19528765e-08 5.25193327e-07 1.1952695e-08 5.25293327e-07 1.19528855e-08 5.25393327e-07 1.19526882e-08 5.25493327e-07 1.19528903e-08 5.25593327e-07 1.19526846e-08 5.25693327e-07 1.19528927e-08
+ 5.25793327e-07 1.19526833e-08 5.25893327e-07 1.1952893e-08 5.25993327e-07 1.19526839e-08 5.26093327e-07 1.19528915e-08 5.26193327e-07 1.19526862e-08 5.26293327e-07 1.19528891e-08 5.26393327e-07 1.19526891e-08 5.26493327e-07 1.19528855e-08
+ 5.26593327e-07 1.19526932e-08 5.26693327e-07 1.19528813e-08 5.26793327e-07 1.19526976e-08 5.26893327e-07 1.19528767e-08 5.26993327e-07 1.19527022e-08 5.27093327e-07 1.19528718e-08 5.27193327e-07 1.19527071e-08 5.27293327e-07 1.19528671e-08
+ 5.27393327e-07 1.1952712e-08 5.27493327e-07 1.19528622e-08 5.27593327e-07 1.19527167e-08 5.27693327e-07 1.19528575e-08 5.27793327e-07 1.19527213e-08 5.27893327e-07 1.1952853e-08 5.27993327e-07 1.19527259e-08 5.28093327e-07 1.19528482e-08
+ 5.28193327e-07 1.19527306e-08 5.28293327e-07 1.19528439e-08 5.28393327e-07 1.19527351e-08 5.28493327e-07 1.19528397e-08 5.28593327e-07 1.19527388e-08 5.28693327e-07 1.1952836e-08 5.28793327e-07 1.19527425e-08 5.28893327e-07 1.19528322e-08
+ 5.28993327e-07 1.19527461e-08 5.29093327e-07 1.1952829e-08 5.29193327e-07 1.19527493e-08 5.29293327e-07 1.19528255e-08 5.29393327e-07 1.19527525e-08 5.29493327e-07 1.19528228e-08 5.29593327e-07 1.19527554e-08 5.29693327e-07 1.195282e-08
+ 5.29793327e-07 1.19527581e-08 5.29893327e-07 1.19528172e-08 5.29993327e-07 1.19527605e-08 5.30093327e-07 1.19528149e-08 5.30193327e-07 1.19527626e-08 5.30293327e-07 1.19528126e-08 5.30393327e-07 1.19527648e-08 5.30493327e-07 1.19528106e-08
+ 5.30593327e-07 1.19527669e-08 5.30693327e-07 1.19528088e-08 5.30793327e-07 1.19527684e-08 5.30893327e-07 1.19528072e-08 5.30993327e-07 1.19527701e-08 5.31093327e-07 1.19528055e-08 5.31193327e-07 1.19527719e-08 5.31293327e-07 1.19528042e-08
+ 5.31393327e-07 1.19527732e-08 5.31493327e-07 1.19528026e-08 5.31593327e-07 1.19527745e-08 5.31693327e-07 1.19528015e-08 5.31793327e-07 1.19527757e-08 5.31893327e-07 1.19528004e-08 5.31993327e-07 1.19527767e-08 5.32093327e-07 1.19527994e-08
+ 5.32193327e-07 1.19527778e-08 5.32293327e-07 1.19527984e-08 5.32393327e-07 1.19527787e-08 5.32493327e-07 1.19527973e-08 5.32593327e-07 1.19527794e-08 5.32693327e-07 1.19527966e-08 5.32793327e-07 1.19527803e-08 5.32893327e-07 1.19527959e-08
+ 5.32993327e-07 1.19527811e-08 5.33093327e-07 1.1952795e-08 5.33193327e-07 1.1952782e-08 5.33293327e-07 1.19527946e-08 5.33393327e-07 1.19527825e-08 5.33493327e-07 1.19527941e-08 5.33593327e-07 1.19527826e-08 5.33693327e-07 1.19527936e-08
+ 5.33793327e-07 1.1952783e-08 5.33893327e-07 1.19527932e-08 5.33993327e-07 1.19527835e-08 5.34093327e-07 1.19527928e-08 5.34193327e-07 1.1952784e-08 5.34293327e-07 1.19527923e-08 5.34393327e-07 1.19527843e-08 5.34493327e-07 1.19527923e-08
+ 5.34593327e-07 1.19527847e-08 5.34693327e-07 1.1952792e-08 5.34793327e-07 1.19527848e-08 5.34893327e-07 1.19527914e-08 5.34993327e-07 1.19527853e-08 5.35093327e-07 1.19527914e-08 5.35193327e-07 1.19527855e-08 5.35293327e-07 1.19527912e-08
+ 5.35393327e-07 1.19527858e-08 5.35493327e-07 1.19527907e-08 5.35593327e-07 1.19527862e-08 5.35693327e-07 1.19527905e-08 5.35793327e-07 1.19527865e-08 5.35893327e-07 1.19527901e-08 5.35993327e-07 1.19527865e-08 5.36093327e-07 1.19527902e-08
+ 5.36193327e-07 1.19527867e-08 5.36293327e-07 1.19527899e-08 5.36393327e-07 1.19527868e-08 5.36493327e-07 1.19527899e-08 5.36593327e-07 1.1952787e-08 5.36693327e-07 1.19527897e-08 5.36793327e-07 1.1952787e-08 5.36893327e-07 1.19527898e-08
+ 5.36993327e-07 1.1952787e-08 5.37093327e-07 1.19527894e-08 5.37193327e-07 1.1952787e-08 5.37293327e-07 1.19527897e-08 5.37393327e-07 1.1952787e-08 5.37493327e-07 1.19527897e-08 5.37593327e-07 1.19527871e-08 5.37693327e-07 1.19527895e-08
+ 5.37793327e-07 1.19527871e-08 5.37893327e-07 1.19527894e-08 5.37993327e-07 1.19527873e-08 5.38093327e-07 1.19527891e-08 5.38193327e-07 1.19527875e-08 5.38293327e-07 1.19527892e-08 5.38393327e-07 1.19527876e-08 5.38493327e-07 1.19527889e-08
+ 5.38593327e-07 1.19527878e-08 5.38693327e-07 1.19527891e-08 5.38793327e-07 1.19527878e-08 5.38893327e-07 1.19527889e-08 5.38993327e-07 1.19527879e-08 5.39093327e-07 1.19527891e-08 5.39193327e-07 1.19527879e-08 5.39293327e-07 1.1952789e-08
+ 5.39393327e-07 1.19527878e-08 5.39493327e-07 1.1952789e-08 5.39593327e-07 1.19527879e-08 5.39693327e-07 1.19527888e-08 5.39793327e-07 1.19527878e-08 5.39893327e-07 1.1952789e-08 5.39993327e-07 1.19527877e-08 5.40093327e-07 1.19527889e-08
+ 5.40193327e-07 1.19527877e-08 5.40293327e-07 1.19527888e-08 5.40393327e-07 1.19527879e-08 5.40493327e-07 1.19527889e-08 5.40593327e-07 1.19527878e-08 5.40693327e-07 1.19527888e-08 5.40793327e-07 1.19527878e-08 5.40893327e-07 1.19527891e-08
+ 5.40993327e-07 1.1952788e-08 5.41093327e-07 1.19527889e-08 5.41193327e-07 1.1952788e-08 5.41293327e-07 1.19527888e-08 5.41393327e-07 1.19527878e-08 5.41493327e-07 1.19527887e-08 5.41593327e-07 1.19527879e-08 5.41693327e-07 1.1952789e-08
+ 5.41793327e-07 1.1952788e-08 5.41893327e-07 1.19527888e-08 5.41993327e-07 1.19527881e-08 5.42093327e-07 1.19527888e-08 5.42193327e-07 1.19527878e-08 5.42293327e-07 1.19527886e-08 5.42393327e-07 1.19527879e-08 5.42493327e-07 1.19527886e-08
+ 5.42593327e-07 1.19527881e-08 5.42693327e-07 1.19527887e-08 5.42793327e-07 1.19527879e-08 5.42893327e-07 1.19527885e-08 5.42993327e-07 1.1952788e-08 5.43093327e-07 1.19527888e-08 5.43193327e-07 1.1952788e-08 5.43293327e-07 1.19527888e-08
+ 5.43393327e-07 1.19527879e-08 5.43493327e-07 1.19527884e-08 5.43593327e-07 1.19527879e-08 5.43693327e-07 1.19527885e-08 5.43793327e-07 1.19527879e-08 5.43893327e-07 1.19527885e-08 5.43993327e-07 1.19527878e-08 5.44093327e-07 1.19527884e-08
+ 5.44193327e-07 1.19527879e-08 5.44293327e-07 1.19527885e-08 5.44393327e-07 1.19527878e-08 5.44493327e-07 1.19527883e-08 5.44593327e-07 1.19527879e-08 5.44693327e-07 1.19527885e-08 5.44793327e-07 1.19527878e-08 5.44893327e-07 1.19527885e-08
+ 5.44993327e-07 1.19527881e-08 5.45093327e-07 1.19527886e-08 5.45193327e-07 1.19527878e-08 5.45293327e-07 1.19527885e-08 5.45393327e-07 1.19527879e-08 5.45493327e-07 1.19527885e-08 5.45593327e-07 1.19527878e-08 5.45693327e-07 1.19527884e-08
+ 5.45793327e-07 1.19527879e-08 5.45893327e-07 1.19527885e-08 5.45993327e-07 1.19527878e-08 5.46093327e-07 1.19527884e-08 5.46193327e-07 1.19527879e-08 5.46293327e-07 1.19527885e-08 5.46393327e-07 1.19527878e-08 5.46493327e-07 1.19527884e-08
+ 5.46593327e-07 1.19527879e-08 5.46693327e-07 1.19527885e-08 5.46793327e-07 1.19527878e-08 5.46893327e-07 1.19527884e-08 5.46993327e-07 1.19527879e-08 5.47093327e-07 1.19527885e-08 5.47193327e-07 1.19527878e-08 5.47293327e-07 1.19527884e-08
+ 5.47393327e-07 1.19527879e-08 5.47493327e-07 1.19527885e-08 5.47593327e-07 1.19527878e-08 5.47693327e-07 1.19527884e-08 5.47793327e-07 1.19527879e-08 5.47893327e-07 1.19527885e-08 5.47993327e-07 1.19527878e-08 5.48093327e-07 1.19527884e-08
+ 5.48193327e-07 1.19527879e-08 5.48293327e-07 1.19527885e-08 5.48393327e-07 1.19527878e-08 5.48493327e-07 1.19527884e-08 5.48593327e-07 1.19527879e-08 5.48693327e-07 1.19527885e-08 5.48793327e-07 1.19527878e-08 5.48893327e-07 1.19527884e-08
+ 5.48993327e-07 1.19527879e-08 5.49093327e-07 1.19527885e-08 5.49193327e-07 1.19527878e-08 5.49293327e-07 1.19527884e-08 5.49393327e-07 1.19527879e-08 5.49493327e-07 1.19527885e-08 5.49593327e-07 1.19527878e-08 5.49693327e-07 1.19527885e-08
+ 5.49793327e-07 1.1952788e-08 5.49893327e-07 1.19527887e-08 5.49993327e-07 1.19527882e-08 5.50093327e-07 1.19527887e-08 5.50193327e-07 1.19527882e-08 5.50293327e-07 1.19527885e-08 5.50393327e-07 1.19527881e-08 5.50493327e-07 1.19527882e-08
+ 5.50593327e-07 1.19527881e-08 5.50693327e-07 1.19527883e-08 5.50793327e-07 1.19527881e-08 5.50893327e-07 1.19527883e-08 5.50993327e-07 1.19527881e-08 5.51e-07 1.19527885e-08 5.5101e-07 1.19399427e-08 5.5103e-07 1.20150115e-08
+ 5.5107e-07 1.18559377e-08 5.5115e-07 1.20621028e-08 5.5125e-07 1.18410989e-08 5.5135e-07 1.20574877e-08 5.5145e-07 1.1863822e-08 5.5155e-07 1.20197035e-08 5.5165e-07 1.1910158e-08 5.5175e-07 1.19686131e-08
+ 5.5185e-07 1.19674862e-08 5.51930828e-07 1.83418271e-07 5.52e-07 1.06002517e-07 5.52008608e-07 -6.35218173e-06 5.52025825e-07 -6.40058733e-06 5.52060258e-07 9.75152962e-06 5.52106188e-07 5.28435492e-06 5.52150118e-07 -1.51923671e-05
+ 5.5219811e-07 6.42629664e-06 5.52255501e-07 9.57222351e-07 5.52312176e-07 -1.57314433e-06 5.52404431e-07 1.13652367e-06 5.52490774e-07 -1.00482103e-06 5.52590774e-07 9.71186727e-07 5.52690774e-07 -8.68547259e-07 5.52790774e-07 8.16808096e-07
+ 5.52890774e-07 -7.24287651e-07 5.52990774e-07 6.88965999e-07 5.53090774e-07 -6.14052292e-07 5.53190774e-07 5.94787164e-07 5.53290774e-07 -5.33642225e-07 5.53390774e-07 5.25529847e-07 5.53490774e-07 -4.73285723e-07 5.53590774e-07 4.7203629e-07
+ 5.53690774e-07 -4.25085269e-07 5.53790774e-07 4.27835408e-07 5.53890774e-07 -3.83953564e-07 5.53990774e-07 3.89048055e-07 5.54090774e-07 -3.4701833e-07 5.54190774e-07 3.53603079e-07 5.54290774e-07 -3.12840629e-07 5.54390774e-07 3.20537789e-07
+ 5.54490774e-07 -2.80809747e-07 5.54590774e-07 2.89491019e-07 5.54690774e-07 -2.50738347e-07 5.54790774e-07 2.60389507e-07 5.54890774e-07 -2.22624131e-07 5.54990774e-07 2.33269734e-07 5.55090774e-07 -1.96520033e-07 5.55190774e-07 2.08185539e-07
+ 5.55290774e-07 -1.72470285e-07 5.55390774e-07 1.85165182e-07 5.55490774e-07 -1.50484079e-07 5.55590774e-07 1.64198319e-07 5.55690774e-07 -1.30531642e-07 5.55790774e-07 1.45236542e-07 5.55890774e-07 -1.12547054e-07 5.55990774e-07 1.28198329e-07
+ 5.56090774e-07 -9.64351095e-08 5.56190774e-07 1.12976947e-07 5.56290774e-07 -8.20795775e-08 5.56390774e-07 9.94489937e-08 5.56490774e-07 -6.93520125e-08 5.56590774e-07 8.74825733e-08 5.56690774e-07 -5.81182253e-08 5.56790774e-07 7.69425248e-08
+ 5.56890774e-07 -4.82432947e-08 5.56990774e-07 6.76957224e-08 5.57090774e-07 -3.959732e-08 5.57190774e-07 5.96159694e-08 5.57290774e-07 -3.20580335e-08 5.57390774e-07 5.2583098e-08 5.57490774e-07 -2.55059463e-08 5.57590774e-07 4.64804055e-08
+ 5.57690774e-07 -1.98288253e-08 5.57790774e-07 4.1200075e-08 5.57890774e-07 -1.49233088e-08 5.57990774e-07 3.66432218e-08 5.58090774e-07 -1.06952402e-08 5.58190774e-07 3.27205768e-08 5.58290774e-07 -7.06015083e-09 5.58390774e-07 2.93521472e-08
+ 5.58490774e-07 -3.94241775e-09 5.58590774e-07 2.64666448e-08 5.58690774e-07 -1.27496946e-09 5.58790774e-07 2.4000838e-08 5.58890774e-07 9.95357963e-10 5.58990774e-07 2.19105883e-08 5.59090774e-07 2.91112168e-09 5.59190774e-07 2.01552989e-08
+ 5.59290774e-07 4.51850521e-09 5.59390774e-07 1.86841679e-08 5.59490774e-07 5.86417118e-09 5.59590774e-07 1.74539928e-08 5.59690774e-07 6.98806962e-09 5.59790774e-07 1.64278643e-08 5.59890774e-07 7.92430507e-09 5.59990774e-07 1.55742175e-08
+ 5.60090774e-07 8.70212047e-09 5.60190774e-07 1.48659897e-08 5.60290774e-07 9.34652492e-09 5.60390774e-07 1.42800906e-08 5.60490774e-07 9.87882104e-09 5.60590774e-07 1.37968806e-08 5.60690774e-07 1.03171052e-08 5.60790774e-07 1.33996929e-08
+ 5.60890774e-07 1.06767188e-08 5.60990774e-07 1.30744149e-08 5.61090774e-07 1.09706387e-08 5.61190774e-07 1.28091175e-08 5.61290774e-07 1.1209824e-08 5.61390774e-07 1.25937394e-08 5.61490774e-07 1.14035098e-08 5.61590774e-07 1.24198065e-08
+ 5.61690774e-07 1.15594666e-08 5.61790774e-07 1.22801992e-08 5.61890774e-07 1.16842192e-08 5.61990774e-07 1.21689275e-08 5.62090774e-07 1.1783264e-08 5.62190774e-07 1.20809674e-08 5.62290774e-07 1.1861181e-08 5.62390774e-07 1.20121454e-08
+ 5.62490774e-07 1.19217766e-08 5.62590774e-07 1.19589735e-08 5.62690774e-07 1.19682666e-08 5.62790774e-07 1.19184841e-08 5.62890774e-07 1.20033725e-08 5.62990774e-07 1.18882069e-08 5.63090774e-07 1.20293195e-08 5.63190774e-07 1.18661405e-08
+ 5.63290774e-07 1.20479116e-08 5.63390774e-07 1.1850656e-08 5.63490774e-07 1.20606221e-08 5.63590774e-07 1.18404172e-08 5.63690774e-07 1.20686623e-08 5.63790774e-07 1.18343279e-08 5.63890774e-07 1.20729713e-08 5.63990774e-07 1.18315197e-08
+ 5.64090774e-07 1.20748511e-08 5.64190774e-07 1.18303283e-08 5.64290774e-07 1.20750054e-08 5.64390774e-07 1.18314565e-08 5.64490774e-07 1.20727117e-08 5.64590774e-07 1.18346005e-08 5.64690774e-07 1.20690052e-08 5.64790774e-07 1.18387675e-08
+ 5.64890774e-07 1.20644241e-08 5.64990774e-07 1.18436872e-08 5.65090774e-07 1.20592382e-08 5.65190774e-07 1.1849077e-08 5.65290774e-07 1.20536968e-08 5.65390774e-07 1.18547525e-08 5.65490774e-07 1.20478535e-08 5.65590774e-07 1.18607524e-08
+ 5.65690774e-07 1.20418265e-08 5.65790774e-07 1.18666782e-08 5.65890774e-07 1.20360327e-08 5.65990774e-07 1.18723564e-08 5.66090774e-07 1.20304578e-08 5.66190774e-07 1.18778301e-08 5.66290774e-07 1.20250903e-08 5.66390774e-07 1.18830854e-08
+ 5.66490774e-07 1.20199509e-08 5.66590774e-07 1.18881048e-08 5.66690774e-07 1.20150554e-08 5.66790774e-07 1.18928744e-08 5.66890774e-07 1.20104132e-08 5.66990774e-07 1.18973873e-08 5.67090774e-07 1.20060307e-08 5.67190774e-07 1.19016378e-08
+ 5.67290774e-07 1.20019122e-08 5.67390774e-07 1.1905626e-08 5.67490774e-07 1.19980544e-08 5.67590774e-07 1.19093532e-08 5.67690774e-07 1.19944567e-08 5.67790774e-07 1.19128237e-08 5.67890774e-07 1.19911097e-08 5.67990774e-07 1.1916051e-08
+ 5.68090774e-07 1.19879989e-08 5.68190774e-07 1.19190478e-08 5.68290774e-07 1.19851135e-08 5.68390774e-07 1.19218413e-08 5.68490774e-07 1.19823907e-08 5.68590774e-07 1.19244633e-08 5.68690774e-07 1.197991e-08 5.68790774e-07 1.19268156e-08
+ 5.68890774e-07 1.19776579e-08 5.68990774e-07 1.19289786e-08 5.69090774e-07 1.19755774e-08 5.69190774e-07 1.19309846e-08 5.69290774e-07 1.19736417e-08 5.69390774e-07 1.19328462e-08 5.69490774e-07 1.19718589e-08 5.69590774e-07 1.19345514e-08
+ 5.69690774e-07 1.19702255e-08 5.69790774e-07 1.19361175e-08 5.69890774e-07 1.19687259e-08 5.69990774e-07 1.19375512e-08 5.70090774e-07 1.19673552e-08 5.70190774e-07 1.19388627e-08 5.70290774e-07 1.19661001e-08 5.70390774e-07 1.19400644e-08
+ 5.70490774e-07 1.19649494e-08 5.70590774e-07 1.19411659e-08 5.70690774e-07 1.1963895e-08 5.70790774e-07 1.19421752e-08 5.70890774e-07 1.19629286e-08 5.70990774e-07 1.19431e-08 5.71090774e-07 1.19620443e-08 5.71190774e-07 1.19439457e-08
+ 5.71290774e-07 1.19612352e-08 5.71390774e-07 1.19447196e-08 5.71490774e-07 1.19604955e-08 5.71590774e-07 1.19454266e-08 5.71690774e-07 1.19598198e-08 5.71790774e-07 1.1946072e-08 5.71890774e-07 1.19592034e-08 5.71990774e-07 1.19466611e-08
+ 5.72090774e-07 1.19586407e-08 5.72190774e-07 1.19471981e-08 5.72290774e-07 1.19581275e-08 5.72390774e-07 1.19476888e-08 5.72490774e-07 1.19576589e-08 5.72590774e-07 1.19481365e-08 5.72690774e-07 1.19572315e-08 5.72790774e-07 1.19485446e-08
+ 5.72890774e-07 1.19568415e-08 5.72990774e-07 1.19489169e-08 5.73090774e-07 1.19564855e-08 5.73190774e-07 1.19492571e-08 5.73290774e-07 1.195616e-08 5.73390774e-07 1.19495683e-08 5.73490774e-07 1.19558631e-08 5.73590774e-07 1.19498513e-08
+ 5.73690774e-07 1.19555934e-08 5.73790774e-07 1.19501089e-08 5.73890774e-07 1.19553473e-08 5.73990774e-07 1.19503444e-08 5.74090774e-07 1.19551221e-08 5.74190774e-07 1.19505598e-08 5.74290774e-07 1.1954916e-08 5.74390774e-07 1.19507567e-08
+ 5.74490774e-07 1.19547276e-08 5.74590774e-07 1.19509369e-08 5.74690774e-07 1.19545556e-08 5.74790774e-07 1.19511012e-08 5.74890774e-07 1.19543982e-08 5.74990774e-07 1.19512519e-08 5.75090774e-07 1.19542544e-08 5.75190774e-07 1.19513892e-08
+ 5.75290774e-07 1.19541231e-08 5.75390774e-07 1.19515147e-08 5.75490774e-07 1.19540033e-08 5.75590774e-07 1.19516284e-08 5.75690774e-07 1.19538953e-08 5.75790774e-07 1.19517322e-08 5.75890774e-07 1.1953796e-08 5.75990774e-07 1.19518267e-08
+ 5.76090774e-07 1.19537056e-08 5.76190774e-07 1.19519136e-08 5.76290774e-07 1.19536225e-08 5.76390774e-07 1.1951993e-08 5.76490774e-07 1.19535467e-08 5.76590774e-07 1.19520653e-08 5.76690774e-07 1.19534775e-08 5.76790774e-07 1.19521313e-08
+ 5.76890774e-07 1.19534143e-08 5.76990774e-07 1.19521916e-08 5.77090774e-07 1.19533566e-08 5.77190774e-07 1.19522467e-08 5.77290774e-07 1.19533045e-08 5.77390774e-07 1.19522967e-08 5.77490774e-07 1.1953257e-08 5.77590774e-07 1.19523422e-08
+ 5.77690774e-07 1.19532133e-08 5.77790774e-07 1.19523836e-08 5.77890774e-07 1.19531738e-08 5.77990774e-07 1.19524212e-08 5.78090774e-07 1.19531379e-08 5.78190774e-07 1.19524554e-08 5.78290774e-07 1.1953105e-08 5.78390774e-07 1.19524866e-08
+ 5.78490774e-07 1.19530754e-08 5.78590774e-07 1.19525148e-08 5.78690774e-07 1.19530485e-08 5.78790774e-07 1.19525404e-08 5.78890774e-07 1.19530241e-08 5.78990774e-07 1.19525635e-08 5.79090774e-07 1.19530022e-08 5.79190774e-07 1.19525844e-08
+ 5.79290774e-07 1.19529827e-08 5.79390774e-07 1.19526031e-08 5.79490774e-07 1.19529645e-08 5.79590774e-07 1.19526204e-08 5.79690774e-07 1.19529481e-08 5.79790774e-07 1.19526362e-08 5.79890774e-07 1.19529332e-08 5.79990774e-07 1.19526502e-08
+ 5.80090774e-07 1.19529197e-08 5.80190774e-07 1.19526631e-08 5.80290774e-07 1.19529075e-08 5.80390774e-07 1.19526747e-08 5.80490774e-07 1.19528965e-08 5.80590774e-07 1.19526853e-08 5.80690774e-07 1.19528864e-08 5.80790774e-07 1.19526949e-08
+ 5.80890774e-07 1.19528773e-08 5.80990774e-07 1.19527034e-08 5.81090774e-07 1.19528691e-08 5.81190774e-07 1.19527112e-08 5.81290774e-07 1.19528617e-08 5.81390774e-07 1.19527183e-08 5.81490774e-07 1.1952855e-08 5.81590774e-07 1.19527247e-08
+ 5.81690774e-07 1.19528489e-08 5.81790774e-07 1.19527304e-08 5.81890774e-07 1.19528434e-08 5.81990774e-07 1.19527359e-08 5.82090774e-07 1.19528384e-08 5.82190774e-07 1.19527405e-08 5.82290774e-07 1.19528337e-08 5.82390774e-07 1.19527447e-08
+ 5.82490774e-07 1.19528299e-08 5.82590774e-07 1.19527487e-08 5.82690774e-07 1.19528258e-08 5.82790774e-07 1.19527524e-08 5.82890774e-07 1.19528226e-08 5.82990774e-07 1.19527553e-08 5.83090774e-07 1.19528197e-08 5.83190774e-07 1.19527588e-08
+ 5.83290774e-07 1.19528165e-08 5.83390774e-07 1.19527615e-08 5.83490774e-07 1.19528138e-08 5.83590774e-07 1.19527638e-08 5.83690774e-07 1.19528115e-08 5.83790774e-07 1.19527657e-08 5.83890774e-07 1.19528096e-08 5.83990774e-07 1.1952768e-08
+ 5.84090774e-07 1.19528078e-08 5.84190774e-07 1.19527698e-08 5.84290774e-07 1.1952806e-08 5.84390774e-07 1.19527715e-08 5.84490774e-07 1.19528044e-08 5.84590774e-07 1.19527728e-08 5.84690774e-07 1.19528029e-08 5.84790774e-07 1.19527741e-08
+ 5.84890774e-07 1.19528017e-08 5.84990774e-07 1.19527755e-08 5.85090774e-07 1.19528005e-08 5.85190774e-07 1.19527765e-08 5.85290774e-07 1.19527996e-08 5.85390774e-07 1.19527776e-08 5.85490774e-07 1.19527986e-08 5.85590774e-07 1.19527786e-08
+ 5.85690774e-07 1.19527976e-08 5.85790774e-07 1.19527793e-08 5.85890774e-07 1.19527968e-08 5.85990774e-07 1.19527802e-08 5.86090774e-07 1.19527959e-08 5.86190774e-07 1.19527809e-08 5.86290774e-07 1.19527953e-08 5.86390774e-07 1.19527815e-08
+ 5.86490774e-07 1.19527948e-08 5.86590774e-07 1.19527823e-08 5.86690774e-07 1.19527941e-08 5.86790774e-07 1.1952783e-08 5.86890774e-07 1.19527936e-08 5.86990774e-07 1.19527832e-08 5.87090774e-07 1.19527931e-08 5.87190774e-07 1.19527835e-08
+ 5.87290774e-07 1.19527927e-08 5.87390774e-07 1.19527839e-08 5.87490774e-07 1.19527923e-08 5.87590774e-07 1.19527844e-08 5.87690774e-07 1.1952792e-08 5.87790774e-07 1.19527847e-08 5.87890774e-07 1.19527917e-08 5.87990774e-07 1.19527851e-08
+ 5.88090774e-07 1.19527917e-08 5.88190774e-07 1.19527853e-08 5.88290774e-07 1.19527913e-08 5.88390774e-07 1.19527856e-08 5.88490774e-07 1.1952791e-08 5.88590774e-07 1.19527857e-08 5.88690774e-07 1.19527908e-08 5.88790774e-07 1.1952786e-08
+ 5.88890774e-07 1.19527905e-08 5.88990774e-07 1.19527863e-08 5.89090774e-07 1.19527903e-08 5.89190774e-07 1.19527864e-08 5.89290774e-07 1.19527903e-08 5.89390774e-07 1.19527865e-08 5.89490774e-07 1.19527901e-08 5.89590774e-07 1.19527868e-08
+ 5.89690774e-07 1.19527898e-08 5.89790774e-07 1.19527868e-08 5.89890774e-07 1.19527899e-08 5.89990774e-07 1.19527868e-08 5.90090774e-07 1.19527898e-08 5.90190774e-07 1.19527869e-08 5.90290774e-07 1.19527897e-08 5.90390774e-07 1.19527869e-08
+ 5.90490774e-07 1.19527898e-08 5.90590774e-07 1.1952787e-08 5.90690774e-07 1.19527896e-08 5.90790774e-07 1.19527871e-08 5.90890774e-07 1.19527894e-08 5.90990774e-07 1.19527871e-08 5.91090774e-07 1.19527893e-08 5.91190774e-07 1.19527873e-08
+ 5.91290774e-07 1.19527893e-08 5.91390774e-07 1.19527874e-08 5.91490774e-07 1.19527893e-08 5.91590774e-07 1.19527875e-08 5.91690774e-07 1.1952789e-08 5.91790774e-07 1.19527875e-08 5.91890774e-07 1.1952789e-08 5.91990774e-07 1.19527876e-08
+ 5.92090774e-07 1.19527891e-08 5.92190774e-07 1.19527876e-08 5.92290774e-07 1.19527889e-08 5.92390774e-07 1.19527878e-08 5.92490774e-07 1.19527889e-08 5.92590774e-07 1.1952788e-08 5.92690774e-07 1.19527888e-08 5.92790774e-07 1.19527881e-08
+ 5.92890774e-07 1.19527887e-08 5.92990774e-07 1.19527882e-08 5.93090774e-07 1.19527883e-08 5.93190774e-07 1.19527878e-08 5.93290774e-07 1.19527885e-08 5.93390774e-07 1.1952788e-08 5.93490774e-07 1.19527883e-08 5.93590774e-07 1.19527879e-08
+ 5.93690774e-07 1.19527884e-08 5.93790774e-07 1.19527879e-08 5.93890774e-07 1.19527885e-08 5.93990774e-07 1.19527878e-08 5.94090774e-07 1.19527885e-08 5.94190774e-07 1.1952788e-08 5.94290774e-07 1.19527888e-08 5.94390774e-07 1.19527881e-08
+ 5.94490774e-07 1.19527888e-08 5.94590774e-07 1.19527881e-08 5.94690774e-07 1.19527886e-08 5.94790774e-07 1.19527881e-08 5.94890774e-07 1.19527887e-08 5.94990774e-07 1.1952788e-08 5.95090774e-07 1.19527888e-08 5.95190774e-07 1.1952788e-08
+ 5.95290774e-07 1.19527887e-08 5.95390774e-07 1.19527879e-08 5.95490774e-07 1.19527886e-08 5.95590774e-07 1.19527881e-08 5.95690774e-07 1.19527887e-08 5.95790774e-07 1.1952788e-08 5.95890774e-07 1.19527885e-08 5.95990774e-07 1.19527881e-08
+ 5.96090774e-07 1.19527888e-08 5.96190774e-07 1.19527881e-08 5.96290774e-07 1.19527886e-08 5.96390774e-07 1.1952788e-08 5.96490774e-07 1.19527888e-08 5.96590774e-07 1.19527881e-08 5.96690774e-07 1.19527886e-08 5.96790774e-07 1.1952788e-08
+ 5.96890774e-07 1.19527883e-08 5.96990774e-07 1.19527879e-08 5.97090774e-07 1.19527883e-08 5.97190774e-07 1.1952788e-08 5.97290774e-07 1.19527883e-08 5.97390774e-07 1.1952788e-08 5.97490774e-07 1.19527882e-08 5.97590774e-07 1.1952788e-08
+ 5.97690774e-07 1.19527883e-08 5.97790774e-07 1.1952788e-08 5.97890774e-07 1.19527883e-08 5.97990774e-07 1.1952788e-08 5.98090774e-07 1.19527884e-08 5.98190774e-07 1.1952788e-08 5.98290774e-07 1.19527883e-08 5.98390774e-07 1.19527881e-08
+ 5.98490774e-07 1.19527883e-08 5.98590774e-07 1.1952788e-08 5.98690774e-07 1.19527884e-08 5.98790774e-07 1.19527879e-08 5.98890774e-07 1.19527885e-08 5.98990774e-07 1.1952788e-08 5.99090774e-07 1.19527884e-08 5.99190774e-07 1.19527881e-08
+ 5.99290774e-07 1.19527883e-08 5.99390774e-07 1.1952788e-08 5.99490774e-07 1.19527885e-08 5.99590774e-07 1.19527879e-08 5.99690774e-07 1.19527885e-08 5.99790774e-07 1.19527881e-08 5.99890774e-07 1.19527882e-08 5.99990774e-07 1.19527881e-08
+ 6e-07 1.19527881e-08 6.0001e-07 1.19810075e-08 6.0003e-07 1.18152684e-08 6.0007e-07 1.21656673e-08 6.0015e-07 1.17141754e-08 6.0025e-07 1.21973735e-08 6.0035e-07 1.17166006e-08 6.0045e-07 1.21670028e-08
+ 6.0055e-07 1.17775964e-08 6.0065e-07 1.18484739e-08 6.0075e-07 2.53191131e-08 6.0085e-07 -4.04759482e-07 6.00932239e-07 6.49708168e-06 6.01e-07 -4.94343878e-05 6.01008502e-07 -5.0992026e-05 6.01025505e-07 -4.39145059e-05
+ 6.01059511e-07 -1.62206912e-05 6.01090728e-07 0.000285043155 6.01143656e-07 0.000513849787 6.01199398e-07 0.00155348227 6.01276452e-07 -0.0180250591 6.01342062e-07 -0.00339007548 6.01411951e-07 3.25710063 6.01487979e-07 4.90275261
+ 6.01566956e-07 5.02684152 6.01643585e-07 4.98988775 6.01743585e-07 5.00539209 6.01843585e-07 4.99682771 6.01943585e-07 5.00195612 6.02043585e-07 4.99873104 6.02143585e-07 5.00083562 6.02243585e-07 4.99943657
+ 6.02343585e-07 5.00037969 6.02443585e-07 4.99974066 6.02543585e-07 5.00017605 6.02643585e-07 4.99987923 6.02743585e-07 5.00008215 6.02843585e-07 4.99994356 6.02943585e-07 5.00003839 6.03043585e-07 4.9999736
+ 6.03143585e-07 5.00001792 6.03243585e-07 4.99998767 6.03343585e-07 5.00000832 6.03443585e-07 4.99999427 6.03543585e-07 5.00000382 6.03643585e-07 4.99999736 6.03743585e-07 5.00000171 6.03843585e-07 4.99999881
+ 6.03943585e-07 5.00000073 6.04043585e-07 4.99999949 6.04143585e-07 5.00000027 6.04243585e-07 4.9999998 6.04343585e-07 5.00000006 6.04443585e-07 4.99999994 6.04543585e-07 4.99999996 6.04643585e-07 5.0
+ 6.04743585e-07 4.99999993 6.04843585e-07 5.00000002 6.04943585e-07 4.99999992 6.05043585e-07 5.00000003 6.05143585e-07 4.99999992 6.05243585e-07 5.00000003 6.05343585e-07 4.99999992 6.05443585e-07 5.00000002
+ 6.05543585e-07 4.99999993 6.05643585e-07 5.00000001 6.05743585e-07 4.99999993 6.05843585e-07 5.00000001 6.05943585e-07 4.99999994 6.06043585e-07 5.0 6.06143585e-07 4.99999994 6.06243585e-07 5.0
+ 6.06343585e-07 4.99999995 6.06443585e-07 4.99999999 6.06543585e-07 4.99999995 6.06643585e-07 4.99999999 6.06743585e-07 4.99999996 6.06843585e-07 4.99999999 6.06943585e-07 4.99999996 6.07043585e-07 4.99999998
+ 6.07143585e-07 4.99999996 6.07243585e-07 4.99999998 6.07343585e-07 4.99999996 6.07443585e-07 4.99999998 6.07543585e-07 4.99999996 6.07643585e-07 4.99999998 6.07743585e-07 4.99999997 6.07843585e-07 4.99999998
+ 6.07943585e-07 4.99999997 6.08043585e-07 4.99999998 6.08143585e-07 4.99999997 6.08243585e-07 4.99999998 6.08343585e-07 4.99999997 6.08443585e-07 4.99999998 6.08543585e-07 4.99999997 6.08643585e-07 4.99999997
+ 6.08743585e-07 4.99999997 6.08843585e-07 4.99999997 6.08943585e-07 4.99999997 6.09043585e-07 4.99999997 6.09143585e-07 4.99999997 6.09243585e-07 4.99999997 6.09343585e-07 4.99999997 6.09443585e-07 4.99999997
+ 6.09543585e-07 4.99999997 6.09643585e-07 4.99999997 6.09743585e-07 4.99999997 6.09843585e-07 4.99999997 6.09943585e-07 4.99999997 6.10043585e-07 4.99999997 6.10143585e-07 4.99999997 6.10243585e-07 4.99999997
+ 6.10343585e-07 4.99999997 6.10443585e-07 4.99999997 6.10543585e-07 4.99999997 6.10643585e-07 4.99999997 6.10743585e-07 4.99999997 6.10843585e-07 4.99999997 6.10943585e-07 4.99999997 6.11043585e-07 4.99999997
+ 6.11143585e-07 4.99999997 6.11243585e-07 4.99999997 6.11343585e-07 4.99999997 6.11443585e-07 4.99999997 6.11543585e-07 4.99999997 6.11643585e-07 4.99999997 6.11743585e-07 4.99999997 6.11843585e-07 4.99999997
+ 6.11943585e-07 4.99999997 6.12043585e-07 4.99999997 6.12143585e-07 4.99999997 6.12243585e-07 4.99999997 6.12343585e-07 4.99999997 6.12443585e-07 4.99999997 6.12543585e-07 4.99999997 6.12643585e-07 4.99999997
+ 6.12743585e-07 4.99999997 6.12843585e-07 4.99999997 6.12943585e-07 4.99999997 6.13043585e-07 4.99999997 6.13143585e-07 4.99999997 6.13243585e-07 4.99999997 6.13343585e-07 4.99999997 6.13443585e-07 4.99999997
+ 6.13543585e-07 4.99999997 6.13643585e-07 4.99999997 6.13743585e-07 4.99999997 6.13843585e-07 4.99999997 6.13943585e-07 4.99999997 6.14043585e-07 4.99999997 6.14143585e-07 4.99999997 6.14243585e-07 4.99999997
+ 6.14343585e-07 4.99999997 6.14443585e-07 4.99999997 6.14543585e-07 4.99999997 6.14643585e-07 4.99999997 6.14743585e-07 4.99999997 6.14843585e-07 4.99999997 6.14943585e-07 4.99999997 6.15043585e-07 4.99999997
+ 6.15143585e-07 4.99999997 6.15243585e-07 4.99999997 6.15343585e-07 4.99999997 6.15443585e-07 4.99999997 6.15543585e-07 4.99999997 6.15643585e-07 4.99999997 6.15743585e-07 4.99999997 6.15843585e-07 4.99999997
+ 6.15943585e-07 4.99999997 6.16043585e-07 4.99999997 6.16143585e-07 4.99999997 6.16243585e-07 4.99999997 6.16343585e-07 4.99999997 6.16443585e-07 4.99999997 6.16543585e-07 4.99999997 6.16643585e-07 4.99999997
+ 6.16743585e-07 4.99999997 6.16843585e-07 4.99999997 6.16943585e-07 4.99999997 6.17043585e-07 4.99999997 6.17143585e-07 4.99999997 6.17243585e-07 4.99999997 6.17343585e-07 4.99999997 6.17443585e-07 4.99999997
+ 6.17543585e-07 4.99999997 6.17643585e-07 4.99999997 6.17743585e-07 4.99999997 6.17843585e-07 4.99999997 6.17943585e-07 4.99999997 6.18043585e-07 4.99999997 6.18143585e-07 4.99999997 6.18243585e-07 4.99999997
+ 6.18343585e-07 4.99999997 6.18443585e-07 4.99999997 6.18543585e-07 4.99999997 6.18643585e-07 4.99999997 6.18743585e-07 4.99999997 6.18843585e-07 4.99999997 6.18943585e-07 4.99999997 6.19043585e-07 4.99999997
+ 6.19143585e-07 4.99999997 6.19243585e-07 4.99999997 6.19343585e-07 4.99999997 6.19443585e-07 4.99999997 6.19543585e-07 4.99999997 6.19643585e-07 4.99999997 6.19743585e-07 4.99999997 6.19843585e-07 4.99999997
+ 6.19943585e-07 4.99999997 6.20043585e-07 4.99999997 6.20143585e-07 4.99999997 6.20243585e-07 4.99999997 6.20343585e-07 4.99999997 6.20443585e-07 4.99999997 6.20543585e-07 4.99999997 6.20643585e-07 4.99999997
+ 6.20743585e-07 4.99999997 6.20843585e-07 4.99999997 6.20943585e-07 4.99999997 6.21043585e-07 4.99999997 6.21143585e-07 4.99999997 6.21243585e-07 4.99999997 6.21343585e-07 4.99999997 6.21443585e-07 4.99999997
+ 6.21543585e-07 4.99999997 6.21643585e-07 4.99999997 6.21743585e-07 4.99999997 6.21843585e-07 4.99999997 6.21943585e-07 4.99999997 6.22043585e-07 4.99999997 6.22143585e-07 4.99999997 6.22243585e-07 4.99999997
+ 6.22343585e-07 4.99999997 6.22443585e-07 4.99999997 6.22543585e-07 4.99999997 6.22643585e-07 4.99999997 6.22743585e-07 4.99999997 6.22843585e-07 4.99999997 6.22943585e-07 4.99999997 6.23043585e-07 4.99999997
+ 6.23143585e-07 4.99999997 6.23243585e-07 4.99999997 6.23343585e-07 4.99999997 6.23443585e-07 4.99999997 6.23543585e-07 4.99999997 6.23643585e-07 4.99999997 6.23743585e-07 4.99999997 6.23843585e-07 4.99999997
+ 6.23943585e-07 4.99999997 6.24043585e-07 4.99999997 6.24143585e-07 4.99999997 6.24243585e-07 4.99999997 6.24343585e-07 4.99999997 6.24443585e-07 4.99999997 6.24543585e-07 4.99999997 6.24643585e-07 4.99999997
+ 6.24743585e-07 4.99999997 6.24843585e-07 4.99999997 6.24943585e-07 4.99999997 6.25043585e-07 4.99999997 6.25143585e-07 4.99999997 6.25243585e-07 4.99999997 6.25343585e-07 4.99999997 6.25443585e-07 4.99999997
+ 6.25543585e-07 4.99999997 6.25643585e-07 4.99999997 6.25743585e-07 4.99999997 6.25843585e-07 4.99999997 6.25943585e-07 4.99999997 6.26043585e-07 4.99999997 6.26143585e-07 4.99999997 6.26243585e-07 4.99999997
+ 6.26343585e-07 4.99999997 6.26443585e-07 4.99999997 6.26543585e-07 4.99999997 6.26643585e-07 4.99999997 6.26743585e-07 4.99999997 6.26843585e-07 4.99999997 6.26943585e-07 4.99999997 6.27043585e-07 4.99999997
+ 6.27143585e-07 4.99999997 6.27243585e-07 4.99999997 6.27343585e-07 4.99999997 6.27443585e-07 4.99999997 6.27543585e-07 4.99999997 6.27643585e-07 4.99999997 6.27743585e-07 4.99999997 6.27843585e-07 4.99999997
+ 6.27943585e-07 4.99999997 6.28043585e-07 4.99999997 6.28143585e-07 4.99999997 6.28243585e-07 4.99999997 6.28343585e-07 4.99999997 6.28443585e-07 4.99999997 6.28543585e-07 4.99999997 6.28643585e-07 4.99999997
+ 6.28743585e-07 4.99999997 6.28843585e-07 4.99999997 6.28943585e-07 4.99999997 6.29043585e-07 4.99999997 6.29143585e-07 4.99999997 6.29243585e-07 4.99999997 6.29343585e-07 4.99999997 6.29443585e-07 4.99999997
+ 6.29543585e-07 4.99999997 6.29643585e-07 4.99999997 6.29743585e-07 4.99999997 6.29843585e-07 4.99999997 6.29943585e-07 4.99999997 6.30043585e-07 4.99999997 6.30143585e-07 4.99999997 6.30243585e-07 4.99999997
+ 6.30343585e-07 4.99999997 6.30443585e-07 4.99999997 6.30543585e-07 4.99999997 6.30643585e-07 4.99999997 6.30743585e-07 4.99999997 6.30843585e-07 4.99999997 6.30943585e-07 4.99999997 6.31043585e-07 4.99999997
+ 6.31143585e-07 4.99999997 6.31243585e-07 4.99999997 6.31343585e-07 4.99999997 6.31443585e-07 4.99999997 6.31543585e-07 4.99999997 6.31643585e-07 4.99999997 6.31743585e-07 4.99999997 6.31843585e-07 4.99999997
+ 6.31943585e-07 4.99999997 6.32043585e-07 4.99999997 6.32143585e-07 4.99999997 6.32243585e-07 4.99999997 6.32343585e-07 4.99999997 6.32443585e-07 4.99999997 6.32543585e-07 4.99999997 6.32643585e-07 4.99999997
+ 6.32743585e-07 4.99999997 6.32843585e-07 4.99999997 6.32943585e-07 4.99999997 6.33043585e-07 4.99999997 6.33143585e-07 4.99999997 6.33243585e-07 4.99999997 6.33343585e-07 4.99999997 6.33443585e-07 4.99999997
+ 6.33543585e-07 4.99999997 6.33643585e-07 4.99999997 6.33743585e-07 4.99999997 6.33843585e-07 4.99999997 6.33943585e-07 4.99999997 6.34043585e-07 4.99999997 6.34143585e-07 4.99999997 6.34243585e-07 4.99999997
+ 6.34343585e-07 4.99999997 6.34443585e-07 4.99999997 6.34543585e-07 4.99999997 6.34643585e-07 4.99999997 6.34743585e-07 4.99999997 6.34843585e-07 4.99999997 6.34943585e-07 4.99999997 6.35043585e-07 4.99999997
+ 6.35143585e-07 4.99999997 6.35243585e-07 4.99999997 6.35343585e-07 4.99999997 6.35443585e-07 4.99999997 6.35543585e-07 4.99999997 6.35643585e-07 4.99999997 6.35743585e-07 4.99999997 6.35843585e-07 4.99999997
+ 6.35943585e-07 4.99999997 6.36043585e-07 4.99999997 6.36143585e-07 4.99999997 6.36243585e-07 4.99999997 6.36343585e-07 4.99999997 6.36443585e-07 4.99999997 6.36543585e-07 4.99999997 6.36643585e-07 4.99999997
+ 6.36743585e-07 4.99999997 6.36843585e-07 4.99999997 6.36943585e-07 4.99999997 6.37043585e-07 4.99999997 6.37143585e-07 4.99999997 6.37243585e-07 4.99999997 6.37343585e-07 4.99999997 6.37443585e-07 4.99999997
+ 6.37543585e-07 4.99999997 6.37643585e-07 4.99999997 6.37743585e-07 4.99999997 6.37843585e-07 4.99999997 6.37943585e-07 4.99999997 6.38043585e-07 4.99999997 6.38143585e-07 4.99999997 6.38243585e-07 4.99999997
+ 6.38343585e-07 4.99999997 6.38443585e-07 4.99999997 6.38543585e-07 4.99999997 6.38643585e-07 4.99999997 6.38743585e-07 4.99999997 6.38843585e-07 4.99999997 6.38943585e-07 4.99999997 6.39043585e-07 4.99999997
+ 6.39143585e-07 4.99999997 6.39243585e-07 4.99999997 6.39343585e-07 4.99999997 6.39443585e-07 4.99999997 6.39543585e-07 4.99999997 6.39643585e-07 4.99999997 6.39743585e-07 4.99999997 6.39843585e-07 4.99999997
+ 6.39943585e-07 4.99999997 6.40043585e-07 4.99999997 6.40143585e-07 4.99999997 6.40243585e-07 4.99999997 6.40343585e-07 4.99999997 6.40443585e-07 4.99999997 6.40543585e-07 4.99999997 6.40643585e-07 4.99999997
+ 6.40743585e-07 4.99999997 6.40843585e-07 4.99999997 6.40943585e-07 4.99999997 6.41043585e-07 4.99999997 6.41143585e-07 4.99999997 6.41243585e-07 4.99999997 6.41343585e-07 4.99999997 6.41443585e-07 4.99999997
+ 6.41543585e-07 4.99999997 6.41643585e-07 4.99999997 6.41743585e-07 4.99999997 6.41843585e-07 4.99999997 6.41943585e-07 4.99999997 6.42043585e-07 4.99999997 6.42143585e-07 4.99999997 6.42243585e-07 4.99999997
+ 6.42343585e-07 4.99999997 6.42443585e-07 4.99999997 6.42543585e-07 4.99999997 6.42643585e-07 4.99999997 6.42743585e-07 4.99999997 6.42843585e-07 4.99999997 6.42943585e-07 4.99999997 6.43043585e-07 4.99999997
+ 6.43143585e-07 4.99999997 6.43243585e-07 4.99999997 6.43343585e-07 4.99999997 6.43443585e-07 4.99999997 6.43543585e-07 4.99999997 6.43643585e-07 4.99999997 6.43743585e-07 4.99999997 6.43843585e-07 4.99999997
+ 6.43943585e-07 4.99999997 6.44043585e-07 4.99999997 6.44143585e-07 4.99999997 6.44243585e-07 4.99999997 6.44343585e-07 4.99999997 6.44443585e-07 4.99999997 6.44543585e-07 4.99999997 6.44643585e-07 4.99999997
+ 6.44743585e-07 4.99999997 6.44843585e-07 4.99999997 6.44943585e-07 4.99999997 6.45043585e-07 4.99999997 6.45143585e-07 4.99999997 6.45243585e-07 4.99999997 6.45343585e-07 4.99999997 6.45443585e-07 4.99999997
+ 6.45543585e-07 4.99999997 6.45643585e-07 4.99999997 6.45743585e-07 4.99999997 6.45843585e-07 4.99999997 6.45943585e-07 4.99999997 6.46043585e-07 4.99999997 6.46143585e-07 4.99999997 6.46243585e-07 4.99999997
+ 6.46343585e-07 4.99999997 6.46443585e-07 4.99999997 6.46543585e-07 4.99999997 6.46643585e-07 4.99999997 6.46743585e-07 4.99999997 6.46843585e-07 4.99999997 6.46943585e-07 4.99999997 6.47043585e-07 4.99999997
+ 6.47143585e-07 4.99999997 6.47243585e-07 4.99999997 6.47343585e-07 4.99999997 6.47443585e-07 4.99999997 6.47543585e-07 4.99999997 6.47643585e-07 4.99999997 6.47743585e-07 4.99999997 6.47843585e-07 4.99999997
+ 6.47943585e-07 4.99999997 6.48043585e-07 4.99999997 6.48143585e-07 4.99999997 6.48243585e-07 4.99999997 6.48343585e-07 4.99999997 6.48443585e-07 4.99999997 6.48543585e-07 4.99999997 6.48643585e-07 4.99999997
+ 6.48743585e-07 4.99999997 6.48843585e-07 4.99999997 6.48943585e-07 4.99999997 6.49043585e-07 4.99999997 6.49143585e-07 4.99999997 6.49243585e-07 4.99999997 6.49343585e-07 4.99999997 6.49443585e-07 4.99999997
+ 6.49543585e-07 4.99999997 6.49643585e-07 4.99999997 6.49743585e-07 4.99999997 6.49843585e-07 4.99999997 6.49943585e-07 4.99999997 6.50043585e-07 4.99999997 6.50143585e-07 4.99999997 6.50243585e-07 4.99999997
+ 6.50343585e-07 4.99999997 6.50443585e-07 4.99999997 6.50543585e-07 4.99999997 6.50643585e-07 4.99999997 6.50743585e-07 4.99999997 6.50843585e-07 4.99999997 6.50943585e-07 4.99999997 6.51e-07 4.99999997
+ 6.5101e-07 4.99999997 6.5103e-07 4.99999997 6.5107e-07 4.99999997 6.5115e-07 4.99999997 6.5125e-07 4.99999997 6.5135e-07 4.99999997 6.5145e-07 4.99999997 6.5155e-07 4.99999997
+ 6.5165e-07 4.99999997 6.5175e-07 4.99999997 6.5185e-07 4.99999997 6.51930828e-07 5.00000127 6.52e-07 5.00000077 6.52008608e-07 4.99998869 6.52025825e-07 4.99996401 6.52060258e-07 5.00000369
+ 6.52106181e-07 5.00005267 6.52150081e-07 4.99998208 6.52198026e-07 4.9999678 6.5225538e-07 5.00001892 6.52312019e-07 4.99999862 6.52404231e-07 5.00000003 6.52504231e-07 5.00000076 6.52604231e-07 4.99999856
+ 6.52704231e-07 5.00000151 6.52804231e-07 4.99999846 6.52904231e-07 5.00000136 6.53004231e-07 4.99999873 6.53104231e-07 5.00000105 6.53204231e-07 4.99999904 6.53304231e-07 5.00000077 6.53404231e-07 4.99999929
+ 6.53504231e-07 5.00000056 6.53604231e-07 4.99999946 6.53704231e-07 5.00000041 6.53804231e-07 4.99999959 6.53904231e-07 5.00000031 6.54004231e-07 4.99999967 6.54104231e-07 5.00000024 6.54204231e-07 4.99999973
+ 6.54304231e-07 5.00000019 6.54404231e-07 4.99999977 6.54504231e-07 5.00000015 6.54604231e-07 4.99999981 6.54704231e-07 5.00000013 6.54804231e-07 4.99999983 6.54904231e-07 5.0000001 6.55004231e-07 4.99999985
+ 6.55104231e-07 5.00000009 6.55204231e-07 4.99999987 6.55304231e-07 5.00000007 6.55404231e-07 4.99999988 6.55504231e-07 5.00000006 6.55604231e-07 4.99999989 6.55704231e-07 5.00000005 6.55804231e-07 4.9999999
+ 6.55904231e-07 5.00000004 6.56004231e-07 4.99999991 6.56104231e-07 5.00000003 6.56204231e-07 4.99999992 6.56304231e-07 5.00000003 6.56404231e-07 4.99999992 6.56504231e-07 5.00000002 6.56604231e-07 4.99999993
+ 6.56704231e-07 5.00000001 6.56804231e-07 4.99999993 6.56904231e-07 5.00000001 6.57004231e-07 4.99999994 6.57104231e-07 5.0 6.57204231e-07 4.99999994 6.57304231e-07 5.0 6.57404231e-07 4.99999994
+ 6.57504231e-07 5.0 6.57604231e-07 4.99999995 6.57704231e-07 4.99999999 6.57804231e-07 4.99999995 6.57904231e-07 4.99999999 6.58004231e-07 4.99999995 6.58104231e-07 4.99999999 6.58204231e-07 4.99999996
+ 6.58304231e-07 4.99999999 6.58404231e-07 4.99999996 6.58504231e-07 4.99999999 6.58604231e-07 4.99999996 6.58704231e-07 4.99999998 6.58804231e-07 4.99999996 6.58904231e-07 4.99999998 6.59004231e-07 4.99999996
+ 6.59104231e-07 4.99999998 6.59204231e-07 4.99999996 6.59304231e-07 4.99999998 6.59404231e-07 4.99999996 6.59504231e-07 4.99999998 6.59604231e-07 4.99999996 6.59704231e-07 4.99999998 6.59804231e-07 4.99999997
+ 6.59904231e-07 4.99999998 6.60004231e-07 4.99999997 6.60104231e-07 4.99999998 6.60204231e-07 4.99999997 6.60304231e-07 4.99999998 6.60404231e-07 4.99999997 6.60504231e-07 4.99999998 6.60604231e-07 4.99999997
+ 6.60704231e-07 4.99999998 6.60804231e-07 4.99999997 6.60904231e-07 4.99999998 6.61004231e-07 4.99999997 6.61104231e-07 4.99999998 6.61204231e-07 4.99999997 6.61304231e-07 4.99999997 6.61404231e-07 4.99999997
+ 6.61504231e-07 4.99999997 6.61604231e-07 4.99999997 6.61704231e-07 4.99999997 6.61804231e-07 4.99999997 6.61904231e-07 4.99999997 6.62004231e-07 4.99999997 6.62104231e-07 4.99999997 6.62204231e-07 4.99999997
+ 6.62304231e-07 4.99999997 6.62404231e-07 4.99999997 6.62504231e-07 4.99999997 6.62604231e-07 4.99999997 6.62704231e-07 4.99999997 6.62804231e-07 4.99999997 6.62904231e-07 4.99999997 6.63004231e-07 4.99999997
+ 6.63104231e-07 4.99999997 6.63204231e-07 4.99999997 6.63304231e-07 4.99999997 6.63404231e-07 4.99999997 6.63504231e-07 4.99999997 6.63604231e-07 4.99999997 6.63704231e-07 4.99999997 6.63804231e-07 4.99999997
+ 6.63904231e-07 4.99999997 6.64004231e-07 4.99999997 6.64104231e-07 4.99999997 6.64204231e-07 4.99999997 6.64304231e-07 4.99999997 6.64404231e-07 4.99999997 6.64504231e-07 4.99999997 6.64604231e-07 4.99999997
+ 6.64704231e-07 4.99999997 6.64804231e-07 4.99999997 6.64904231e-07 4.99999997 6.65004231e-07 4.99999997 6.65104231e-07 4.99999997 6.65204231e-07 4.99999997 6.65304231e-07 4.99999997 6.65404231e-07 4.99999997
+ 6.65504231e-07 4.99999997 6.65604231e-07 4.99999997 6.65704231e-07 4.99999997 6.65804231e-07 4.99999997 6.65904231e-07 4.99999997 6.66004231e-07 4.99999997 6.66104231e-07 4.99999997 6.66204231e-07 4.99999997
+ 6.66304231e-07 4.99999997 6.66404231e-07 4.99999997 6.66504231e-07 4.99999997 6.66604231e-07 4.99999997 6.66704231e-07 4.99999997 6.66804231e-07 4.99999997 6.66904231e-07 4.99999997 6.67004231e-07 4.99999997
+ 6.67104231e-07 4.99999997 6.67204231e-07 4.99999997 6.67304231e-07 4.99999997 6.67404231e-07 4.99999997 6.67504231e-07 4.99999997 6.67604231e-07 4.99999997 6.67704231e-07 4.99999997 6.67804231e-07 4.99999997
+ 6.67904231e-07 4.99999997 6.68004231e-07 4.99999997 6.68104231e-07 4.99999997 6.68204231e-07 4.99999997 6.68304231e-07 4.99999997 6.68404231e-07 4.99999997 6.68504231e-07 4.99999997 6.68604231e-07 4.99999997
+ 6.68704231e-07 4.99999997 6.68804231e-07 4.99999997 6.68904231e-07 4.99999997 6.69004231e-07 4.99999997 6.69104231e-07 4.99999997 6.69204231e-07 4.99999997 6.69304231e-07 4.99999997 6.69404231e-07 4.99999997
+ 6.69504231e-07 4.99999997 6.69604231e-07 4.99999997 6.69704231e-07 4.99999997 6.69804231e-07 4.99999997 6.69904231e-07 4.99999997 6.70004231e-07 4.99999997 6.70104231e-07 4.99999997 6.70204231e-07 4.99999997
+ 6.70304231e-07 4.99999997 6.70404231e-07 4.99999997 6.70504231e-07 4.99999997 6.70604231e-07 4.99999997 6.70704231e-07 4.99999997 6.70804231e-07 4.99999997 6.70904231e-07 4.99999997 6.71004231e-07 4.99999997
+ 6.71104231e-07 4.99999997 6.71204231e-07 4.99999997 6.71304231e-07 4.99999997 6.71404231e-07 4.99999997 6.71504231e-07 4.99999997 6.71604231e-07 4.99999997 6.71704231e-07 4.99999997 6.71804231e-07 4.99999997
+ 6.71904231e-07 4.99999997 6.72004231e-07 4.99999997 6.72104231e-07 4.99999997 6.72204231e-07 4.99999997 6.72304231e-07 4.99999997 6.72404231e-07 4.99999997 6.72504231e-07 4.99999997 6.72604231e-07 4.99999997
+ 6.72704231e-07 4.99999997 6.72804231e-07 4.99999997 6.72904231e-07 4.99999997 6.73004231e-07 4.99999997 6.73104231e-07 4.99999997 6.73204231e-07 4.99999997 6.73304231e-07 4.99999997 6.73404231e-07 4.99999997
+ 6.73504231e-07 4.99999997 6.73604231e-07 4.99999997 6.73704231e-07 4.99999997 6.73804231e-07 4.99999997 6.73904231e-07 4.99999997 6.74004231e-07 4.99999997 6.74104231e-07 4.99999997 6.74204231e-07 4.99999997
+ 6.74304231e-07 4.99999997 6.74404231e-07 4.99999997 6.74504231e-07 4.99999997 6.74604231e-07 4.99999997 6.74704231e-07 4.99999997 6.74804231e-07 4.99999997 6.74904231e-07 4.99999997 6.75004231e-07 4.99999997
+ 6.75104231e-07 4.99999997 6.75204231e-07 4.99999997 6.75304231e-07 4.99999997 6.75404231e-07 4.99999997 6.75504231e-07 4.99999997 6.75604231e-07 4.99999997 6.75704231e-07 4.99999997 6.75804231e-07 4.99999997
+ 6.75904231e-07 4.99999997 6.76004231e-07 4.99999997 6.76104231e-07 4.99999997 6.76204231e-07 4.99999997 6.76304231e-07 4.99999997 6.76404231e-07 4.99999997 6.76504231e-07 4.99999997 6.76604231e-07 4.99999997
+ 6.76704231e-07 4.99999997 6.76804231e-07 4.99999997 6.76904231e-07 4.99999997 6.77004231e-07 4.99999997 6.77104231e-07 4.99999997 6.77204231e-07 4.99999997 6.77304231e-07 4.99999997 6.77404231e-07 4.99999997
+ 6.77504231e-07 4.99999997 6.77604231e-07 4.99999997 6.77704231e-07 4.99999997 6.77804231e-07 4.99999997 6.77904231e-07 4.99999997 6.78004231e-07 4.99999997 6.78104231e-07 4.99999997 6.78204231e-07 4.99999997
+ 6.78304231e-07 4.99999997 6.78404231e-07 4.99999997 6.78504231e-07 4.99999997 6.78604231e-07 4.99999997 6.78704231e-07 4.99999997 6.78804231e-07 4.99999997 6.78904231e-07 4.99999997 6.79004231e-07 4.99999997
+ 6.79104231e-07 4.99999997 6.79204231e-07 4.99999997 6.79304231e-07 4.99999997 6.79404231e-07 4.99999997 6.79504231e-07 4.99999997 6.79604231e-07 4.99999997 6.79704231e-07 4.99999997 6.79804231e-07 4.99999997
+ 6.79904231e-07 4.99999997 6.80004231e-07 4.99999997 6.80104231e-07 4.99999997 6.80204231e-07 4.99999997 6.80304231e-07 4.99999997 6.80404231e-07 4.99999997 6.80504231e-07 4.99999997 6.80604231e-07 4.99999997
+ 6.80704231e-07 4.99999997 6.80804231e-07 4.99999997 6.80904231e-07 4.99999997 6.81004231e-07 4.99999997 6.81104231e-07 4.99999997 6.81204231e-07 4.99999997 6.81304231e-07 4.99999997 6.81404231e-07 4.99999997
+ 6.81504231e-07 4.99999997 6.81604231e-07 4.99999997 6.81704231e-07 4.99999997 6.81804231e-07 4.99999997 6.81904231e-07 4.99999997 6.82004231e-07 4.99999997 6.82104231e-07 4.99999997 6.82204231e-07 4.99999997
+ 6.82304231e-07 4.99999997 6.82404231e-07 4.99999997 6.82504231e-07 4.99999997 6.82604231e-07 4.99999997 6.82704231e-07 4.99999997 6.82804231e-07 4.99999997 6.82904231e-07 4.99999997 6.83004231e-07 4.99999997
+ 6.83104231e-07 4.99999997 6.83204231e-07 4.99999997 6.83304231e-07 4.99999997 6.83404231e-07 4.99999997 6.83504231e-07 4.99999997 6.83604231e-07 4.99999997 6.83704231e-07 4.99999997 6.83804231e-07 4.99999997
+ 6.83904231e-07 4.99999997 6.84004231e-07 4.99999997 6.84104231e-07 4.99999997 6.84204231e-07 4.99999997 6.84304231e-07 4.99999997 6.84404231e-07 4.99999997 6.84504231e-07 4.99999997 6.84604231e-07 4.99999997
+ 6.84704231e-07 4.99999997 6.84804231e-07 4.99999997 6.84904231e-07 4.99999997 6.85004231e-07 4.99999997 6.85104231e-07 4.99999997 6.85204231e-07 4.99999997 6.85304231e-07 4.99999997 6.85404231e-07 4.99999997
+ 6.85504231e-07 4.99999997 6.85604231e-07 4.99999997 6.85704231e-07 4.99999997 6.85804231e-07 4.99999997 6.85904231e-07 4.99999997 6.86004231e-07 4.99999997 6.86104231e-07 4.99999997 6.86204231e-07 4.99999997
+ 6.86304231e-07 4.99999997 6.86404231e-07 4.99999997 6.86504231e-07 4.99999997 6.86604231e-07 4.99999997 6.86704231e-07 4.99999997 6.86804231e-07 4.99999997 6.86904231e-07 4.99999997 6.87004231e-07 4.99999997
+ 6.87104231e-07 4.99999997 6.87204231e-07 4.99999997 6.87304231e-07 4.99999997 6.87404231e-07 4.99999997 6.87504231e-07 4.99999997 6.87604231e-07 4.99999997 6.87704231e-07 4.99999997 6.87804231e-07 4.99999997
+ 6.87904231e-07 4.99999997 6.88004231e-07 4.99999997 6.88104231e-07 4.99999997 6.88204231e-07 4.99999997 6.88304231e-07 4.99999997 6.88404231e-07 4.99999997 6.88504231e-07 4.99999997 6.88604231e-07 4.99999997
+ 6.88704231e-07 4.99999997 6.88804231e-07 4.99999997 6.88904231e-07 4.99999997 6.89004231e-07 4.99999997 6.89104231e-07 4.99999997 6.89204231e-07 4.99999997 6.89304231e-07 4.99999997 6.89404231e-07 4.99999997
+ 6.89504231e-07 4.99999997 6.89604231e-07 4.99999997 6.89704231e-07 4.99999997 6.89804231e-07 4.99999997 6.89904231e-07 4.99999997 6.90004231e-07 4.99999997 6.90104231e-07 4.99999997 6.90204231e-07 4.99999997
+ 6.90304231e-07 4.99999997 6.90404231e-07 4.99999997 6.90504231e-07 4.99999997 6.90604231e-07 4.99999997 6.90704231e-07 4.99999997 6.90804231e-07 4.99999997 6.90904231e-07 4.99999997 6.91004231e-07 4.99999997
+ 6.91104231e-07 4.99999997 6.91204231e-07 4.99999997 6.91304231e-07 4.99999997 6.91404231e-07 4.99999997 6.91504231e-07 4.99999997 6.91604231e-07 4.99999997 6.91704231e-07 4.99999997 6.91804231e-07 4.99999997
+ 6.91904231e-07 4.99999997 6.92004231e-07 4.99999997 6.92104231e-07 4.99999997 6.92204231e-07 4.99999997 6.92304231e-07 4.99999997 6.92404231e-07 4.99999997 6.92504231e-07 4.99999997 6.92604231e-07 4.99999997
+ 6.92704231e-07 4.99999997 6.92804231e-07 4.99999997 6.92904231e-07 4.99999997 6.93004231e-07 4.99999997 6.93104231e-07 4.99999997 6.93204231e-07 4.99999997 6.93304231e-07 4.99999997 6.93404231e-07 4.99999997
+ 6.93504231e-07 4.99999997 6.93604231e-07 4.99999997 6.93704231e-07 4.99999997 6.93804231e-07 4.99999997 6.93904231e-07 4.99999997 6.94004231e-07 4.99999997 6.94104231e-07 4.99999997 6.94204231e-07 4.99999997
+ 6.94304231e-07 4.99999997 6.94404231e-07 4.99999997 6.94504231e-07 4.99999997 6.94604231e-07 4.99999997 6.94704231e-07 4.99999997 6.94804231e-07 4.99999997 6.94904231e-07 4.99999997 6.95004231e-07 4.99999997
+ 6.95104231e-07 4.99999997 6.95204231e-07 4.99999997 6.95304231e-07 4.99999997 6.95404231e-07 4.99999997 6.95504231e-07 4.99999997 6.95604231e-07 4.99999997 6.95704231e-07 4.99999997 6.95804231e-07 4.99999997
+ 6.95904231e-07 4.99999997 6.96004231e-07 4.99999997 6.96104231e-07 4.99999997 6.96204231e-07 4.99999997 6.96304231e-07 4.99999997 6.96404231e-07 4.99999997 6.96504231e-07 4.99999997 6.96604231e-07 4.99999997
+ 6.96704231e-07 4.99999997 6.96804231e-07 4.99999997 6.96904231e-07 4.99999997 6.97004231e-07 4.99999997 6.97104231e-07 4.99999997 6.97204231e-07 4.99999997 6.97304231e-07 4.99999997 6.97404231e-07 4.99999997
+ 6.97504231e-07 4.99999997 6.97604231e-07 4.99999997 6.97704231e-07 4.99999997 6.97804231e-07 4.99999997 6.97904231e-07 4.99999997 6.98004231e-07 4.99999997 6.98104231e-07 4.99999997 6.98204231e-07 4.99999997
+ 6.98304231e-07 4.99999997 6.98404231e-07 4.99999997 6.98504231e-07 4.99999997 6.98604231e-07 4.99999997 6.98704231e-07 4.99999997 6.98804231e-07 4.99999997 6.98904231e-07 4.99999997 6.99004231e-07 4.99999997
+ 6.99104231e-07 4.99999997 6.99204231e-07 4.99999997 6.99304231e-07 4.99999997 6.99404231e-07 4.99999997 6.99504231e-07 4.99999997 6.99604231e-07 4.99999997 6.99704231e-07 4.99999997 6.99804231e-07 4.99999997
+ 6.99904231e-07 4.99999997 7e-07 4.99999997 7.0001e-07 4.99999997 7.0003e-07 4.99999997 7.0007e-07 4.99999997 7.0015e-07 4.99999997 7.0025e-07 4.99999997 7.0035e-07 4.99999997
+ 7.0045e-07 4.99999997 7.0055e-07 4.99999997 7.0065e-07 4.99999997 7.0075e-07 5.00000001 7.0085e-07 4.99999814 7.00931988e-07 5.00001158 7.01e-07 4.99997651 7.01008484e-07 4.99997816
+ 7.01025451e-07 4.99999556 7.01059385e-07 5.00001851 7.01090588e-07 5.00001181 7.01143428e-07 5.00000049 7.011991e-07 5.00001369 7.012991e-07 4.99978337 7.013991e-07 5.00014046 7.014991e-07 5.00032641
+ 7.01578678e-07 4.99987228 7.01663998e-07 4.99960593 7.01763998e-07 5.00049059 7.01858547e-07 4.99953494 7.01958547e-07 5.000381 7.02058547e-07 4.99971267 7.02158547e-07 5.00020063 7.02258547e-07 4.99986803
+ 7.02358547e-07 5.00007856 7.02458547e-07 4.99995925 7.02558547e-07 5.00001358 7.02658547e-07 5.00000443 7.02758547e-07 4.99998371 7.02858547e-07 5.00002377 7.02958547e-07 4.99997188 7.03058547e-07 5.0000303
+ 7.03158547e-07 4.99996886 7.03258547e-07 5.00003095 7.03358547e-07 4.99996972 7.03458547e-07 5.00002911 7.03558547e-07 4.99997213 7.03658547e-07 5.00002639 7.03758547e-07 4.99997499 7.03858547e-07 5.0000235
+ 7.03958547e-07 4.99997783 7.04058547e-07 5.00002075 7.04158547e-07 4.99998047 7.04258547e-07 5.00001824 7.04358547e-07 4.99998284 7.04458547e-07 5.000016 7.04558547e-07 4.99998495 7.04658547e-07 5.00001403
+ 7.04758547e-07 4.99998681 7.04858547e-07 5.00001229 7.04958547e-07 4.99998843 7.05058547e-07 5.00001077 7.05158547e-07 4.99998986 7.05258547e-07 5.00000943 7.05358547e-07 4.99999111 7.05458547e-07 5.00000826
+ 7.05558547e-07 4.99999221 7.05658547e-07 5.00000724 7.05758547e-07 4.99999317 7.05858547e-07 5.00000634 7.05958547e-07 4.99999401 7.06058547e-07 5.00000555 7.06158547e-07 4.99999474 7.06258547e-07 5.00000486
+ 7.06358547e-07 4.99999539 7.06458547e-07 5.00000426 7.06558547e-07 4.99999595 7.06658547e-07 5.00000373 7.06758547e-07 4.99999645 7.06858547e-07 5.00000327 7.06958547e-07 4.99999688 7.07058547e-07 5.00000286
+ 7.07158547e-07 4.99999727 7.07258547e-07 5.00000251 7.07358547e-07 4.9999976 7.07458547e-07 5.00000219 7.07558547e-07 4.99999789 7.07658547e-07 5.00000192 7.07758547e-07 4.99999815 7.07858547e-07 5.00000168
+ 7.07958547e-07 4.99999837 7.08058547e-07 5.00000147 7.08158547e-07 4.99999857 7.08258547e-07 5.00000128 7.08358547e-07 4.99999874 7.08458547e-07 5.00000112 7.08558547e-07 4.99999889 7.08658547e-07 5.00000098
+ 7.08758547e-07 4.99999903 7.08858547e-07 5.00000086 7.08958547e-07 4.99999914 7.09058547e-07 5.00000075 7.09158547e-07 4.99999925 7.09258547e-07 5.00000065 7.09358547e-07 4.99999934 7.09458547e-07 5.00000057
+ 7.09558547e-07 4.99999941 7.09658547e-07 5.00000049 7.09758547e-07 4.99999948 7.09858547e-07 5.00000043 7.09958547e-07 4.99999954 7.10058547e-07 5.00000037 7.10158547e-07 4.9999996 7.10258547e-07 5.00000032
+ 7.10358547e-07 4.99999964 7.10458547e-07 5.00000028 7.10558547e-07 4.99999968 7.10658547e-07 5.00000024 7.10758547e-07 4.99999972 7.10858547e-07 5.00000021 7.10958547e-07 4.99999975 7.11058547e-07 5.00000018
+ 7.11158547e-07 4.99999977 7.11258547e-07 5.00000015 7.11358547e-07 4.9999998 7.11458547e-07 5.00000013 7.11558547e-07 4.99999982 7.11658547e-07 5.00000011 7.11758547e-07 4.99999984 7.11858547e-07 5.00000009
+ 7.11958547e-07 4.99999986 7.12058547e-07 5.00000008 7.12158547e-07 4.99999987 7.12258547e-07 5.00000006 7.12358547e-07 4.99999988 7.12458547e-07 5.00000005 7.12558547e-07 4.99999989 7.12658547e-07 5.00000004
+ 7.12758547e-07 4.9999999 7.12858547e-07 5.00000003 7.12958547e-07 4.99999991 7.13058547e-07 5.00000003 7.13158547e-07 4.99999992 7.13258547e-07 5.00000002 7.13358547e-07 4.99999993 7.13458547e-07 5.00000001
+ 7.13558547e-07 4.99999993 7.13658547e-07 5.00000001 7.13758547e-07 4.99999994 7.13858547e-07 5.0 7.13958547e-07 4.99999994 7.14058547e-07 5.0 7.14158547e-07 4.99999995 7.14258547e-07 5.0
+ 7.14358547e-07 4.99999995 7.14458547e-07 4.99999999 7.14558547e-07 4.99999995 7.14658547e-07 4.99999999 7.14758547e-07 4.99999995 7.14858547e-07 4.99999999 7.14958547e-07 4.99999996 7.15058547e-07 4.99999999
+ 7.15158547e-07 4.99999996 7.15258547e-07 4.99999998 7.15358547e-07 4.99999996 7.15458547e-07 4.99999998 7.15558547e-07 4.99999996 7.15658547e-07 4.99999998 7.15758547e-07 4.99999996 7.15858547e-07 4.99999998
+ 7.15958547e-07 4.99999996 7.16058547e-07 4.99999998 7.16158547e-07 4.99999997 7.16258547e-07 4.99999998 7.16358547e-07 4.99999997 7.16458547e-07 4.99999998 7.16558547e-07 4.99999997 7.16658547e-07 4.99999998
+ 7.16758547e-07 4.99999997 7.16858547e-07 4.99999998 7.16958547e-07 4.99999997 7.17058547e-07 4.99999998 7.17158547e-07 4.99999997 7.17258547e-07 4.99999998 7.17358547e-07 4.99999997 7.17458547e-07 4.99999998
+ 7.17558547e-07 4.99999997 7.17658547e-07 4.99999997 7.17758547e-07 4.99999997 7.17858547e-07 4.99999997 7.17958547e-07 4.99999997 7.18058547e-07 4.99999997 7.18158547e-07 4.99999997 7.18258547e-07 4.99999997
+ 7.18358547e-07 4.99999997 7.18458547e-07 4.99999997 7.18558547e-07 4.99999997 7.18658547e-07 4.99999997 7.18758547e-07 4.99999997 7.18858547e-07 4.99999997 7.18958547e-07 4.99999997 7.19058547e-07 4.99999997
+ 7.19158547e-07 4.99999997 7.19258547e-07 4.99999997 7.19358547e-07 4.99999997 7.19458547e-07 4.99999997 7.19558547e-07 4.99999997 7.19658547e-07 4.99999997 7.19758547e-07 4.99999997 7.19858547e-07 4.99999997
+ 7.19958547e-07 4.99999997 7.20058547e-07 4.99999997 7.20158547e-07 4.99999997 7.20258547e-07 4.99999997 7.20358547e-07 4.99999997 7.20458547e-07 4.99999997 7.20558547e-07 4.99999997 7.20658547e-07 4.99999997
+ 7.20758547e-07 4.99999997 7.20858547e-07 4.99999997 7.20958547e-07 4.99999997 7.21058547e-07 4.99999997 7.21158547e-07 4.99999997 7.21258547e-07 4.99999997 7.21358547e-07 4.99999997 7.21458547e-07 4.99999997
+ 7.21558547e-07 4.99999997 7.21658547e-07 4.99999997 7.21758547e-07 4.99999997 7.21858547e-07 4.99999997 7.21958547e-07 4.99999997 7.22058547e-07 4.99999997 7.22158547e-07 4.99999997 7.22258547e-07 4.99999997
+ 7.22358547e-07 4.99999997 7.22458547e-07 4.99999997 7.22558547e-07 4.99999997 7.22658547e-07 4.99999997 7.22758547e-07 4.99999997 7.22858547e-07 4.99999997 7.22958547e-07 4.99999997 7.23058547e-07 4.99999997
+ 7.23158547e-07 4.99999997 7.23258547e-07 4.99999997 7.23358547e-07 4.99999997 7.23458547e-07 4.99999997 7.23558547e-07 4.99999997 7.23658547e-07 4.99999997 7.23758547e-07 4.99999997 7.23858547e-07 4.99999997
+ 7.23958547e-07 4.99999997 7.24058547e-07 4.99999997 7.24158547e-07 4.99999997 7.24258547e-07 4.99999997 7.24358547e-07 4.99999997 7.24458547e-07 4.99999997 7.24558547e-07 4.99999997 7.24658547e-07 4.99999997
+ 7.24758547e-07 4.99999997 7.24858547e-07 4.99999997 7.24958547e-07 4.99999997 7.25058547e-07 4.99999997 7.25158547e-07 4.99999997 7.25258547e-07 4.99999997 7.25358547e-07 4.99999997 7.25458547e-07 4.99999997
+ 7.25558547e-07 4.99999997 7.25658547e-07 4.99999997 7.25758547e-07 4.99999997 7.25858547e-07 4.99999997 7.25958547e-07 4.99999997 7.26058547e-07 4.99999997 7.26158547e-07 4.99999997 7.26258547e-07 4.99999997
+ 7.26358547e-07 4.99999997 7.26458547e-07 4.99999997 7.26558547e-07 4.99999997 7.26658547e-07 4.99999997 7.26758547e-07 4.99999997 7.26858547e-07 4.99999997 7.26958547e-07 4.99999997 7.27058547e-07 4.99999997
+ 7.27158547e-07 4.99999997 7.27258547e-07 4.99999997 7.27358547e-07 4.99999997 7.27458547e-07 4.99999997 7.27558547e-07 4.99999997 7.27658547e-07 4.99999997 7.27758547e-07 4.99999997 7.27858547e-07 4.99999997
+ 7.27958547e-07 4.99999997 7.28058547e-07 4.99999997 7.28158547e-07 4.99999997 7.28258547e-07 4.99999997 7.28358547e-07 4.99999997 7.28458547e-07 4.99999997 7.28558547e-07 4.99999997 7.28658547e-07 4.99999997
+ 7.28758547e-07 4.99999997 7.28858547e-07 4.99999997 7.28958547e-07 4.99999997 7.29058547e-07 4.99999997 7.29158547e-07 4.99999997 7.29258547e-07 4.99999997 7.29358547e-07 4.99999997 7.29458547e-07 4.99999997
+ 7.29558547e-07 4.99999997 7.29658547e-07 4.99999997 7.29758547e-07 4.99999997 7.29858547e-07 4.99999997 7.29958547e-07 4.99999997 7.30058547e-07 4.99999997 7.30158547e-07 4.99999997 7.30258547e-07 4.99999997
+ 7.30358547e-07 4.99999997 7.30458547e-07 4.99999997 7.30558547e-07 4.99999997 7.30658547e-07 4.99999997 7.30758547e-07 4.99999997 7.30858547e-07 4.99999997 7.30958547e-07 4.99999997 7.31058547e-07 4.99999997
+ 7.31158547e-07 4.99999997 7.31258547e-07 4.99999997 7.31358547e-07 4.99999997 7.31458547e-07 4.99999997 7.31558547e-07 4.99999997 7.31658547e-07 4.99999997 7.31758547e-07 4.99999997 7.31858547e-07 4.99999997
+ 7.31958547e-07 4.99999997 7.32058547e-07 4.99999997 7.32158547e-07 4.99999997 7.32258547e-07 4.99999997 7.32358547e-07 4.99999997 7.32458547e-07 4.99999997 7.32558547e-07 4.99999997 7.32658547e-07 4.99999997
+ 7.32758547e-07 4.99999997 7.32858547e-07 4.99999997 7.32958547e-07 4.99999997 7.33058547e-07 4.99999997 7.33158547e-07 4.99999997 7.33258547e-07 4.99999997 7.33358547e-07 4.99999997 7.33458547e-07 4.99999997
+ 7.33558547e-07 4.99999997 7.33658547e-07 4.99999997 7.33758547e-07 4.99999997 7.33858547e-07 4.99999997 7.33958547e-07 4.99999997 7.34058547e-07 4.99999997 7.34158547e-07 4.99999997 7.34258547e-07 4.99999997
+ 7.34358547e-07 4.99999997 7.34458547e-07 4.99999997 7.34558547e-07 4.99999997 7.34658547e-07 4.99999997 7.34758547e-07 4.99999997 7.34858547e-07 4.99999997 7.34958547e-07 4.99999997 7.35058547e-07 4.99999997
+ 7.35158547e-07 4.99999997 7.35258547e-07 4.99999997 7.35358547e-07 4.99999997 7.35458547e-07 4.99999997 7.35558547e-07 4.99999997 7.35658547e-07 4.99999997 7.35758547e-07 4.99999997 7.35858547e-07 4.99999997
+ 7.35958547e-07 4.99999997 7.36058547e-07 4.99999997 7.36158547e-07 4.99999997 7.36258547e-07 4.99999997 7.36358547e-07 4.99999997 7.36458547e-07 4.99999997 7.36558547e-07 4.99999997 7.36658547e-07 4.99999997
+ 7.36758547e-07 4.99999997 7.36858547e-07 4.99999997 7.36958547e-07 4.99999997 7.37058547e-07 4.99999997 7.37158547e-07 4.99999997 7.37258547e-07 4.99999997 7.37358547e-07 4.99999997 7.37458547e-07 4.99999997
+ 7.37558547e-07 4.99999997 7.37658547e-07 4.99999997 7.37758547e-07 4.99999997 7.37858547e-07 4.99999997 7.37958547e-07 4.99999997 7.38058547e-07 4.99999997 7.38158547e-07 4.99999997 7.38258547e-07 4.99999997
+ 7.38358547e-07 4.99999997 7.38458547e-07 4.99999997 7.38558547e-07 4.99999997 7.38658547e-07 4.99999997 7.38758547e-07 4.99999997 7.38858547e-07 4.99999997 7.38958547e-07 4.99999997 7.39058547e-07 4.99999997
+ 7.39158547e-07 4.99999997 7.39258547e-07 4.99999997 7.39358547e-07 4.99999997 7.39458547e-07 4.99999997 7.39558547e-07 4.99999997 7.39658547e-07 4.99999997 7.39758547e-07 4.99999997 7.39858547e-07 4.99999997
+ 7.39958547e-07 4.99999997 7.40058547e-07 4.99999997 7.40158547e-07 4.99999997 7.40258547e-07 4.99999997 7.40358547e-07 4.99999997 7.40458547e-07 4.99999997 7.40558547e-07 4.99999997 7.40658547e-07 4.99999997
+ 7.40758547e-07 4.99999997 7.40858547e-07 4.99999997 7.40958547e-07 4.99999997 7.41058547e-07 4.99999997 7.41158547e-07 4.99999997 7.41258547e-07 4.99999997 7.41358547e-07 4.99999997 7.41458547e-07 4.99999997
+ 7.41558547e-07 4.99999997 7.41658547e-07 4.99999997 7.41758547e-07 4.99999997 7.41858547e-07 4.99999997 7.41958547e-07 4.99999997 7.42058547e-07 4.99999997 7.42158547e-07 4.99999997 7.42258547e-07 4.99999997
+ 7.42358547e-07 4.99999997 7.42458547e-07 4.99999997 7.42558547e-07 4.99999997 7.42658547e-07 4.99999997 7.42758547e-07 4.99999997 7.42858547e-07 4.99999997 7.42958547e-07 4.99999997 7.43058547e-07 4.99999997
+ 7.43158547e-07 4.99999997 7.43258547e-07 4.99999997 7.43358547e-07 4.99999997 7.43458547e-07 4.99999997 7.43558547e-07 4.99999997 7.43658547e-07 4.99999997 7.43758547e-07 4.99999997 7.43858547e-07 4.99999997
+ 7.43958547e-07 4.99999997 7.44058547e-07 4.99999997 7.44158547e-07 4.99999997 7.44258547e-07 4.99999997 7.44358547e-07 4.99999997 7.44458547e-07 4.99999997 7.44558547e-07 4.99999997 7.44658547e-07 4.99999997
+ 7.44758547e-07 4.99999997 7.44858547e-07 4.99999997 7.44958547e-07 4.99999997 7.45058547e-07 4.99999997 7.45158547e-07 4.99999997 7.45258547e-07 4.99999997 7.45358547e-07 4.99999997 7.45458547e-07 4.99999997
+ 7.45558547e-07 4.99999997 7.45658547e-07 4.99999997 7.45758547e-07 4.99999997 7.45858547e-07 4.99999997 7.45958547e-07 4.99999997 7.46058547e-07 4.99999997 7.46158547e-07 4.99999997 7.46258547e-07 4.99999997
+ 7.46358547e-07 4.99999997 7.46458547e-07 4.99999997 7.46558547e-07 4.99999997 7.46658547e-07 4.99999997 7.46758547e-07 4.99999997 7.46858547e-07 4.99999997 7.46958547e-07 4.99999997 7.47058547e-07 4.99999997
+ 7.47158547e-07 4.99999997 7.47258547e-07 4.99999997 7.47358547e-07 4.99999997 7.47458547e-07 4.99999997 7.47558547e-07 4.99999997 7.47658547e-07 4.99999997 7.47758547e-07 4.99999997 7.47858547e-07 4.99999997
+ 7.47958547e-07 4.99999997 7.48058547e-07 4.99999997 7.48158547e-07 4.99999997 7.48258547e-07 4.99999997 7.48358547e-07 4.99999997 7.48458547e-07 4.99999997 7.48558547e-07 4.99999997 7.48658547e-07 4.99999997
+ 7.48758547e-07 4.99999997 7.48858547e-07 4.99999997 7.48958547e-07 4.99999997 7.49058547e-07 4.99999997 7.49158547e-07 4.99999997 7.49258547e-07 4.99999997 7.49358547e-07 4.99999997 7.49458547e-07 4.99999997
+ 7.49558547e-07 4.99999997 7.49658547e-07 4.99999997 7.49758547e-07 4.99999997 7.49858547e-07 4.99999997 7.49958547e-07 4.99999997 7.50058547e-07 4.99999997 7.50158547e-07 4.99999997 7.50258547e-07 4.99999997
+ 7.50358547e-07 4.99999997 7.50458547e-07 4.99999997 7.50558547e-07 4.99999997 7.50658547e-07 4.99999997 7.50758547e-07 4.99999997 7.50858547e-07 4.99999997 7.50958547e-07 4.99999997 7.51e-07 4.99999997
+ 7.5101e-07 4.99999997 7.5103e-07 4.99999997 7.5107e-07 4.99999997 7.5115e-07 4.99999997 7.5125e-07 4.99999997 7.5135e-07 4.99999997 7.5145e-07 4.99999997 7.5155e-07 4.99999997
+ 7.5165e-07 4.99999997 7.5175e-07 4.99999997 7.5185e-07 4.99999997 7.51930828e-07 5.00000123 7.52e-07 5.00000148 7.52008608e-07 4.99998858 7.52025825e-07 4.99996426 7.52060258e-07 5.00000424
+ 7.52106188e-07 5.00004614 7.52150118e-07 4.99998884 7.5219811e-07 4.99996906 7.522555e-07 5.0000164 7.52312176e-07 4.99999727 7.52404431e-07 5.00000287 7.52490759e-07 4.99999775 7.52590759e-07 5.0000011
+ 7.52690759e-07 4.99999973 7.52790759e-07 4.99999956 7.52890759e-07 5.00000078 7.52990759e-07 4.99999897 7.53090759e-07 5.00000104 7.53190759e-07 4.99999892 7.53290759e-07 5.00000096 7.53390759e-07 4.99999906
+ 7.53490759e-07 5.00000079 7.53590759e-07 4.99999924 7.53690759e-07 5.00000062 7.53790759e-07 4.99999939 7.53890759e-07 5.00000049 7.53990759e-07 4.99999951 7.54090759e-07 5.00000038 7.54190759e-07 4.9999996
+ 7.54290759e-07 5.00000031 7.54390759e-07 4.99999966 7.54490759e-07 5.00000025 7.54590759e-07 4.99999971 7.54690759e-07 5.00000021 7.54790759e-07 4.99999975 7.54890759e-07 5.00000018 7.54990759e-07 4.99999978
+ 7.55090759e-07 5.00000015 7.55190759e-07 4.9999998 7.55290759e-07 5.00000013 7.55390759e-07 4.99999983 7.55490759e-07 5.00000011 7.55590759e-07 4.99999984 7.55690759e-07 5.00000009 7.55790759e-07 4.99999986
+ 7.55890759e-07 5.00000008 7.55990759e-07 4.99999987 7.56090759e-07 5.00000007 7.56190759e-07 4.99999988 7.56290759e-07 5.00000006 7.56390759e-07 4.99999989 7.56490759e-07 5.00000005 7.56590759e-07 4.9999999
+ 7.56690759e-07 5.00000004 7.56790759e-07 4.99999991 7.56890759e-07 5.00000003 7.56990759e-07 4.99999992 7.57090759e-07 5.00000002 7.57190759e-07 4.99999992 7.57290759e-07 5.00000001 7.57390759e-07 4.99999993
+ 7.57490759e-07 5.00000001 7.57590759e-07 4.99999994 7.57690759e-07 5.00000001 7.57790759e-07 4.99999994 7.57890759e-07 5.0 7.57990759e-07 4.99999994 7.58090759e-07 5.0 7.58190759e-07 4.99999995
+ 7.58290759e-07 4.99999999 7.58390759e-07 4.99999995 7.58490759e-07 4.99999999 7.58590759e-07 4.99999995 7.58690759e-07 4.99999999 7.58790759e-07 4.99999996 7.58890759e-07 4.99999999 7.58990759e-07 4.99999996
+ 7.59090759e-07 4.99999999 7.59190759e-07 4.99999996 7.59290759e-07 4.99999998 7.59390759e-07 4.99999996 7.59490759e-07 4.99999998 7.59590759e-07 4.99999996 7.59690759e-07 4.99999998 7.59790759e-07 4.99999996
+ 7.59890759e-07 4.99999998 7.59990759e-07 4.99999996 7.60090759e-07 4.99999998 7.60190759e-07 4.99999997 7.60290759e-07 4.99999998 7.60390759e-07 4.99999997 7.60490759e-07 4.99999998 7.60590759e-07 4.99999997
+ 7.60690759e-07 4.99999998 7.60790759e-07 4.99999997 7.60890759e-07 4.99999998 7.60990759e-07 4.99999997 7.61090759e-07 4.99999998 7.61190759e-07 4.99999997 7.61290759e-07 4.99999998 7.61390759e-07 4.99999997
+ 7.61490759e-07 4.99999997 7.61590759e-07 4.99999997 7.61690759e-07 4.99999997 7.61790759e-07 4.99999997 7.61890759e-07 4.99999997 7.61990759e-07 4.99999997 7.62090759e-07 4.99999997 7.62190759e-07 4.99999997
+ 7.62290759e-07 4.99999997 7.62390759e-07 4.99999997 7.62490759e-07 4.99999997 7.62590759e-07 4.99999997 7.62690759e-07 4.99999997 7.62790759e-07 4.99999997 7.62890759e-07 4.99999997 7.62990759e-07 4.99999997
+ 7.63090759e-07 4.99999997 7.63190759e-07 4.99999997 7.63290759e-07 4.99999997 7.63390759e-07 4.99999997 7.63490759e-07 4.99999997 7.63590759e-07 4.99999997 7.63690759e-07 4.99999997 7.63790759e-07 4.99999997
+ 7.63890759e-07 4.99999997 7.63990759e-07 4.99999997 7.64090759e-07 4.99999997 7.64190759e-07 4.99999997 7.64290759e-07 4.99999997 7.64390759e-07 4.99999997 7.64490759e-07 4.99999997 7.64590759e-07 4.99999997
+ 7.64690759e-07 4.99999997 7.64790759e-07 4.99999997 7.64890759e-07 4.99999997 7.64990759e-07 4.99999997 7.65090759e-07 4.99999997 7.65190759e-07 4.99999997 7.65290759e-07 4.99999997 7.65390759e-07 4.99999997
+ 7.65490759e-07 4.99999997 7.65590759e-07 4.99999997 7.65690759e-07 4.99999997 7.65790759e-07 4.99999997 7.65890759e-07 4.99999997 7.65990759e-07 4.99999997 7.66090759e-07 4.99999997 7.66190759e-07 4.99999997
+ 7.66290759e-07 4.99999997 7.66390759e-07 4.99999997 7.66490759e-07 4.99999997 7.66590759e-07 4.99999997 7.66690759e-07 4.99999997 7.66790759e-07 4.99999997 7.66890759e-07 4.99999997 7.66990759e-07 4.99999997
+ 7.67090759e-07 4.99999997 7.67190759e-07 4.99999997 7.67290759e-07 4.99999997 7.67390759e-07 4.99999997 7.67490759e-07 4.99999997 7.67590759e-07 4.99999997 7.67690759e-07 4.99999997 7.67790759e-07 4.99999997
+ 7.67890759e-07 4.99999997 7.67990759e-07 4.99999997 7.68090759e-07 4.99999997 7.68190759e-07 4.99999997 7.68290759e-07 4.99999997 7.68390759e-07 4.99999997 7.68490759e-07 4.99999997 7.68590759e-07 4.99999997
+ 7.68690759e-07 4.99999997 7.68790759e-07 4.99999997 7.68890759e-07 4.99999997 7.68990759e-07 4.99999997 7.69090759e-07 4.99999997 7.69190759e-07 4.99999997 7.69290759e-07 4.99999997 7.69390759e-07 4.99999997
+ 7.69490759e-07 4.99999997 7.69590759e-07 4.99999997 7.69690759e-07 4.99999997 7.69790759e-07 4.99999997 7.69890759e-07 4.99999997 7.69990759e-07 4.99999997 7.70090759e-07 4.99999997 7.70190759e-07 4.99999997
+ 7.70290759e-07 4.99999997 7.70390759e-07 4.99999997 7.70490759e-07 4.99999997 7.70590759e-07 4.99999997 7.70690759e-07 4.99999997 7.70790759e-07 4.99999997 7.70890759e-07 4.99999997 7.70990759e-07 4.99999997
+ 7.71090759e-07 4.99999997 7.71190759e-07 4.99999997 7.71290759e-07 4.99999997 7.71390759e-07 4.99999997 7.71490759e-07 4.99999997 7.71590759e-07 4.99999997 7.71690759e-07 4.99999997 7.71790759e-07 4.99999997
+ 7.71890759e-07 4.99999997 7.71990759e-07 4.99999997 7.72090759e-07 4.99999997 7.72190759e-07 4.99999997 7.72290759e-07 4.99999997 7.72390759e-07 4.99999997 7.72490759e-07 4.99999997 7.72590759e-07 4.99999997
+ 7.72690759e-07 4.99999997 7.72790759e-07 4.99999997 7.72890759e-07 4.99999997 7.72990759e-07 4.99999997 7.73090759e-07 4.99999997 7.73190759e-07 4.99999997 7.73290759e-07 4.99999997 7.73390759e-07 4.99999997
+ 7.73490759e-07 4.99999997 7.73590759e-07 4.99999997 7.73690759e-07 4.99999997 7.73790759e-07 4.99999997 7.73890759e-07 4.99999997 7.73990759e-07 4.99999997 7.74090759e-07 4.99999997 7.74190759e-07 4.99999997
+ 7.74290759e-07 4.99999997 7.74390759e-07 4.99999997 7.74490759e-07 4.99999997 7.74590759e-07 4.99999997 7.74690759e-07 4.99999997 7.74790759e-07 4.99999997 7.74890759e-07 4.99999997 7.74990759e-07 4.99999997
+ 7.75090759e-07 4.99999997 7.75190759e-07 4.99999997 7.75290759e-07 4.99999997 7.75390759e-07 4.99999997 7.75490759e-07 4.99999997 7.75590759e-07 4.99999997 7.75690759e-07 4.99999997 7.75790759e-07 4.99999997
+ 7.75890759e-07 4.99999997 7.75990759e-07 4.99999997 7.76090759e-07 4.99999997 7.76190759e-07 4.99999997 7.76290759e-07 4.99999997 7.76390759e-07 4.99999997 7.76490759e-07 4.99999997 7.76590759e-07 4.99999997
+ 7.76690759e-07 4.99999997 7.76790759e-07 4.99999997 7.76890759e-07 4.99999997 7.76990759e-07 4.99999997 7.77090759e-07 4.99999997 7.77190759e-07 4.99999997 7.77290759e-07 4.99999997 7.77390759e-07 4.99999997
+ 7.77490759e-07 4.99999997 7.77590759e-07 4.99999997 7.77690759e-07 4.99999997 7.77790759e-07 4.99999997 7.77890759e-07 4.99999997 7.77990759e-07 4.99999997 7.78090759e-07 4.99999997 7.78190759e-07 4.99999997
+ 7.78290759e-07 4.99999997 7.78390759e-07 4.99999997 7.78490759e-07 4.99999997 7.78590759e-07 4.99999997 7.78690759e-07 4.99999997 7.78790759e-07 4.99999997 7.78890759e-07 4.99999997 7.78990759e-07 4.99999997
+ 7.79090759e-07 4.99999997 7.79190759e-07 4.99999997 7.79290759e-07 4.99999997 7.79390759e-07 4.99999997 7.79490759e-07 4.99999997 7.79590759e-07 4.99999997 7.79690759e-07 4.99999997 7.79790759e-07 4.99999997
+ 7.79890759e-07 4.99999997 7.79990759e-07 4.99999997 7.80090759e-07 4.99999997 7.80190759e-07 4.99999997 7.80290759e-07 4.99999997 7.80390759e-07 4.99999997 7.80490759e-07 4.99999997 7.80590759e-07 4.99999997
+ 7.80690759e-07 4.99999997 7.80790759e-07 4.99999997 7.80890759e-07 4.99999997 7.80990759e-07 4.99999997 7.81090759e-07 4.99999997 7.81190759e-07 4.99999997 7.81290759e-07 4.99999997 7.81390759e-07 4.99999997
+ 7.81490759e-07 4.99999997 7.81590759e-07 4.99999997 7.81690759e-07 4.99999997 7.81790759e-07 4.99999997 7.81890759e-07 4.99999997 7.81990759e-07 4.99999997 7.82090759e-07 4.99999997 7.82190759e-07 4.99999997
+ 7.82290759e-07 4.99999997 7.82390759e-07 4.99999997 7.82490759e-07 4.99999997 7.82590759e-07 4.99999997 7.82690759e-07 4.99999997 7.82790759e-07 4.99999997 7.82890759e-07 4.99999997 7.82990759e-07 4.99999997
+ 7.83090759e-07 4.99999997 7.83190759e-07 4.99999997 7.83290759e-07 4.99999997 7.83390759e-07 4.99999997 7.83490759e-07 4.99999997 7.83590759e-07 4.99999997 7.83690759e-07 4.99999997 7.83790759e-07 4.99999997
+ 7.83890759e-07 4.99999997 7.83990759e-07 4.99999997 7.84090759e-07 4.99999997 7.84190759e-07 4.99999997 7.84290759e-07 4.99999997 7.84390759e-07 4.99999997 7.84490759e-07 4.99999997 7.84590759e-07 4.99999997
+ 7.84690759e-07 4.99999997 7.84790759e-07 4.99999997 7.84890759e-07 4.99999997 7.84990759e-07 4.99999997 7.85090759e-07 4.99999997 7.85190759e-07 4.99999997 7.85290759e-07 4.99999997 7.85390759e-07 4.99999997
+ 7.85490759e-07 4.99999997 7.85590759e-07 4.99999997 7.85690759e-07 4.99999997 7.85790759e-07 4.99999997 7.85890759e-07 4.99999997 7.85990759e-07 4.99999997 7.86090759e-07 4.99999997 7.86190759e-07 4.99999997
+ 7.86290759e-07 4.99999997 7.86390759e-07 4.99999997 7.86490759e-07 4.99999997 7.86590759e-07 4.99999997 7.86690759e-07 4.99999997 7.86790759e-07 4.99999997 7.86890759e-07 4.99999997 7.86990759e-07 4.99999997
+ 7.87090759e-07 4.99999997 7.87190759e-07 4.99999997 7.87290759e-07 4.99999997 7.87390759e-07 4.99999997 7.87490759e-07 4.99999997 7.87590759e-07 4.99999997 7.87690759e-07 4.99999997 7.87790759e-07 4.99999997
+ 7.87890759e-07 4.99999997 7.87990759e-07 4.99999997 7.88090759e-07 4.99999997 7.88190759e-07 4.99999997 7.88290759e-07 4.99999997 7.88390759e-07 4.99999997 7.88490759e-07 4.99999997 7.88590759e-07 4.99999997
+ 7.88690759e-07 4.99999997 7.88790759e-07 4.99999997 7.88890759e-07 4.99999997 7.88990759e-07 4.99999997 7.89090759e-07 4.99999997 7.89190759e-07 4.99999997 7.89290759e-07 4.99999997 7.89390759e-07 4.99999997
+ 7.89490759e-07 4.99999997 7.89590759e-07 4.99999997 7.89690759e-07 4.99999997 7.89790759e-07 4.99999997 7.89890759e-07 4.99999997 7.89990759e-07 4.99999997 7.90090759e-07 4.99999997 7.90190759e-07 4.99999997
+ 7.90290759e-07 4.99999997 7.90390759e-07 4.99999997 7.90490759e-07 4.99999997 7.90590759e-07 4.99999997 7.90690759e-07 4.99999997 7.90790759e-07 4.99999997 7.90890759e-07 4.99999997 7.90990759e-07 4.99999997
+ 7.91090759e-07 4.99999997 7.91190759e-07 4.99999997 7.91290759e-07 4.99999997 7.91390759e-07 4.99999997 7.91490759e-07 4.99999997 7.91590759e-07 4.99999997 7.91690759e-07 4.99999997 7.91790759e-07 4.99999997
+ 7.91890759e-07 4.99999997 7.91990759e-07 4.99999997 7.92090759e-07 4.99999997 7.92190759e-07 4.99999997 7.92290759e-07 4.99999997 7.92390759e-07 4.99999997 7.92490759e-07 4.99999997 7.92590759e-07 4.99999997
+ 7.92690759e-07 4.99999997 7.92790759e-07 4.99999997 7.92890759e-07 4.99999997 7.92990759e-07 4.99999997 7.93090759e-07 4.99999997 7.93190759e-07 4.99999997 7.93290759e-07 4.99999997 7.93390759e-07 4.99999997
+ 7.93490759e-07 4.99999997 7.93590759e-07 4.99999997 7.93690759e-07 4.99999997 7.93790759e-07 4.99999997 7.93890759e-07 4.99999997 7.93990759e-07 4.99999997 7.94090759e-07 4.99999997 7.94190759e-07 4.99999997
+ 7.94290759e-07 4.99999997 7.94390759e-07 4.99999997 7.94490759e-07 4.99999997 7.94590759e-07 4.99999997 7.94690759e-07 4.99999997 7.94790759e-07 4.99999997 7.94890759e-07 4.99999997 7.94990759e-07 4.99999997
+ 7.95090759e-07 4.99999997 7.95190759e-07 4.99999997 7.95290759e-07 4.99999997 7.95390759e-07 4.99999997 7.95490759e-07 4.99999997 7.95590759e-07 4.99999997 7.95690759e-07 4.99999997 7.95790759e-07 4.99999997
+ 7.95890759e-07 4.99999997 7.95990759e-07 4.99999997 7.96090759e-07 4.99999997 7.96190759e-07 4.99999997 7.96290759e-07 4.99999997 7.96390759e-07 4.99999997 7.96490759e-07 4.99999997 7.96590759e-07 4.99999997
+ 7.96690759e-07 4.99999997 7.96790759e-07 4.99999997 7.96890759e-07 4.99999997 7.96990759e-07 4.99999997 7.97090759e-07 4.99999997 7.97190759e-07 4.99999997 7.97290759e-07 4.99999997 7.97390759e-07 4.99999997
+ 7.97490759e-07 4.99999997 7.97590759e-07 4.99999997 7.97690759e-07 4.99999997 7.97790759e-07 4.99999997 7.97890759e-07 4.99999997 7.97990759e-07 4.99999997 7.98090759e-07 4.99999997 7.98190759e-07 4.99999997
+ 7.98290759e-07 4.99999997 7.98390759e-07 4.99999997 7.98490759e-07 4.99999997 7.98590759e-07 4.99999997 7.98690759e-07 4.99999997 7.98790759e-07 4.99999997 7.98890759e-07 4.99999997 7.98990759e-07 4.99999997
+ 7.99090759e-07 4.99999997 7.99190759e-07 4.99999997 7.99290759e-07 4.99999997 7.99390759e-07 4.99999997 7.99490759e-07 4.99999997 7.99590759e-07 4.99999997 7.99690759e-07 4.99999997 7.99790759e-07 4.99999997
+ 7.99890759e-07 4.99999997 7.99990759e-07 4.99999997 8e-07 4.99999997 8.0001e-07 4.99999997 8.0003e-07 4.99999997 8.0007e-07 4.99999997 8.0015e-07 4.99999997 8.0025e-07 4.99999997
+ 8.0035e-07 4.99999997 8.0045e-07 4.99999997 8.0055e-07 4.99999997 8.0065e-07 4.99999997 8.0075e-07 5.00000001 8.0085e-07 4.99999686 8.00931913e-07 5.00000385 8.01e-07 5.00010633
+ 8.01008477e-07 5.00014453 8.01025432e-07 5.00027393 8.01059342e-07 4.99937073 8.01090545e-07 4.99743534 8.01143412e-07 4.99875515 8.01199108e-07 5.05834962 8.01266691e-07 4.82390127 8.01329415e-07 1.08191107
+ 8.01394829e-07 -0.0834648083 8.01464618e-07 0.122803197 8.01533535e-07 -0.0865031891 8.01610366e-07 0.0799022498 8.01709241e-07 -0.071357353 8.01809241e-07 0.0656628381 8.01909241e-07 -0.0593137472 8.02009241e-07 0.0545273436
+ 8.02109241e-07 -0.0493042956 8.02209241e-07 0.0453245048 8.02309241e-07 -0.0410570554 8.02409241e-07 0.037700894 8.02509241e-07 -0.0342011994 8.02609241e-07 0.0313787965 8.02709241e-07 -0.0285001312 8.02809241e-07 0.0261309755
+ 8.02909241e-07 -0.0237572942 8.03009241e-07 0.0217710974 8.03109241e-07 -0.0198097687 8.03209241e-07 0.0181460851 8.03309241e-07 -0.0165226519 8.03409241e-07 0.0151299819 8.03509241e-07 -0.0137842547 8.03609241e-07 0.0126189805
+ 8.03709241e-07 -0.0115020691 8.03809241e-07 0.0105273918 8.03909241e-07 -0.00959941956 8.04009241e-07 0.00878437449 8.04109241e-07 -0.0080127004 8.04209241e-07 0.00733127901 8.04309241e-07 -0.00668910201 8.04409241e-07 0.00611948647
+ 8.04509241e-07 -0.00558474235 8.04609241e-07 0.00510864727 8.04709241e-07 -0.00466313017 8.04809241e-07 0.00426524119 8.04909241e-07 -0.00389389982 8.05009241e-07 0.00356139756 8.05109241e-07 -0.00325176812 8.05209241e-07 0.00297392599
+ 8.05309241e-07 -0.00271567297 8.05409241e-07 0.00248351831 8.05509241e-07 -0.00226806096 8.05609241e-07 0.00207409017 8.05709241e-07 -0.00189429747 8.05809241e-07 0.00173223667 8.05909241e-07 -0.00158217745 8.06009241e-07 0.00144678179
+ 8.06109241e-07 -0.00132151935 8.06209241e-07 0.00120840479 8.06309241e-07 -0.00110382775 8.06409241e-07 0.0010093302 8.06509241e-07 -0.000922012818 8.06609241e-07 0.000843070142 8.06709241e-07 -0.00077015679 8.06809241e-07 0.000704210127
+ 8.06909241e-07 -0.000641698121 8.07009241e-07 0.000588620508 8.07109241e-07 -0.000537460404 8.07209241e-07 0.00049143601 8.07309241e-07 -0.000448954494 8.07409241e-07 0.000410509151 8.07509241e-07 -0.00037502548 8.07609241e-07 0.000342912489
+ 8.07709241e-07 -0.000313272133 8.07809241e-07 0.000286449239 8.07909241e-07 -0.000260434291 8.08009241e-07 0.000239494613 8.08109241e-07 -0.000217572043 8.08209241e-07 0.000200138431 8.08309241e-07 -0.000181776513 8.08409241e-07 0.000168412028
+ 8.08509241e-07 -0.000151700166 8.08609241e-07 0.000140636669 8.08709241e-07 -0.000126668718 8.08809241e-07 0.000117445566 8.08909241e-07 -0.00010577273 8.09009241e-07 9.80823968e-05 8.09109241e-07 -8.83271665e-05 8.09209241e-07 8.19142604e-05
+ 8.09309241e-07 -7.37611653e-05 8.09409241e-07 6.84132514e-05 8.09509241e-07 -6.15986662e-05 8.09609241e-07 5.71389142e-05 8.09709241e-07 -5.14425502e-05 8.09809241e-07 4.77236794e-05 8.09909241e-07 -4.29614712e-05 8.10009241e-07 3.98607554e-05
+ 8.10109241e-07 -3.5878914e-05 8.10209241e-07 3.32940479e-05 8.10309241e-07 -2.99640861e-05 8.10409241e-07 2.78097581e-05 8.10509241e-07 -2.50243268e-05 8.10609241e-07 2.32293653e-05 8.10709241e-07 -2.08987797e-05 8.10809241e-07 1.94038161e-05
+ 8.10909241e-07 -1.7453167e-05 8.11009241e-07 1.62086675e-05 8.11109241e-07 -1.45753822e-05 8.11209241e-07 1.35400087e-05 8.11309241e-07 -1.21718182e-05 8.11409241e-07 1.13110661e-05 8.11509241e-07 -1.01643087e-05 8.11609241e-07 9.44937439e-06
+ 8.11709241e-07 -8.48757837e-06 8.11809241e-07 7.89441434e-06 8.11909241e-07 -7.08713851e-06 8.12009241e-07 6.59570205e-06 8.12109241e-07 -5.91746374e-06 8.12209241e-07 5.51092447e-06 8.12309241e-07 -4.94046151e-06 8.12409241e-07 4.60484172e-06
+ 8.12509241e-07 -4.12441064e-06 8.12609241e-07 3.84802635e-06 8.12709241e-07 -3.44279985e-06 8.12809241e-07 3.21589029e-06 8.12909241e-07 -2.8734813e-06 8.13009241e-07 2.68789385e-06 8.13109241e-07 -2.39795499e-06 8.13209241e-07 2.2468806e-06
+ 8.13309241e-07 -2.00076871e-06 8.13409241e-07 1.87852049e-06 8.13509241e-07 -1.66901602e-06 8.13609241e-07 1.57084431e-06 8.13709241e-07 -1.39191691e-06 8.13809241e-07 1.31385476e-06 8.13909241e-07 -1.16046737e-06 8.14009241e-07 1.09920149e-06
+ 8.14109241e-07 -9.67146834e-07 8.14209241e-07 9.19909936e-07 8.14309241e-07 -8.05673783e-07 8.14409241e-07 7.70154473e-07 8.14509241e-07 -6.7080149e-07 8.14609241e-07 6.45069407e-07 8.14709241e-07 -5.58147936e-07 8.14809241e-07 5.40590661e-07
+ 8.14909241e-07 -4.64052764e-07 8.15009241e-07 4.53323507e-07 8.15109241e-07 -3.8545863e-07 8.15209241e-07 3.80432504e-07 8.15309241e-07 -3.19811887e-07 8.15409241e-07 3.1954934e-07 8.15509241e-07 -2.64979597e-07 8.15609241e-07 2.68695866e-07
+ 8.15709241e-07 -2.19180201e-07 8.15809241e-07 2.26219815e-07 8.15909241e-07 -1.8092564e-07 8.16009241e-07 1.90741111e-07 8.16109241e-07 -1.48972995e-07 8.16209241e-07 1.6110703e-07 8.16309241e-07 -1.22284104e-07 8.16409241e-07 1.36354746e-07
+ 8.16509241e-07 -9.99918294e-08 8.16609241e-07 1.15680046e-07 8.16709241e-07 -8.13718872e-08 8.16809241e-07 9.84112048e-08 8.16909241e-07 -6.58223735e-08 8.17009241e-07 8.39929852e-08 8.17109241e-07 -5.284004e-08 8.17209241e-07 7.19556155e-08
+ 8.17309241e-07 -4.2001428e-08 8.17409241e-07 6.19059217e-08 8.17509241e-07 -3.29525416e-08 8.17609241e-07 5.35156812e-08 8.17709241e-07 -2.53978474e-08 8.17809241e-07 4.65108739e-08 8.17909241e-07 -1.90906164e-08 8.18009241e-07 4.06627303e-08
+ 8.18109241e-07 -1.38111839e-08 8.18209241e-07 3.57678313e-08 8.18309241e-07 -9.41798312e-09 8.18409241e-07 3.16941589e-08 8.18509241e-07 -5.74987449e-09 8.18609241e-07 2.82930291e-08 8.18709241e-07 -2.68736194e-09 8.18809241e-07 2.54534265e-08
+ 8.18909241e-07 -1.30473965e-10 8.19009241e-07 2.30826486e-08 8.19109241e-07 2.00426414e-09 8.19209241e-07 2.11293848e-08 8.19309241e-07 3.76433651e-09 8.19409241e-07 1.95203311e-08 8.19509241e-07 5.21432736e-09 8.19609241e-07 1.81947456e-08
+ 8.19709241e-07 6.40887901e-09 8.19809241e-07 1.71026802e-08 8.19909241e-07 7.39299602e-09 8.20009241e-07 1.62029947e-08 8.20109241e-07 8.2037514e-09 8.20209241e-07 1.53618154e-08 8.20309241e-07 8.85747617e-09 8.20409241e-07 1.4763059e-08
+ 8.20509241e-07 9.40108796e-09 8.20609241e-07 1.42694719e-08 8.20709241e-07 9.84925336e-09 8.20809241e-07 1.38625607e-08 8.20909241e-07 1.0218713e-08 8.21009241e-07 1.35271143e-08 8.21109241e-07 1.05232837e-08 8.21209241e-07 1.3250585e-08
+ 8.21309241e-07 1.07743599e-08 8.21409241e-07 1.30226259e-08 8.21509241e-07 1.09813364e-08 8.21609241e-07 1.28347068e-08 8.21709241e-07 1.11519594e-08 8.21809241e-07 1.26797948e-08 8.21909241e-07 1.12926135e-08 8.22009241e-07 1.25520923e-08
+ 8.22109241e-07 1.14085627e-08 8.22209241e-07 1.24468203e-08 8.22309241e-07 1.15041462e-08 8.22409241e-07 1.23600388e-08 8.22509241e-07 1.15829411e-08 8.22609241e-07 1.22885005e-08 8.22709241e-07 1.16478963e-08 8.22809241e-07 1.2229528e-08
+ 8.22909241e-07 1.17014426e-08 8.23009241e-07 1.21809137e-08 8.23109241e-07 1.17455837e-08 8.23209241e-07 1.21408381e-08 8.23309241e-07 1.17819722e-08 8.23409241e-07 1.2107802e-08 8.23509241e-07 1.18119693e-08 8.23609241e-07 1.2080569e-08
+ 8.23709241e-07 1.18366978e-08 8.23809241e-07 1.20581192e-08 8.23909241e-07 1.18570828e-08 8.24009241e-07 1.20396129e-08 8.24109241e-07 1.18738876e-08 8.24209241e-07 1.20243571e-08 8.24309241e-07 1.18877407e-08 8.24409241e-07 1.20117812e-08
+ 8.24509241e-07 1.18991606e-08 8.24609241e-07 1.20014143e-08 8.24709241e-07 1.1908575e-08 8.24809241e-07 1.19928685e-08 8.24909241e-07 1.19163359e-08 8.25009241e-07 1.19858236e-08 8.25109241e-07 1.19227341e-08 8.25209241e-07 1.19800164e-08
+ 8.25309241e-07 1.1928008e-08 8.25409241e-07 1.19752293e-08 8.25509241e-07 1.19323559e-08 8.25609241e-07 1.19712832e-08 8.25709241e-07 1.19359404e-08 8.25809241e-07 1.19680302e-08 8.25909241e-07 1.19388954e-08 8.26009241e-07 1.19653485e-08
+ 8.26109241e-07 1.19413315e-08 8.26209241e-07 1.19631381e-08 8.26309241e-07 1.19433398e-08 8.26409241e-07 1.19613162e-08 8.26509241e-07 1.19449956e-08 8.26609241e-07 1.19598141e-08 8.26709241e-07 1.19463605e-08 8.26809241e-07 1.19585763e-08
+ 8.26909241e-07 1.19474855e-08 8.27009241e-07 1.19575561e-08 8.27109241e-07 1.19484131e-08 8.27209241e-07 1.19567148e-08 8.27309241e-07 1.19491778e-08 8.27409241e-07 1.19560217e-08 8.27509241e-07 1.19498085e-08 8.27609241e-07 1.19554503e-08
+ 8.27709241e-07 1.19503282e-08 8.27809241e-07 1.19549795e-08 8.27909241e-07 1.19507569e-08 8.28009241e-07 1.19545911e-08 8.28109241e-07 1.19511105e-08 8.28209241e-07 1.19542709e-08 8.28309241e-07 1.19514016e-08 8.28409241e-07 1.19540074e-08
+ 8.28509241e-07 1.19516422e-08 8.28609241e-07 1.19537903e-08 8.28709241e-07 1.19518405e-08 8.28809241e-07 1.19536113e-08 8.28909241e-07 1.19520038e-08 8.29009241e-07 1.19534637e-08 8.29109241e-07 1.19521385e-08 8.29209241e-07 1.19533421e-08
+ 8.29309241e-07 1.19522498e-08 8.29409241e-07 1.19532421e-08 8.29509241e-07 1.19523414e-08 8.29609241e-07 1.19531597e-08 8.29709241e-07 1.19524171e-08 8.29809241e-07 1.19530916e-08 8.29909241e-07 1.19524796e-08 8.30009241e-07 1.19530356e-08
+ 8.30109241e-07 1.19525311e-08 8.30209241e-07 1.19529897e-08 8.30309241e-07 1.19525737e-08 8.30409241e-07 1.19529515e-08 8.30509241e-07 1.19526087e-08 8.30609241e-07 1.19529204e-08 8.30709241e-07 1.19526377e-08 8.30809241e-07 1.19528948e-08
+ 8.30909241e-07 1.19526615e-08 8.31009241e-07 1.19528738e-08 8.31109241e-07 1.19526815e-08 8.31209241e-07 1.19528562e-08 8.31309241e-07 1.19526979e-08 8.31409241e-07 1.19528421e-08 8.31509241e-07 1.19527115e-08 8.31609241e-07 1.19528304e-08
+ 8.31709241e-07 1.19527227e-08 8.31809241e-07 1.19528206e-08 8.31909241e-07 1.19527322e-08 8.32009241e-07 1.19528127e-08 8.32109241e-07 1.19527401e-08 8.32209241e-07 1.1952806e-08 8.32309241e-07 1.19527463e-08 8.32409241e-07 1.1952801e-08
+ 8.32509241e-07 1.19527518e-08 8.32609241e-07 1.19527966e-08 8.32709241e-07 1.19527563e-08 8.32809241e-07 1.19527932e-08 8.32909241e-07 1.19527596e-08 8.33009241e-07 1.19527904e-08 8.33109241e-07 1.19527629e-08 8.33209241e-07 1.1952788e-08
+ 8.33309241e-07 1.19527654e-08 8.33409241e-07 1.1952786e-08 8.33509241e-07 1.19527677e-08 8.33609241e-07 1.19527845e-08 8.33709241e-07 1.19527694e-08 8.33809241e-07 1.19527834e-08 8.33909241e-07 1.19527708e-08 8.34009241e-07 1.19527826e-08
+ 8.34109241e-07 1.19527722e-08 8.34209241e-07 1.19527817e-08 8.34309241e-07 1.19527729e-08 8.34409241e-07 1.19527811e-08 8.34509241e-07 1.19527741e-08 8.34609241e-07 1.19527807e-08 8.34709241e-07 1.19527749e-08 8.34809241e-07 1.19527804e-08
+ 8.34909241e-07 1.19527755e-08 8.35009241e-07 1.195278e-08 8.35109241e-07 1.19527762e-08 8.35209241e-07 1.19527801e-08 8.35309241e-07 1.19527767e-08 8.35409241e-07 1.19527799e-08 8.35509241e-07 1.19527771e-08 8.35609241e-07 1.19527799e-08
+ 8.35709241e-07 1.19527775e-08 8.35809241e-07 1.19527798e-08 8.35909241e-07 1.19527777e-08 8.36009241e-07 1.195278e-08 8.36109241e-07 1.1952778e-08 8.36209241e-07 1.195278e-08 8.36309241e-07 1.19527784e-08 8.36409241e-07 1.195278e-08
+ 8.36509241e-07 1.19527786e-08 8.36609241e-07 1.195278e-08 8.36709241e-07 1.19527789e-08 8.36809241e-07 1.19527799e-08 8.36909241e-07 1.19527795e-08 8.37009241e-07 1.19527802e-08 8.37109241e-07 1.19527794e-08 8.37209241e-07 1.19527799e-08
+ 8.37309241e-07 1.19527797e-08 8.37409241e-07 1.195278e-08 8.37509241e-07 1.19527802e-08 8.37609241e-07 1.19527804e-08 8.37709241e-07 1.19527803e-08 8.37809241e-07 1.19527802e-08 8.37909241e-07 1.19527804e-08 8.38009241e-07 1.19527807e-08
+ 8.38109241e-07 1.19527803e-08 8.38209241e-07 1.19527807e-08 8.38309241e-07 1.19527809e-08 8.38409241e-07 1.19527805e-08 8.38509241e-07 1.19527805e-08 8.38609241e-07 1.19527808e-08 8.38709241e-07 1.1952781e-08 8.38809241e-07 1.19527808e-08
+ 8.38909241e-07 1.19527809e-08 8.39009241e-07 1.19527808e-08 8.39109241e-07 1.19527813e-08 8.39209241e-07 1.19527812e-08 8.39309241e-07 1.19527815e-08 8.39409241e-07 1.19527815e-08 8.39509241e-07 1.19527814e-08 8.39609241e-07 1.19527815e-08
+ 8.39709241e-07 1.19527816e-08 8.39809241e-07 1.19527814e-08 8.39909241e-07 1.19527816e-08 8.40009241e-07 1.19527818e-08 8.40109241e-07 1.19527818e-08 8.40209241e-07 1.1952782e-08 8.40309241e-07 1.19527818e-08 8.40409241e-07 1.1952782e-08
+ 8.40509241e-07 1.19527819e-08 8.40609241e-07 1.19527821e-08 8.40709241e-07 1.19527822e-08 8.40809241e-07 1.19527823e-08 8.40909241e-07 1.19527819e-08 8.41009241e-07 1.19527821e-08 8.41109241e-07 1.19527823e-08 8.41209241e-07 1.1952782e-08
+ 8.41309241e-07 1.19527822e-08 8.41409241e-07 1.19527824e-08 8.41509241e-07 1.19527823e-08 8.41609241e-07 1.19527826e-08 8.41709241e-07 1.19527826e-08 8.41809241e-07 1.19527823e-08 8.41909241e-07 1.19527826e-08 8.42009241e-07 1.19527828e-08
+ 8.42109241e-07 1.19527826e-08 8.42209241e-07 1.19527825e-08 8.42309241e-07 1.19527829e-08 8.42409241e-07 1.19527826e-08 8.42509241e-07 1.19527827e-08 8.42609241e-07 1.19527831e-08 8.42709241e-07 1.19527826e-08 8.42809241e-07 1.19527828e-08
+ 8.42909241e-07 1.1952783e-08 8.43009241e-07 1.19527831e-08 8.43109241e-07 1.19527831e-08 8.43209241e-07 1.1952783e-08 8.43309241e-07 1.19527833e-08 8.43409241e-07 1.19527833e-08 8.43509241e-07 1.19527833e-08 8.43609241e-07 1.19527831e-08
+ 8.43709241e-07 1.19527832e-08 8.43809241e-07 1.19527835e-08 8.43909241e-07 1.19527833e-08 8.44009241e-07 1.19527835e-08 8.44109241e-07 1.19527834e-08 8.44209241e-07 1.19527837e-08 8.44309241e-07 1.19527835e-08 8.44409241e-07 1.19527836e-08
+ 8.44509241e-07 1.19527835e-08 8.44609241e-07 1.19527837e-08 8.44709241e-07 1.19527834e-08 8.44809241e-07 1.1952784e-08 8.44909241e-07 1.19527837e-08 8.45009241e-07 1.1952784e-08 8.45109241e-07 1.19527837e-08 8.45209241e-07 1.19527839e-08
+ 8.45309241e-07 1.19527836e-08 8.45409241e-07 1.19527838e-08 8.45509241e-07 1.19527838e-08 8.45609241e-07 1.19527843e-08 8.45709241e-07 1.1952784e-08 8.45809241e-07 1.1952784e-08 8.45909241e-07 1.19527841e-08 8.46009241e-07 1.19527844e-08
+ 8.46109241e-07 1.19527841e-08 8.46209241e-07 1.19527843e-08 8.46309241e-07 1.1952784e-08 8.46409241e-07 1.19527843e-08 8.46509241e-07 1.19527844e-08 8.46609241e-07 1.19527841e-08 8.46709241e-07 1.19527842e-08 8.46809241e-07 1.19527843e-08
+ 8.46909241e-07 1.19527845e-08 8.47009241e-07 1.19527842e-08 8.47109241e-07 1.19527845e-08 8.47209241e-07 1.19527842e-08 8.47309241e-07 1.19527844e-08 8.47409241e-07 1.19527845e-08 8.47509241e-07 1.19527847e-08 8.47609241e-07 1.19527846e-08
+ 8.47709241e-07 1.19527847e-08 8.47809241e-07 1.19527844e-08 8.47909241e-07 1.19527847e-08 8.48009241e-07 1.19527845e-08 8.48109241e-07 1.19527845e-08 8.48209241e-07 1.19527847e-08 8.48309241e-07 1.19527848e-08 8.48409241e-07 1.19527847e-08
+ 8.48509241e-07 1.19527847e-08 8.48609241e-07 1.19527845e-08 8.48709241e-07 1.19527849e-08 8.48809241e-07 1.19527847e-08 8.48909241e-07 1.19527849e-08 8.49009241e-07 1.19527846e-08 8.49109241e-07 1.1952785e-08 8.49209241e-07 1.19527847e-08
+ 8.49309241e-07 1.19527852e-08 8.49409241e-07 1.19527848e-08 8.49509241e-07 1.19527853e-08 8.49609241e-07 1.1952785e-08 8.49709241e-07 1.19527849e-08 8.49809241e-07 1.19527848e-08 8.49909241e-07 1.19527852e-08 8.50009241e-07 1.19527848e-08
+ 8.50109241e-07 1.19527852e-08 8.50209241e-07 1.19527852e-08 8.50309241e-07 1.1952785e-08 8.50409241e-07 1.19527852e-08 8.50509241e-07 1.19527852e-08 8.50609241e-07 1.1952785e-08 8.50709241e-07 1.19527854e-08 8.50809241e-07 1.19527852e-08
+ 8.50909241e-07 1.19527851e-08 8.51e-07 1.19527852e-08 8.5101e-07 1.1939096e-08 8.5103e-07 1.20196142e-08 8.5107e-07 1.18477351e-08 8.5115e-07 1.20721806e-08 8.5125e-07 1.18298608e-08 8.5135e-07 1.20694676e-08
+ 8.5145e-07 1.18519292e-08 8.5155e-07 1.20304652e-08 8.5165e-07 1.19012721e-08 8.5175e-07 1.19750946e-08 8.5185e-07 1.19638079e-08 8.51930828e-07 1.89264353e-07 8.52e-07 2.6011952e-07 8.52008608e-07 -7.14340553e-06
+ 8.52025825e-07 -6.92152579e-06 8.52060258e-07 1.22318635e-05 8.52106181e-07 -2.07308553e-07 8.52150081e-07 -6.86147133e-06 8.52198026e-07 -7.40021862e-07 8.5225538e-07 5.62676254e-06 8.52312019e-07 -4.8081976e-06 8.52404232e-07 3.76387955e-06
+ 8.52504232e-07 -3.03362411e-06 8.52604232e-07 2.49152677e-06 8.52704232e-07 -2.0066143e-06 8.52804232e-07 1.66419859e-06 8.52904232e-07 -1.34587456e-06 8.53004232e-07 1.13667787e-06 8.53104232e-07 -9.25169787e-07 8.53204232e-07 7.99904053e-07
+ 8.53304232e-07 -6.55185529e-07 8.53404232e-07 5.82278078e-07 8.53504232e-07 -4.79264614e-07 8.53604232e-07 4.39148788e-07 8.53704232e-07 -3.62367893e-07 8.53804232e-07 3.42983277e-07 8.53904232e-07 -2.82863542e-07 8.54004232e-07 2.7670735e-07
+ 8.54104232e-07 -2.27290234e-07 8.54204232e-07 2.29706838e-07 8.54304232e-07 -1.87298528e-07 8.54404232e-07 1.95374429e-07 8.54504232e-07 -1.5762143e-07 8.54604232e-07 1.69487684e-07 8.54704232e-07 -1.34878216e-07 8.54804232e-07 1.49328817e-07
+ 8.54904232e-07 -1.16888777e-07 8.55004232e-07 1.33147156e-07 8.55104232e-07 -1.02245866e-07 8.55204232e-07 1.19804709e-07 8.55304232e-07 -9.00265232e-08 8.55404232e-07 1.08549071e-07 8.55504232e-07 -7.96164004e-08 8.55604232e-07 9.88760457e-08
+ 8.55704232e-07 -7.05996945e-08 8.55804232e-07 9.04391845e-08 8.55904232e-07 -6.26865411e-08 8.56004232e-07 8.29959184e-08 8.56104232e-07 -5.56733953e-08 8.56204232e-07 7.63728477e-08 8.56304232e-07 -4.94109318e-08 8.56404232e-07 7.04403302e-08
+ 8.56504232e-07 -4.37857094e-08 8.56604232e-07 6.50985336e-08 8.56704232e-07 -3.87103505e-08 8.56804232e-07 6.02708226e-08 8.56904232e-07 -3.41165904e-08 8.57004232e-07 5.58953142e-08 8.57104232e-07 -2.99479537e-08 8.57204232e-07 5.19203753e-08
+ 8.57304232e-07 -2.61574241e-08 8.57404232e-07 4.83032379e-08 8.57504232e-07 -2.27059202e-08 8.57604232e-07 4.50079064e-08 8.57704232e-07 -1.95601254e-08 8.57804232e-07 4.20039857e-08 8.57904232e-07 -1.66928493e-08 8.58004232e-07 3.92662433e-08
+ 8.58104232e-07 -1.40797466e-08 8.58204232e-07 3.67710487e-08 8.58304232e-07 -1.16977539e-08 8.58404232e-07 3.44962388e-08 8.58504232e-07 -9.52592208e-09 8.58604232e-07 3.24219686e-08 8.58704232e-07 -7.54543122e-09 8.58804232e-07 3.05303505e-08
+ 8.58904232e-07 -5.73924311e-09 8.59004232e-07 2.88051113e-08 8.59104232e-07 -4.09181397e-09 8.59204232e-07 2.72314284e-08 8.59304232e-07 -2.58904997e-09 8.59404232e-07 2.57959147e-08 8.59504232e-07 -1.2182356e-09 8.59604232e-07 2.44864712e-08
+ 8.59704232e-07 3.19395066e-11 8.59804232e-07 2.32925139e-08 8.59904232e-07 1.16462462e-09 8.60004232e-07 2.22173191e-08 8.60104232e-07 2.18546928e-09 8.60204232e-07 2.12478758e-08 8.60304232e-07 3.10627829e-09 8.60404232e-07 2.03731003e-08
+ 8.60504232e-07 3.93746677e-09 8.60604232e-07 1.9583196e-08 8.60704232e-07 4.68825639e-09 8.60804232e-07 1.88694752e-08 8.60904232e-07 5.36683803e-09 8.61004232e-07 1.82242124e-08 8.61104232e-07 5.98050098e-09 8.61204232e-07 1.76405259e-08
+ 8.61304232e-07 6.53574517e-09 8.61404232e-07 1.7112274e-08 8.61504232e-07 7.03837574e-09 8.61604232e-07 1.66339684e-08 8.61704232e-07 7.49358273e-09 8.61804232e-07 1.62006999e-08 8.61904232e-07 7.90601179e-09 8.62004232e-07 1.58080698e-08
+ 8.62104232e-07 8.27982868e-09 8.62204232e-07 1.54521328e-08 8.62304232e-07 8.61876895e-09 8.62404232e-07 1.51293526e-08 8.62504232e-07 8.9261824e-09 8.62604232e-07 1.48365569e-08 8.62704232e-07 9.20506371e-09 8.62804232e-07 1.45709316e-08
+ 8.62904232e-07 9.45804962e-09 8.63004232e-07 1.43299974e-08 8.63104232e-07 9.68749889e-09 8.63204232e-07 1.41114864e-08 8.63304232e-07 9.8955979e-09 8.63404232e-07 1.39132948e-08 8.63504232e-07 1.00843647e-08 8.63604232e-07 1.3733493e-08
+ 8.63704232e-07 1.02556396e-08 8.63804232e-07 1.35703292e-08 8.63904232e-07 1.04110868e-08 8.64004232e-07 1.34221845e-08 8.64104232e-07 1.05522192e-08 8.64204232e-07 1.32880898e-08 8.64304232e-07 1.06794394e-08 8.64404232e-07 1.3166998e-08
+ 8.64504232e-07 1.07951332e-08 8.64604232e-07 1.30563922e-08 8.64704232e-07 1.09007877e-08 8.64804232e-07 1.29555431e-08 8.64904232e-07 1.09969994e-08 8.65004232e-07 1.28637763e-08 8.65104232e-07 1.10845362e-08 8.65204232e-07 1.27802766e-08
+ 8.65304232e-07 1.11641363e-08 8.65404232e-07 1.27044498e-08 8.65504232e-07 1.12363762e-08 8.65604232e-07 1.26355459e-08 8.65704232e-07 1.13021392e-08 8.65804232e-07 1.25728631e-08 8.65904232e-07 1.13617872e-08 8.66004232e-07 1.2516119e-08
+ 8.66104232e-07 1.14157952e-08 8.66204232e-07 1.24646918e-08 8.66304232e-07 1.14647825e-08 8.66404232e-07 1.24180176e-08 8.66504232e-07 1.15092592e-08 8.66604232e-07 1.23756302e-08 8.66704232e-07 1.1549659e-08 8.66804232e-07 1.23371224e-08
+ 8.66904232e-07 1.15863663e-08 8.67004232e-07 1.23021311e-08 8.67104232e-07 1.16197208e-08 8.67204232e-07 1.22703342e-08 8.67304232e-07 1.1650073e-08 8.67404232e-07 1.22412999e-08 8.67504232e-07 1.1677812e-08 8.67604232e-07 1.22148983e-08
+ 8.67704232e-07 1.17029104e-08 8.67804232e-07 1.21910169e-08 8.67904232e-07 1.17256512e-08 8.68004232e-07 1.21693517e-08 8.68104232e-07 1.17462983e-08 8.68204232e-07 1.21496707e-08 8.68304232e-07 1.17650611e-08 8.68404232e-07 1.21317818e-08
+ 8.68504232e-07 1.17821176e-08 8.68604232e-07 1.21155185e-08 8.68704232e-07 1.17976254e-08 8.68804232e-07 1.2100731e-08 8.68904232e-07 1.18117254e-08 8.69004232e-07 1.20872868e-08 8.69104232e-07 1.18245444e-08 8.69204232e-07 1.20750639e-08
+ 8.69304232e-07 1.18361992e-08 8.69404232e-07 1.20639507e-08 8.69504232e-07 1.1846796e-08 8.69604232e-07 1.20538463e-08 8.69704232e-07 1.18564304e-08 8.69804232e-07 1.204466e-08 8.69904232e-07 1.18651896e-08 8.70004232e-07 1.20363081e-08
+ 8.70104232e-07 1.18731534e-08 8.70204232e-07 1.20287149e-08 8.70304232e-07 1.18803934e-08 8.70404232e-07 1.20218112e-08 8.70504232e-07 1.1886976e-08 8.70604232e-07 1.20155351e-08 8.70704232e-07 1.18929603e-08 8.70804232e-07 1.20098293e-08
+ 8.70904232e-07 1.1898401e-08 8.71004232e-07 1.20046417e-08 8.71104232e-07 1.19033473e-08 8.71204232e-07 1.19999249e-08 8.71304232e-07 1.19078448e-08 8.71404232e-07 1.19956369e-08 8.71504232e-07 1.19119332e-08 8.71604232e-07 1.19917385e-08
+ 8.71704232e-07 1.191565e-08 8.71804232e-07 1.1988195e-08 8.71904232e-07 1.19190287e-08 8.72004232e-07 1.19849735e-08 8.72104232e-07 1.19221003e-08 8.72204232e-07 1.19820448e-08 8.72304232e-07 1.19248928e-08 8.72404232e-07 1.19793827e-08
+ 8.72504232e-07 1.19274312e-08 8.72604232e-07 1.19769624e-08 8.72704232e-07 1.19297385e-08 8.72804232e-07 1.19747623e-08 8.72904232e-07 1.19318362e-08 8.73004232e-07 1.19727623e-08 8.73104232e-07 1.19337436e-08 8.73204232e-07 1.1970944e-08
+ 8.73304232e-07 1.19354769e-08 8.73404232e-07 1.19692911e-08 8.73504232e-07 1.19370528e-08 8.73604232e-07 1.19677885e-08 8.73704232e-07 1.19384858e-08 8.73804232e-07 1.19664224e-08 8.73904232e-07 1.19397881e-08 8.74004232e-07 1.19651806e-08
+ 8.74104232e-07 1.19409723e-08 8.74204232e-07 1.19640516e-08 8.74304232e-07 1.19420486e-08 8.74404232e-07 1.19630253e-08 8.74504232e-07 1.19430267e-08 8.74604232e-07 1.19620927e-08 8.74704232e-07 1.19439165e-08 8.74804232e-07 1.19612445e-08
+ 8.74904232e-07 1.1944725e-08 8.75004232e-07 1.19604737e-08 8.75104232e-07 1.19454599e-08 8.75204232e-07 1.19597725e-08 8.75304232e-07 1.19461282e-08 8.75404232e-07 1.19591356e-08 8.75504232e-07 1.1946736e-08 8.75604232e-07 1.19585565e-08
+ 8.75704232e-07 1.19472882e-08 8.75804232e-07 1.19580296e-08 8.75904232e-07 1.19477901e-08 8.76004232e-07 1.19575514e-08 8.76104232e-07 1.19482464e-08 8.76204232e-07 1.1957116e-08 8.76304232e-07 1.19486612e-08 8.76404232e-07 1.19567207e-08
+ 8.76504232e-07 1.19490384e-08 8.76604232e-07 1.19563608e-08 8.76704232e-07 1.19493813e-08 8.76804232e-07 1.19560341e-08 8.76904232e-07 1.1949693e-08 8.77004232e-07 1.19557371e-08 8.77104232e-07 1.1949976e-08 8.77204232e-07 1.19554669e-08
+ 8.77304232e-07 1.19502337e-08 8.77404232e-07 1.19552215e-08 8.77504232e-07 1.19504676e-08 8.77604232e-07 1.19549983e-08 8.77704232e-07 1.19506808e-08 8.77804232e-07 1.19547953e-08 8.77904232e-07 1.19508739e-08 8.78004232e-07 1.19546109e-08
+ 8.78104232e-07 1.19510499e-08 8.78204232e-07 1.19544433e-08 8.78304232e-07 1.19512097e-08 8.78404232e-07 1.19542909e-08 8.78504232e-07 1.19513548e-08 8.78604232e-07 1.19541528e-08 8.78704232e-07 1.19514867e-08 8.78804232e-07 1.19540273e-08
+ 8.78904232e-07 1.19516066e-08 8.79004232e-07 1.1953913e-08 8.79104232e-07 1.1951715e-08 8.79204232e-07 1.19538095e-08 8.79304232e-07 1.19518137e-08 8.79404232e-07 1.19537153e-08 8.79504232e-07 1.19519035e-08 8.79604232e-07 1.19536299e-08
+ 8.79704232e-07 1.19519847e-08 8.79804232e-07 1.19535525e-08 8.79904232e-07 1.19520585e-08 8.80004232e-07 1.19534822e-08 8.80104232e-07 1.19521253e-08 8.80204232e-07 1.19534188e-08 8.80304232e-07 1.19521864e-08 8.80404232e-07 1.19533604e-08
+ 8.80504232e-07 1.19522416e-08 8.80604232e-07 1.19533082e-08 8.80704232e-07 1.19522917e-08 8.80804232e-07 1.19532601e-08 8.80904232e-07 1.19523371e-08 8.81004232e-07 1.19532169e-08 8.81104232e-07 1.19523785e-08 8.81204232e-07 1.19531776e-08
+ 8.81304232e-07 1.1952416e-08 8.81404232e-07 1.19531418e-08 8.81504232e-07 1.195245e-08 8.81604232e-07 1.19531093e-08 8.81704232e-07 1.19524809e-08 8.81804232e-07 1.19530799e-08 8.81904232e-07 1.1952509e-08 8.82004232e-07 1.19530532e-08
+ 8.82104232e-07 1.19525344e-08 8.82204232e-07 1.19530287e-08 8.82304232e-07 1.19525577e-08 8.82404232e-07 1.19530068e-08 8.82504232e-07 1.19525784e-08 8.82604232e-07 1.19529871e-08 8.82704232e-07 1.19525976e-08 8.82804232e-07 1.1952969e-08
+ 8.82904232e-07 1.19526148e-08 8.83004232e-07 1.19529523e-08 8.83104232e-07 1.19526307e-08 8.83204232e-07 1.19529374e-08 8.83304232e-07 1.1952645e-08 8.83404232e-07 1.19529235e-08 8.83504232e-07 1.19526579e-08 8.83604232e-07 1.19529114e-08
+ 8.83704232e-07 1.195267e-08 8.83804232e-07 1.19529e-08 8.83904232e-07 1.19526803e-08 8.84004232e-07 1.195289e-08 8.84104232e-07 1.19526904e-08 8.84204232e-07 1.19528807e-08 8.84304232e-07 1.1952699e-08 8.84404232e-07 1.19528722e-08
+ 8.84504232e-07 1.19527073e-08 8.84604232e-07 1.19528643e-08 8.84704232e-07 1.19527148e-08 8.84804232e-07 1.19528572e-08 8.84904232e-07 1.19527212e-08 8.85004232e-07 1.1952851e-08 8.85104232e-07 1.19527273e-08 8.85204232e-07 1.19528455e-08
+ 8.85304232e-07 1.19527329e-08 8.85404232e-07 1.19528399e-08 8.85504232e-07 1.19527379e-08 8.85604232e-07 1.19528353e-08 8.85704232e-07 1.19527426e-08 8.85804232e-07 1.19528309e-08 8.85904232e-07 1.19527464e-08 8.86004232e-07 1.1952827e-08
+ 8.86104232e-07 1.19527503e-08 8.86204232e-07 1.19528234e-08 8.86304232e-07 1.1952754e-08 8.86404232e-07 1.19528198e-08 8.86504232e-07 1.19527571e-08 8.86604232e-07 1.19528169e-08 8.86704232e-07 1.19527598e-08 8.86804232e-07 1.19528142e-08
+ 8.86904232e-07 1.19527623e-08 8.87004232e-07 1.19528118e-08 8.87104232e-07 1.19527647e-08 8.87204232e-07 1.19528098e-08 8.87304232e-07 1.19527666e-08 8.87404232e-07 1.19528078e-08 8.87504232e-07 1.19527685e-08 8.87604232e-07 1.19528058e-08
+ 8.87704232e-07 1.19527705e-08 8.87804232e-07 1.19528042e-08 8.87904232e-07 1.19527723e-08 8.88004232e-07 1.19528026e-08 8.88104232e-07 1.19527737e-08 8.88204232e-07 1.19528012e-08 8.88304232e-07 1.1952775e-08 8.88404232e-07 1.19528e-08
+ 8.88504232e-07 1.19527759e-08 8.88604232e-07 1.19527991e-08 8.88704232e-07 1.19527771e-08 8.88804232e-07 1.19527979e-08 8.88904232e-07 1.1952778e-08 8.89004232e-07 1.19527972e-08 8.89104232e-07 1.19527789e-08 8.89204232e-07 1.19527962e-08
+ 8.89304232e-07 1.19527797e-08 8.89404232e-07 1.19527954e-08 8.89504232e-07 1.19527806e-08 8.89604232e-07 1.19527946e-08 8.89704232e-07 1.19527813e-08 8.89804232e-07 1.19527938e-08 8.89904232e-07 1.19527817e-08 8.90004232e-07 1.19527935e-08
+ 8.90104232e-07 1.19527822e-08 8.90204232e-07 1.19527932e-08 8.90304232e-07 1.19527829e-08 8.90404232e-07 1.19527923e-08 8.90504232e-07 1.19527834e-08 8.90604232e-07 1.19527919e-08 8.90704232e-07 1.19527837e-08 8.90804232e-07 1.19527919e-08
+ 8.90904232e-07 1.19527841e-08 8.91004232e-07 1.19527914e-08 8.91104232e-07 1.19527847e-08 8.91204232e-07 1.19527907e-08 8.91304232e-07 1.19527851e-08 8.91404232e-07 1.19527907e-08 8.91504232e-07 1.19527851e-08 8.91604232e-07 1.19527901e-08
+ 8.91704232e-07 1.19527855e-08 8.91804232e-07 1.19527898e-08 8.91904232e-07 1.19527858e-08 8.92004232e-07 1.19527896e-08 8.92104232e-07 1.1952786e-08 8.92204232e-07 1.19527898e-08 8.92304232e-07 1.19527861e-08 8.92404232e-07 1.19527894e-08
+ 8.92504232e-07 1.19527863e-08 8.92604232e-07 1.19527894e-08 8.92704232e-07 1.19527864e-08 8.92804232e-07 1.19527892e-08 8.92904232e-07 1.19527867e-08 8.93004232e-07 1.19527889e-08 8.93104232e-07 1.19527869e-08 8.93204232e-07 1.19527889e-08
+ 8.93304232e-07 1.19527867e-08 8.93404232e-07 1.19527887e-08 8.93504232e-07 1.19527871e-08 8.93604232e-07 1.19527884e-08 8.93704232e-07 1.19527873e-08 8.93804232e-07 1.19527886e-08 8.93904232e-07 1.19527873e-08 8.94004232e-07 1.19527883e-08
+ 8.94104232e-07 1.19527874e-08 8.94204232e-07 1.19527885e-08 8.94304232e-07 1.19527871e-08 8.94404232e-07 1.19527885e-08 8.94504232e-07 1.19527874e-08 8.94604232e-07 1.19527881e-08 8.94704232e-07 1.19527874e-08 8.94804232e-07 1.19527883e-08
+ 8.94904232e-07 1.19527878e-08 8.95004232e-07 1.1952788e-08 8.95104232e-07 1.19527877e-08 8.95204232e-07 1.19527881e-08 8.95304232e-07 1.19527875e-08 8.95404232e-07 1.1952788e-08 8.95504232e-07 1.19527878e-08 8.95604232e-07 1.1952788e-08
+ 8.95704232e-07 1.19527875e-08 8.95804232e-07 1.19527881e-08 8.95904232e-07 1.19527876e-08 8.96004232e-07 1.19527881e-08 8.96104232e-07 1.19527877e-08 8.96204232e-07 1.1952788e-08 8.96304232e-07 1.19527878e-08 8.96404232e-07 1.1952788e-08
+ 8.96504232e-07 1.19527878e-08 8.96604232e-07 1.19527879e-08 8.96704232e-07 1.19527877e-08 8.96804232e-07 1.19527881e-08 8.96904232e-07 1.19527878e-08 8.97004232e-07 1.19527881e-08 8.97104232e-07 1.1952788e-08 8.97204232e-07 1.19527877e-08
+ 8.97304232e-07 1.19527879e-08 8.97404232e-07 1.1952788e-08 8.97504232e-07 1.1952788e-08 8.97604232e-07 1.19527879e-08 8.97704232e-07 1.1952788e-08 8.97804232e-07 1.19527879e-08 8.97904232e-07 1.19527877e-08 8.98004232e-07 1.19527881e-08
+ 8.98104232e-07 1.19527877e-08 8.98204232e-07 1.19527881e-08 8.98304232e-07 1.19527877e-08 8.98404232e-07 1.19527881e-08 8.98504232e-07 1.19527878e-08 8.98604232e-07 1.19527883e-08 8.98704232e-07 1.19527877e-08 8.98804232e-07 1.1952788e-08
+ 8.98904232e-07 1.19527877e-08 8.99004232e-07 1.19527882e-08 8.99104232e-07 1.19527876e-08 8.99204232e-07 1.19527884e-08 8.99304232e-07 1.19527877e-08 8.99404232e-07 1.19527881e-08 8.99504232e-07 1.19527877e-08 8.99604232e-07 1.19527885e-08
+ 8.99704232e-07 1.19527874e-08 8.99804232e-07 1.1952788e-08 8.99904232e-07 1.19527876e-08 9e-07 1.19527882e-08 9.0001e-07 1.19847867e-08 9.0003e-07 1.17957476e-08 9.0007e-07 1.21960664e-08 9.0015e-07 1.16790212e-08
+ 9.0025e-07 1.22357528e-08 9.0035e-07 1.16768705e-08 9.0045e-07 1.22053472e-08 9.0055e-07 1.17434326e-08 9.0065e-07 1.18632202e-08 9.0075e-07 2.60700188e-08 9.0085e-07 -6.67652971e-07 9.00932051e-07 4.41565399e-06
+ 9.01e-07 -1.00425785e-05 9.01008488e-07 -1.02352439e-05 9.01025463e-07 4.62438714e-06 9.01059414e-07 6.10068297e-06 9.0109062e-07 2.93430931e-06 9.0114347e-07 -1.23168869e-07 9.01199151e-07 8.33058792e-06 9.01299151e-07 -3.00514879e-05
+ 9.01399151e-07 0.000133952605 9.01499151e-07 -0.000207264225 9.01599151e-07 0.000192426471 9.01699151e-07 -0.000285523601 9.01799151e-07 0.000366852825 9.01893327e-07 -0.00036846974 9.01993327e-07 0.000376973588 9.02093327e-07 -0.000371315116
+ 9.02193327e-07 0.000359140809 9.02293327e-07 -0.000341874797 9.02393327e-07 0.000321770317 9.02493327e-07 -0.000299895372 9.02593327e-07 0.000277811836 9.02693327e-07 -0.000255845433 9.02793327e-07 0.000234952298 9.02893327e-07 -0.000215003446
+ 9.02993327e-07 0.000196566982 9.03093327e-07 -0.000179310692 9.03193327e-07 0.000163591693 9.03293327e-07 -0.000149019485 9.03393327e-07 0.0001358423 9.03493327e-07 -0.00012367801 9.03593327e-07 0.000112719887 9.03693327e-07 -0.000102618211
+ 9.03793327e-07 9.35370426e-05 9.03893327e-07 -8.51645593e-05 9.03993327e-07 7.76479395e-05 9.04093327e-07 -7.07110531e-05 9.04193327e-07 6.44902504e-05 9.04293327e-07 -5.87404539e-05 9.04393327e-07 5.35903595e-05 9.04493327e-07 -4.88209881e-05
+ 9.04593327e-07 4.45552201e-05 9.04693327e-07 -4.05956834e-05 9.04793327e-07 3.70606357e-05 9.04893327e-07 -3.37704863e-05 9.04993327e-07 3.08397242e-05 9.05093327e-07 -2.81033671e-05 9.05193327e-07 2.56727906e-05 9.05293327e-07 -2.33950168e-05
+ 9.05393327e-07 2.13788324e-05 9.05493327e-07 -1.94811354e-05 9.05593327e-07 1.78085526e-05 9.05693327e-07 -1.62261184e-05 9.05793327e-07 1.48386552e-05 9.05893327e-07 -1.35179108e-05 9.05993327e-07 1.23671987e-05 9.06093327e-07 -1.12638134e-05
+ 9.06193327e-07 1.03098066e-05 9.06293327e-07 -9.38706102e-06 9.06393327e-07 8.59657348e-06 9.06493327e-07 -7.824026e-06 9.06593327e-07 7.16953335e-06 9.06693327e-07 -6.48075399e-06 9.06793327e-07 5.98664906e-06 9.06893327e-07 -5.40521902e-06
+ 9.06993327e-07 4.99725389e-06 9.07093327e-07 -4.50840114e-06 9.07193327e-07 4.17217679e-06 9.07293327e-07 -3.76047466e-06 9.07393327e-07 3.48401778e-06 9.07493327e-07 -3.13661854e-06 9.07593327e-07 2.90996505e-06 9.07693327e-07 -2.61617076e-06
+ 9.07793327e-07 2.43102733e-06 9.07893327e-07 -2.18192815e-06 9.07993327e-07 2.04442042e-06 9.08093327e-07 -1.81749786e-06 9.08193327e-07 1.70770947e-06 9.08293327e-07 -1.51444849e-06 9.08393327e-07 1.42684781e-06 9.08493327e-07 -1.26166668e-06
+ 9.08593327e-07 1.1925578e-06 9.08693327e-07 -1.05078906e-06 9.08793327e-07 9.97096861e-07 9.08893327e-07 -8.74852071e-07 9.08993327e-07 8.34014161e-07 9.09093327e-07 -7.28053117e-07 9.09193327e-07 6.97935565e-07 9.09293327e-07 -6.05557653e-07
+ 9.09393327e-07 5.84381408e-07 9.09493327e-07 -5.03334641e-07 9.09593327e-07 4.89616695e-07 9.09693327e-07 -4.18023602e-07 9.09793327e-07 4.10527791e-07 9.09893327e-07 -3.46822422e-07 9.09993327e-07 3.44517445e-07 9.10093327e-07 -2.87393596e-07
+ 9.10193327e-07 2.89419645e-07 9.10293327e-07 -2.37788026e-07 9.10393327e-07 2.4342808e-07 9.10493327e-07 -1.96380018e-07 9.10593327e-07 2.05035977e-07 9.10693327e-07 -1.61813343e-07 9.10793327e-07 1.72986221e-07 9.10893327e-07 -1.32956444e-07
+ 9.10993327e-07 1.4622993e-07 9.11093327e-07 -1.08865152e-07 9.11193327e-07 1.23891857e-07 9.11293327e-07 -8.87516065e-08 9.11393327e-07 1.05241666e-07 9.11493327e-07 -7.19604539e-08 9.11593327e-07 8.96740331e-08 9.11693327e-07 -5.79459548e-08
+ 9.11793327e-07 7.668191e-08 9.11893327e-07 -4.62495987e-08 9.11993327e-07 6.58388038e-08 9.12093327e-07 -3.64880343e-08 9.12193327e-07 5.6789147e-08 9.12293327e-07 -2.83407877e-08 9.12393327e-07 4.92359388e-08 9.12493327e-07 -2.15406662e-08
+ 9.12593327e-07 4.29315531e-08 9.12693327e-07 -1.58507322e-08 9.12793327e-07 3.76566189e-08 9.12893327e-07 -1.11162829e-08 9.12993327e-07 3.32669802e-08 9.13093327e-07 -7.16407419e-09 9.13193327e-07 2.96027728e-08 9.13293327e-07 -3.86498894e-09
+ 9.13393327e-07 2.65440784e-08 9.13493327e-07 -1.11106224e-09 9.13593327e-07 2.39907998e-08 9.13693327e-07 1.1878297e-09 9.13793327e-07 2.18748402e-08 9.13893327e-07 3.09374734e-09 9.13993327e-07 2.01325726e-08 9.14093327e-07 4.66365546e-09
+ 9.14193327e-07 1.86974617e-08 9.14293327e-07 5.95680449e-09 9.14393327e-07 1.75153376e-08 9.14493327e-07 7.02199823e-09 9.14593327e-07 1.65415939e-08 9.14693327e-07 7.89942517e-09 9.14793327e-07 1.57394953e-08 9.14893327e-07 8.62218708e-09
+ 9.14993327e-07 1.49812768e-08 9.15093327e-07 9.20369131e-09 9.15193327e-07 1.44482747e-08 9.15293327e-07 9.68756114e-09 9.15393327e-07 1.40089631e-08 9.15493327e-07 1.00864089e-08 9.15593327e-07 1.36468572e-08 9.15693327e-07 1.04151539e-08
+ 9.15793327e-07 1.3348402e-08 9.15893327e-07 1.06861086e-08 9.15993327e-07 1.31024162e-08 9.16093327e-07 1.0909425e-08 9.16193327e-07 1.28996817e-08 9.16293327e-07 1.10934721e-08 9.16393327e-07 1.27326005e-08 9.16493327e-07 1.12451503e-08
+ 9.16593327e-07 1.25949073e-08 9.16693327e-07 1.13701465e-08 9.16793327e-07 1.24814388e-08 9.16893327e-07 1.1473149e-08 9.16993327e-07 1.23879381e-08 9.17093327e-07 1.15580224e-08 9.17193327e-07 1.23108973e-08 9.17293327e-07 1.16279524e-08
+ 9.17393327e-07 1.22474232e-08 9.17493327e-07 1.1685565e-08 9.17593327e-07 1.21951317e-08 9.17693327e-07 1.17330255e-08 9.17793327e-07 1.21520569e-08 9.17893327e-07 1.17721189e-08 9.17993327e-07 1.21165785e-08 9.18093327e-07 1.18043161e-08
+ 9.18193327e-07 1.20873597e-08 9.18293327e-07 1.18308303e-08 9.18393327e-07 1.20633014e-08 9.18493327e-07 1.18526595e-08 9.18593327e-07 1.20434953e-08 9.18693327e-07 1.18706288e-08 9.18793327e-07 1.20271934e-08 9.18893327e-07 1.1885417e-08
+ 9.18993327e-07 1.20137792e-08 9.19093327e-07 1.18975841e-08 9.19193327e-07 1.20027444e-08 9.19293327e-07 1.19075909e-08 9.19393327e-07 1.19936706e-08 9.19493327e-07 1.19158184e-08 9.19593327e-07 1.19862109e-08 9.19693327e-07 1.19225815e-08
+ 9.19793327e-07 1.19800805e-08 9.19893327e-07 1.19281375e-08 9.19993327e-07 1.19750458e-08 9.20093327e-07 1.19326991e-08 9.20193327e-07 1.19709136e-08 9.20293327e-07 1.19364418e-08 9.20393327e-07 1.19675242e-08 9.20493327e-07 1.19395104e-08
+ 9.20593327e-07 1.19647463e-08 9.20693327e-07 1.1942025e-08 9.20793327e-07 1.19624707e-08 9.20893327e-07 1.19440839e-08 9.20993327e-07 1.19606084e-08 9.21093327e-07 1.19457679e-08 9.21193327e-07 1.1959086e-08 9.21293327e-07 1.19471435e-08
+ 9.21393327e-07 1.19578434e-08 9.21493327e-07 1.1948266e-08 9.21593327e-07 1.19568301e-08 9.21693327e-07 1.19491802e-08 9.21793327e-07 1.19560053e-08 9.21893327e-07 1.19499239e-08 9.21993327e-07 1.19553351e-08 9.22093327e-07 1.19505276e-08
+ 9.22193327e-07 1.19547912e-08 9.22293327e-07 1.19510175e-08 9.22393327e-07 1.19543507e-08 9.22493327e-07 1.19514132e-08 9.22593327e-07 1.19539953e-08 9.22693327e-07 1.19517324e-08 9.22793327e-07 1.19537091e-08 9.22893327e-07 1.19519889e-08
+ 9.22993327e-07 1.19534794e-08 9.23093327e-07 1.19521943e-08 9.23193327e-07 1.19532955e-08 9.23293327e-07 1.19523583e-08 9.23393327e-07 1.19531493e-08 9.23493327e-07 1.19524883e-08 9.23593327e-07 1.1953034e-08 9.23693327e-07 1.19525906e-08
+ 9.23793327e-07 1.19529433e-08 9.23893327e-07 1.19526711e-08 9.23993327e-07 1.19528726e-08 9.24093327e-07 1.19527333e-08 9.24193327e-07 1.19528178e-08 9.24293327e-07 1.19527808e-08 9.24393327e-07 1.19527766e-08 9.24493327e-07 1.19528168e-08
+ 9.24593327e-07 1.19527452e-08 9.24693327e-07 1.19528438e-08 9.24793327e-07 1.19527225e-08 9.24893327e-07 1.19528631e-08 9.24993327e-07 1.19527063e-08 9.25093327e-07 1.19528764e-08 9.25193327e-07 1.19526952e-08 9.25293327e-07 1.19528853e-08
+ 9.25393327e-07 1.1952688e-08 9.25493327e-07 1.19528903e-08 9.25593327e-07 1.19526845e-08 9.25693327e-07 1.19528927e-08 9.25793327e-07 1.19526833e-08 9.25893327e-07 1.1952893e-08 9.25993327e-07 1.1952684e-08 9.26093327e-07 1.19528913e-08
+ 9.26193327e-07 1.19526863e-08 9.26293327e-07 1.19528888e-08 9.26393327e-07 1.19526892e-08 9.26493327e-07 1.19528853e-08 9.26593327e-07 1.19526931e-08 9.26693327e-07 1.19528814e-08 9.26793327e-07 1.19526976e-08 9.26893327e-07 1.19528767e-08
+ 9.26993327e-07 1.19527021e-08 9.27093327e-07 1.19528718e-08 9.27193327e-07 1.19527072e-08 9.27293327e-07 1.19528671e-08 9.27393327e-07 1.19527118e-08 9.27493327e-07 1.19528623e-08 9.27593327e-07 1.19527166e-08 9.27693327e-07 1.19528576e-08
+ 9.27793327e-07 1.19527213e-08 9.27893327e-07 1.1952853e-08 9.27993327e-07 1.19527259e-08 9.28093327e-07 1.19528482e-08 9.28193327e-07 1.19527305e-08 9.28293327e-07 1.19528438e-08 9.28393327e-07 1.19527349e-08 9.28493327e-07 1.19528397e-08
+ 9.28593327e-07 1.1952739e-08 9.28693327e-07 1.19528358e-08 9.28793327e-07 1.19527428e-08 9.28893327e-07 1.19528323e-08 9.28993327e-07 1.1952746e-08 9.29093327e-07 1.19528291e-08 9.29193327e-07 1.19527492e-08 9.29293327e-07 1.19528259e-08
+ 9.29393327e-07 1.19527525e-08 9.29493327e-07 1.19528227e-08 9.29593327e-07 1.19527555e-08 9.29693327e-07 1.195282e-08 9.29793327e-07 1.19527582e-08 9.29893327e-07 1.19528171e-08 9.29993327e-07 1.19527606e-08 9.30093327e-07 1.19528147e-08
+ 9.30193327e-07 1.19527628e-08 9.30293327e-07 1.19528125e-08 9.30393327e-07 1.19527651e-08 9.30493327e-07 1.19528103e-08 9.30593327e-07 1.1952767e-08 9.30693327e-07 1.19528086e-08 9.30793327e-07 1.19527689e-08 9.30893327e-07 1.19528068e-08
+ 9.30993327e-07 1.19527705e-08 9.31093327e-07 1.19528051e-08 9.31193327e-07 1.1952772e-08 9.31293327e-07 1.19528039e-08 9.31393327e-07 1.19527735e-08 9.31493327e-07 1.19528026e-08 9.31593327e-07 1.19527745e-08 9.31693327e-07 1.19528012e-08
+ 9.31793327e-07 1.19527758e-08 9.31893327e-07 1.19528002e-08 9.31993327e-07 1.19527769e-08 9.32093327e-07 1.19527993e-08 9.32193327e-07 1.19527777e-08 9.32293327e-07 1.19527985e-08 9.32393327e-07 1.19527785e-08 9.32493327e-07 1.19527976e-08
+ 9.32593327e-07 1.19527795e-08 9.32693327e-07 1.19527966e-08 9.32793327e-07 1.19527802e-08 9.32893327e-07 1.19527959e-08 9.32993327e-07 1.19527811e-08 9.33093327e-07 1.19527952e-08 9.33193327e-07 1.19527817e-08 9.33293327e-07 1.19527947e-08
+ 9.33393327e-07 1.19527823e-08 9.33493327e-07 1.19527941e-08 9.33593327e-07 1.19527828e-08 9.33693327e-07 1.19527935e-08 9.33793327e-07 1.19527831e-08 9.33893327e-07 1.19527932e-08 9.33993327e-07 1.19527837e-08 9.34093327e-07 1.19527928e-08
+ 9.34193327e-07 1.1952784e-08 9.34293327e-07 1.19527925e-08 9.34393327e-07 1.19527843e-08 9.34493327e-07 1.19527922e-08 9.34593327e-07 1.19527847e-08 9.34693327e-07 1.19527917e-08 9.34793327e-07 1.1952785e-08 9.34893327e-07 1.19527914e-08
+ 9.34993327e-07 1.19527853e-08 9.35093327e-07 1.19527912e-08 9.35193327e-07 1.19527857e-08 9.35293327e-07 1.19527911e-08 9.35393327e-07 1.19527858e-08 9.35493327e-07 1.19527906e-08 9.35593327e-07 1.19527862e-08 9.35693327e-07 1.19527905e-08
+ 9.35793327e-07 1.19527864e-08 9.35893327e-07 1.19527902e-08 9.35993327e-07 1.19527864e-08 9.36093327e-07 1.19527902e-08 9.36193327e-07 1.19527867e-08 9.36293327e-07 1.19527897e-08 9.36393327e-07 1.19527868e-08 9.36493327e-07 1.19527899e-08
+ 9.36593327e-07 1.19527868e-08 9.36693327e-07 1.19527898e-08 9.36793327e-07 1.19527868e-08 9.36893327e-07 1.19527898e-08 9.36993327e-07 1.19527869e-08 9.37093327e-07 1.19527895e-08 9.37193327e-07 1.1952787e-08 9.37293327e-07 1.19527895e-08
+ 9.37393327e-07 1.19527872e-08 9.37493327e-07 1.19527895e-08 9.37593327e-07 1.19527872e-08 9.37693327e-07 1.19527895e-08 9.37793327e-07 1.19527874e-08 9.37893327e-07 1.19527891e-08 9.37993327e-07 1.19527874e-08 9.38093327e-07 1.19527891e-08
+ 9.38193327e-07 1.19527873e-08 9.38293327e-07 1.19527894e-08 9.38393327e-07 1.19527875e-08 9.38493327e-07 1.1952789e-08 9.38593327e-07 1.19527876e-08 9.38693327e-07 1.19527889e-08 9.38793327e-07 1.19527877e-08 9.38893327e-07 1.19527888e-08
+ 9.38993327e-07 1.19527879e-08 9.39093327e-07 1.19527886e-08 9.39193327e-07 1.1952788e-08 9.39293327e-07 1.19527888e-08 9.39393327e-07 1.19527881e-08 9.39493327e-07 1.19527887e-08 9.39593327e-07 1.19527879e-08 9.39693327e-07 1.19527885e-08
+ 9.39793327e-07 1.19527879e-08 9.39893327e-07 1.19527886e-08 9.39993327e-07 1.19527879e-08 9.40093327e-07 1.19527889e-08 9.40193327e-07 1.19527878e-08 9.40293327e-07 1.1952789e-08 9.40393327e-07 1.19527878e-08 9.40493327e-07 1.19527887e-08
+ 9.40593327e-07 1.19527878e-08 9.40693327e-07 1.1952789e-08 9.40793327e-07 1.19527876e-08 9.40893327e-07 1.19527886e-08 9.40993327e-07 1.19527878e-08 9.41093327e-07 1.19527885e-08 9.41193327e-07 1.19527881e-08 9.41293327e-07 1.19527883e-08
+ 9.41393327e-07 1.19527878e-08 9.41493327e-07 1.19527886e-08 9.41593327e-07 1.19527881e-08 9.41693327e-07 1.19527886e-08 9.41793327e-07 1.19527881e-08 9.41893327e-07 1.19527888e-08 9.41993327e-07 1.1952788e-08 9.42093327e-07 1.19527888e-08
+ 9.42193327e-07 1.19527878e-08 9.42293327e-07 1.19527887e-08 9.42393327e-07 1.1952788e-08 9.42493327e-07 1.19527888e-08 9.42593327e-07 1.19527878e-08 9.42693327e-07 1.19527883e-08 9.42793327e-07 1.19527879e-08 9.42893327e-07 1.19527884e-08
+ 9.42993327e-07 1.19527878e-08 9.43093327e-07 1.19527883e-08 9.43193327e-07 1.19527879e-08 9.43293327e-07 1.19527884e-08 9.43393327e-07 1.19527879e-08 9.43493327e-07 1.19527884e-08 9.43593327e-07 1.19527878e-08 9.43693327e-07 1.19527884e-08
+ 9.43793327e-07 1.19527879e-08 9.43893327e-07 1.19527885e-08 9.43993327e-07 1.19527878e-08 9.44093327e-07 1.19527883e-08 9.44193327e-07 1.1952788e-08 9.44293327e-07 1.19527883e-08 9.44393327e-07 1.1952788e-08 9.44493327e-07 1.19527883e-08
+ 9.44593327e-07 1.19527881e-08 9.44693327e-07 1.19527883e-08 9.44793327e-07 1.19527878e-08 9.44893327e-07 1.19527883e-08 9.44993327e-07 1.19527881e-08 9.45093327e-07 1.19527884e-08 9.45193327e-07 1.1952788e-08 9.45293327e-07 1.19527885e-08
+ 9.45393327e-07 1.1952788e-08 9.45493327e-07 1.19527884e-08 9.45593327e-07 1.19527881e-08 9.45693327e-07 1.19527884e-08 9.45793327e-07 1.1952788e-08 9.45893327e-07 1.19527885e-08 9.45993327e-07 1.19527879e-08 9.46093327e-07 1.19527885e-08
+ 9.46193327e-07 1.19527878e-08 9.46293327e-07 1.19527885e-08 9.46393327e-07 1.19527879e-08 9.46493327e-07 1.19527885e-08 9.46593327e-07 1.19527878e-08 9.46693327e-07 1.19527885e-08 9.46793327e-07 1.1952788e-08 9.46893327e-07 1.19527886e-08
+ 9.46993327e-07 1.19527882e-08 9.47093327e-07 1.19527886e-08 9.47193327e-07 1.19527882e-08 9.47293327e-07 1.19527885e-08 9.47393327e-07 1.19527881e-08 9.47493327e-07 1.19527882e-08 9.47593327e-07 1.19527879e-08 9.47693327e-07 1.19527883e-08
+ 9.47793327e-07 1.19527881e-08 9.47893327e-07 1.19527882e-08 9.47993327e-07 1.19527879e-08 9.48093327e-07 1.19527883e-08 9.48193327e-07 1.19527879e-08 9.48293327e-07 1.19527885e-08 9.48393327e-07 1.1952788e-08 9.48493327e-07 1.19527884e-08
+ 9.48593327e-07 1.19527881e-08 9.48693327e-07 1.19527882e-08 9.48793327e-07 1.1952788e-08 9.48893327e-07 1.19527882e-08 9.48993327e-07 1.19527881e-08 9.49093327e-07 1.19527882e-08 9.49193327e-07 1.19527882e-08 9.49293327e-07 1.19527883e-08
+ 9.49393327e-07 1.19527881e-08 9.49493327e-07 1.19527883e-08 9.49593327e-07 1.19527881e-08 9.49693327e-07 1.1952788e-08 9.49793327e-07 1.19527881e-08 9.49893327e-07 1.19527881e-08 9.49993327e-07 1.19527882e-08 9.50093327e-07 1.19527881e-08
+ 9.50193327e-07 1.19527881e-08 9.50293327e-07 1.19527881e-08 9.50393327e-07 1.19527882e-08 9.50493327e-07 1.19527881e-08 9.50593327e-07 1.19527882e-08 9.50693327e-07 1.19527881e-08 9.50793327e-07 1.19527883e-08 9.50893327e-07 1.19527881e-08
+ 9.50993327e-07 1.19527882e-08 9.51e-07 1.19527874e-08 9.5101e-07 1.19399424e-08 9.5103e-07 1.20150128e-08 9.5107e-07 1.18559368e-08 9.5115e-07 1.20621033e-08 9.5125e-07 1.18410984e-08 9.5135e-07 1.20574882e-08
+ 9.5145e-07 1.18638216e-08 9.5155e-07 1.20197039e-08 9.5165e-07 1.19101577e-08 9.5175e-07 1.19686134e-08 9.5185e-07 1.1967486e-08 9.51930828e-07 1.83418271e-07 9.52e-07 1.06002517e-07 9.52008608e-07 -6.35218173e-06
+ 9.52025825e-07 -6.40058733e-06 9.52060258e-07 9.75152962e-06 9.52106188e-07 5.28435492e-06 9.52150118e-07 -1.51923671e-05 9.5219811e-07 6.42629664e-06 9.52255501e-07 9.57222351e-07 9.52312176e-07 -1.57314433e-06 9.52404431e-07 1.13652367e-06
+ 9.52490774e-07 -1.00482103e-06 9.52590774e-07 9.71186728e-07 9.52690774e-07 -8.68547259e-07 9.52790774e-07 8.16808096e-07 9.52890774e-07 -7.24287651e-07 9.52990774e-07 6.88965999e-07 9.53090774e-07 -6.14052292e-07 9.53190774e-07 5.94787164e-07
+ 9.53290774e-07 -5.33642225e-07 9.53390774e-07 5.25529847e-07 9.53490774e-07 -4.73285723e-07 9.53590774e-07 4.72036289e-07 9.53690774e-07 -4.25085269e-07 9.53790774e-07 4.27835408e-07 9.53890774e-07 -3.83953563e-07 9.53990774e-07 3.89048055e-07
+ 9.54090774e-07 -3.4701833e-07 9.54190774e-07 3.53603078e-07 9.54290774e-07 -3.12840629e-07 9.54390774e-07 3.20537789e-07 9.54490774e-07 -2.80809747e-07 9.54590774e-07 2.89491019e-07 9.54690774e-07 -2.50738347e-07 9.54790774e-07 2.60389507e-07
+ 9.54890774e-07 -2.2262413e-07 9.54990774e-07 2.33269734e-07 9.55090774e-07 -1.96520033e-07 9.55190774e-07 2.08185539e-07 9.55290774e-07 -1.72470285e-07 9.55390774e-07 1.85165182e-07 9.55490774e-07 -1.50484079e-07 9.55590774e-07 1.64198319e-07
+ 9.55690774e-07 -1.30531642e-07 9.55790774e-07 1.45236542e-07 9.55890774e-07 -1.12547054e-07 9.55990774e-07 1.28198328e-07 9.56090774e-07 -9.64351094e-08 9.56190774e-07 1.12976947e-07 9.56290774e-07 -8.20795775e-08 9.56390774e-07 9.94489937e-08
+ 9.56490774e-07 -6.93520122e-08 9.56590774e-07 8.74825732e-08 9.56690774e-07 -5.81182252e-08 9.56790774e-07 7.69425247e-08 9.56890774e-07 -4.82432947e-08 9.56990774e-07 6.76957224e-08 9.57090774e-07 -3.95973199e-08 9.57190774e-07 5.96159692e-08
+ 9.57290774e-07 -3.20580335e-08 9.57390774e-07 5.2583098e-08 9.57490774e-07 -2.55059463e-08 9.57590774e-07 4.64804052e-08 9.57690774e-07 -1.98288253e-08 9.57790774e-07 4.12000749e-08 9.57890774e-07 -1.49233088e-08 9.57990774e-07 3.6643222e-08
+ 9.58090774e-07 -1.06952403e-08 9.58190774e-07 3.27205767e-08 9.58290774e-07 -7.06015074e-09 9.58390774e-07 2.93521472e-08 9.58490774e-07 -3.94241798e-09 9.58590774e-07 2.64666448e-08 9.58690774e-07 -1.27496944e-09 9.58790774e-07 2.40008381e-08
+ 9.58890774e-07 9.95358129e-10 9.58990774e-07 2.19105881e-08 9.59090774e-07 2.9111219e-09 9.59190774e-07 2.01552985e-08 9.59290774e-07 4.51850554e-09 9.59390774e-07 1.86841675e-08 9.59490774e-07 5.86417134e-09 9.59590774e-07 1.74539926e-08
+ 9.59690774e-07 6.98806979e-09 9.59790774e-07 1.64278639e-08 9.59890774e-07 7.9243051e-09 9.59990774e-07 1.55742174e-08 9.60090774e-07 8.70212052e-09 9.60190774e-07 1.48659897e-08 9.60290774e-07 9.346525e-09 9.60390774e-07 1.42800906e-08
+ 9.60490774e-07 9.87882079e-09 9.60590774e-07 1.37968806e-08 9.60690774e-07 1.03171054e-08 9.60790774e-07 1.33996929e-08 9.60890774e-07 1.06767188e-08 9.60990774e-07 1.30744149e-08 9.61090774e-07 1.0970639e-08 9.61190774e-07 1.28091175e-08
+ 9.61290774e-07 1.1209824e-08 9.61390774e-07 1.25937396e-08 9.61490774e-07 1.14035097e-08 9.61590774e-07 1.24198065e-08 9.61690774e-07 1.15594665e-08 9.61790774e-07 1.22801993e-08 9.61890774e-07 1.16842191e-08 9.61990774e-07 1.21689277e-08
+ 9.62090774e-07 1.17832642e-08 9.62190774e-07 1.20809675e-08 9.62290774e-07 1.18611809e-08 9.62390774e-07 1.20121453e-08 9.62490774e-07 1.19217768e-08 9.62590774e-07 1.19589732e-08 9.62690774e-07 1.19682666e-08 9.62790774e-07 1.19184844e-08
+ 9.62890774e-07 1.20033726e-08 9.62990774e-07 1.18882068e-08 9.63090774e-07 1.20293198e-08 9.63190774e-07 1.18661404e-08 9.63290774e-07 1.20479118e-08 9.63390774e-07 1.18506557e-08 9.63490774e-07 1.20606223e-08 9.63590774e-07 1.1840417e-08
+ 9.63690774e-07 1.20686623e-08 9.63790774e-07 1.18343279e-08 9.63890774e-07 1.20729713e-08 9.63990774e-07 1.18315196e-08 9.64090774e-07 1.20748511e-08 9.64190774e-07 1.18303283e-08 9.64290774e-07 1.20750052e-08 9.64390774e-07 1.18314565e-08
+ 9.64490774e-07 1.20727117e-08 9.64590774e-07 1.18346006e-08 9.64690774e-07 1.20690051e-08 9.64790774e-07 1.18387676e-08 9.64890774e-07 1.20644243e-08 9.64990774e-07 1.18436873e-08 9.65090774e-07 1.2059238e-08 9.65190774e-07 1.18490772e-08
+ 9.65290774e-07 1.20536964e-08 9.65390774e-07 1.18547528e-08 9.65490774e-07 1.20478533e-08 9.65590774e-07 1.18607527e-08 9.65690774e-07 1.2041826e-08 9.65790774e-07 1.18666786e-08 9.65890774e-07 1.20360324e-08 9.65990774e-07 1.18723566e-08
+ 9.66090774e-07 1.20304576e-08 9.66190774e-07 1.18778302e-08 9.66290774e-07 1.20250903e-08 9.66390774e-07 1.18830857e-08 9.66490774e-07 1.20199506e-08 9.66590774e-07 1.18881049e-08 9.66690774e-07 1.20150551e-08 9.66790774e-07 1.18928746e-08
+ 9.66890774e-07 1.2010413e-08 9.66990774e-07 1.18973874e-08 9.67090774e-07 1.20060305e-08 9.67190774e-07 1.19016379e-08 9.67290774e-07 1.20019122e-08 9.67390774e-07 1.19056261e-08 9.67490774e-07 1.19980542e-08 9.67590774e-07 1.19093532e-08
+ 9.67690774e-07 1.19944569e-08 9.67790774e-07 1.19128236e-08 9.67890774e-07 1.19911095e-08 9.67990774e-07 1.19160511e-08 9.68090774e-07 1.19879988e-08 9.68190774e-07 1.1919048e-08 9.68290774e-07 1.19851133e-08 9.68390774e-07 1.19218414e-08
+ 9.68490774e-07 1.19823906e-08 9.68590774e-07 1.19244632e-08 9.68690774e-07 1.19799102e-08 9.68790774e-07 1.19268154e-08 9.68890774e-07 1.19776581e-08 9.68990774e-07 1.19289784e-08 9.69090774e-07 1.19755773e-08 9.69190774e-07 1.19309846e-08
+ 9.69290774e-07 1.19736416e-08 9.69390774e-07 1.19328462e-08 9.69490774e-07 1.19718592e-08 9.69590774e-07 1.19345513e-08 9.69690774e-07 1.19702255e-08 9.69790774e-07 1.19361176e-08 9.69890774e-07 1.19687261e-08 9.69990774e-07 1.1937551e-08
+ 9.70090774e-07 1.19673551e-08 9.70190774e-07 1.19388626e-08 9.70290774e-07 1.19661e-08 9.70390774e-07 1.19400644e-08 9.70490774e-07 1.19649494e-08 9.70590774e-07 1.19411661e-08 9.70690774e-07 1.19638948e-08 9.70790774e-07 1.19421753e-08
+ 9.70890774e-07 1.19629286e-08 9.70990774e-07 1.19431e-08 9.71090774e-07 1.19620445e-08 9.71190774e-07 1.19439457e-08 9.71290774e-07 1.19612351e-08 9.71390774e-07 1.19447195e-08 9.71490774e-07 1.19604954e-08 9.71590774e-07 1.19454268e-08
+ 9.71690774e-07 1.19598198e-08 9.71790774e-07 1.19460721e-08 9.71890774e-07 1.19592033e-08 9.71990774e-07 1.19466611e-08 9.72090774e-07 1.19586407e-08 9.72190774e-07 1.1947198e-08 9.72290774e-07 1.19581278e-08 9.72390774e-07 1.19476887e-08
+ 9.72490774e-07 1.1957659e-08 9.72590774e-07 1.19481361e-08 9.72690774e-07 1.19572318e-08 9.72790774e-07 1.19485442e-08 9.72890774e-07 1.19568417e-08 9.72990774e-07 1.19489169e-08 9.73090774e-07 1.19564857e-08 9.73190774e-07 1.1949257e-08
+ 9.73290774e-07 1.19561603e-08 9.73390774e-07 1.19495684e-08 9.73490774e-07 1.19558632e-08 9.73590774e-07 1.19498513e-08 9.73690774e-07 1.19555937e-08 9.73790774e-07 1.1950109e-08 9.73890774e-07 1.19553472e-08 9.73990774e-07 1.19503444e-08
+ 9.74090774e-07 1.1955122e-08 9.74190774e-07 1.195056e-08 9.74290774e-07 1.19549159e-08 9.74390774e-07 1.19507568e-08 9.74490774e-07 1.19547275e-08 9.74590774e-07 1.1950937e-08 9.74690774e-07 1.19545553e-08 9.74790774e-07 1.19511016e-08
+ 9.74890774e-07 1.19543979e-08 9.74990774e-07 1.19512522e-08 9.75090774e-07 1.1954254e-08 9.75190774e-07 1.19513895e-08 9.75290774e-07 1.19541227e-08 9.75390774e-07 1.1951515e-08 9.75490774e-07 1.19540033e-08 9.75590774e-07 1.19516285e-08
+ 9.75690774e-07 1.1953895e-08 9.75790774e-07 1.19517321e-08 9.75890774e-07 1.19537962e-08 9.75990774e-07 1.19518265e-08 9.76090774e-07 1.19537055e-08 9.76190774e-07 1.19519135e-08 9.76290774e-07 1.19536224e-08 9.76390774e-07 1.1951993e-08
+ 9.76490774e-07 1.19535465e-08 9.76590774e-07 1.19520654e-08 9.76690774e-07 1.19534775e-08 9.76790774e-07 1.19521316e-08 9.76890774e-07 1.19534143e-08 9.76990774e-07 1.19521916e-08 9.77090774e-07 1.19533568e-08 9.77190774e-07 1.19522465e-08
+ 9.77290774e-07 1.19533047e-08 9.77390774e-07 1.19522965e-08 9.77490774e-07 1.19532568e-08 9.77590774e-07 1.19523424e-08 9.77690774e-07 1.19532131e-08 9.77790774e-07 1.19523835e-08 9.77890774e-07 1.19531735e-08 9.77990774e-07 1.19524214e-08
+ 9.78090774e-07 1.19531376e-08 9.78190774e-07 1.19524555e-08 9.78290774e-07 1.19531049e-08 9.78390774e-07 1.19524867e-08 9.78490774e-07 1.19530757e-08 9.78590774e-07 1.19525148e-08 9.78690774e-07 1.19530487e-08 9.78790774e-07 1.19525405e-08
+ 9.78890774e-07 1.19530241e-08 9.78990774e-07 1.19525636e-08 9.79090774e-07 1.19530023e-08 9.79190774e-07 1.19525846e-08 9.79290774e-07 1.19529825e-08 9.79390774e-07 1.19526033e-08 9.79490774e-07 1.19529643e-08 9.79590774e-07 1.19526207e-08
+ 9.79690774e-07 1.19529481e-08 9.79790774e-07 1.19526363e-08 9.79890774e-07 1.19529331e-08 9.79990774e-07 1.19526503e-08 9.80090774e-07 1.19529196e-08 9.80190774e-07 1.19526631e-08 9.80290774e-07 1.19529073e-08 9.80390774e-07 1.19526749e-08
+ 9.80490774e-07 1.19528963e-08 9.80590774e-07 1.19526855e-08 9.80690774e-07 1.19528865e-08 9.80790774e-07 1.19526948e-08 9.80890774e-07 1.19528774e-08 9.80990774e-07 1.19527034e-08 9.81090774e-07 1.1952869e-08 9.81190774e-07 1.19527114e-08
+ 9.81290774e-07 1.19528616e-08 9.81390774e-07 1.19527184e-08 9.81490774e-07 1.19528551e-08 9.81590774e-07 1.19527247e-08 9.81690774e-07 1.19528489e-08 9.81790774e-07 1.19527306e-08 9.81890774e-07 1.19528435e-08 9.81990774e-07 1.19527359e-08
+ 9.82090774e-07 1.19528386e-08 9.82190774e-07 1.19527405e-08 9.82290774e-07 1.19528339e-08 9.82390774e-07 1.1952745e-08 9.82490774e-07 1.19528296e-08 9.82590774e-07 1.19527488e-08 9.82690774e-07 1.1952826e-08 9.82790774e-07 1.19527527e-08
+ 9.82890774e-07 1.19528223e-08 9.82990774e-07 1.19527558e-08 9.83090774e-07 1.19528193e-08 9.83190774e-07 1.19527588e-08 9.83290774e-07 1.19528165e-08 9.83390774e-07 1.19527613e-08 9.83490774e-07 1.19528138e-08 9.83590774e-07 1.19527638e-08
+ 9.83690774e-07 1.19528118e-08 9.83790774e-07 1.19527658e-08 9.83890774e-07 1.19528094e-08 9.83990774e-07 1.19527682e-08 9.84090774e-07 1.19528076e-08 9.84190774e-07 1.19527697e-08 9.84290774e-07 1.19528059e-08 9.84390774e-07 1.19527714e-08
+ 9.84490774e-07 1.19528044e-08 9.84590774e-07 1.19527728e-08 9.84690774e-07 1.19528029e-08 9.84790774e-07 1.19527743e-08 9.84890774e-07 1.19528014e-08 9.84990774e-07 1.19527757e-08 9.85090774e-07 1.19528004e-08 9.85190774e-07 1.19527767e-08
+ 9.85290774e-07 1.19527994e-08 9.85390774e-07 1.19527778e-08 9.85490774e-07 1.19527985e-08 9.85590774e-07 1.19527787e-08 9.85690774e-07 1.19527974e-08 9.85790774e-07 1.19527794e-08 9.85890774e-07 1.19527966e-08 9.85990774e-07 1.19527803e-08
+ 9.86090774e-07 1.19527959e-08 9.86190774e-07 1.1952781e-08 9.86290774e-07 1.19527952e-08 9.86390774e-07 1.19527815e-08 9.86490774e-07 1.19527946e-08 9.86590774e-07 1.19527822e-08 9.86690774e-07 1.19527941e-08 9.86790774e-07 1.19527825e-08
+ 9.86890774e-07 1.19527936e-08 9.86990774e-07 1.1952783e-08 9.87090774e-07 1.19527932e-08 9.87190774e-07 1.19527835e-08 9.87290774e-07 1.19527929e-08 9.87390774e-07 1.1952784e-08 9.87490774e-07 1.19527924e-08 9.87590774e-07 1.19527844e-08
+ 9.87690774e-07 1.1952792e-08 9.87790774e-07 1.19527846e-08 9.87890774e-07 1.1952792e-08 9.87990774e-07 1.19527848e-08 9.88090774e-07 1.19527917e-08 9.88190774e-07 1.1952785e-08 9.88290774e-07 1.19527916e-08 9.88390774e-07 1.19527853e-08
+ 9.88490774e-07 1.19527913e-08 9.88590774e-07 1.19527856e-08 9.88690774e-07 1.1952791e-08 9.88790774e-07 1.19527858e-08 9.88890774e-07 1.19527907e-08 9.88990774e-07 1.19527861e-08 9.89090774e-07 1.19527905e-08 9.89190774e-07 1.19527862e-08
+ 9.89290774e-07 1.19527901e-08 9.89390774e-07 1.19527866e-08 9.89490774e-07 1.19527899e-08 9.89590774e-07 1.19527869e-08 9.89690774e-07 1.19527899e-08 9.89790774e-07 1.19527868e-08 9.89890774e-07 1.19527899e-08 9.89990774e-07 1.19527868e-08
+ 9.90090774e-07 1.19527898e-08 9.90190774e-07 1.19527869e-08 9.90290774e-07 1.19527897e-08 9.90390774e-07 1.1952787e-08 9.90490774e-07 1.19527896e-08 9.90590774e-07 1.1952787e-08 9.90690774e-07 1.19527897e-08 9.90790774e-07 1.19527871e-08
+ 9.90890774e-07 1.19527893e-08 9.90990774e-07 1.19527873e-08 9.91090774e-07 1.19527892e-08 9.91190774e-07 1.19527874e-08 9.91290774e-07 1.19527892e-08 9.91390774e-07 1.19527875e-08 9.91490774e-07 1.19527891e-08 9.91590774e-07 1.19527877e-08
+ 9.91690774e-07 1.1952789e-08 9.91790774e-07 1.19527877e-08 9.91890774e-07 1.19527889e-08 9.91990774e-07 1.19527875e-08 9.92090774e-07 1.19527889e-08 9.92190774e-07 1.19527877e-08 9.92290774e-07 1.19527891e-08 9.92390774e-07 1.19527878e-08
+ 9.92490774e-07 1.1952789e-08 9.92590774e-07 1.19527877e-08 9.92690774e-07 1.19527887e-08 9.92790774e-07 1.19527879e-08 9.92890774e-07 1.19527889e-08 9.92990774e-07 1.19527878e-08 9.93090774e-07 1.19527887e-08 9.93190774e-07 1.19527878e-08
+ 9.93290774e-07 1.1952789e-08 9.93390774e-07 1.19527877e-08 9.93490774e-07 1.19527891e-08 9.93590774e-07 1.19527876e-08 9.93690774e-07 1.1952789e-08 9.93790774e-07 1.19527876e-08 9.93890774e-07 1.19527888e-08 9.93990774e-07 1.19527877e-08
+ 9.94090774e-07 1.19527891e-08 9.94190774e-07 1.19527877e-08 9.94290774e-07 1.19527891e-08 9.94390774e-07 1.19527875e-08 9.94490774e-07 1.19527886e-08 9.94590774e-07 1.19527878e-08 9.94690774e-07 1.19527886e-08 9.94790774e-07 1.19527881e-08
+ 9.94890774e-07 1.19527887e-08 9.94990774e-07 1.19527881e-08 9.95090774e-07 1.19527886e-08 9.95190774e-07 1.1952788e-08 9.95290774e-07 1.19527885e-08 9.95390774e-07 1.19527878e-08 9.95490774e-07 1.19527885e-08 9.95590774e-07 1.19527879e-08
+ 9.95690774e-07 1.19527884e-08 9.95790774e-07 1.19527879e-08 9.95890774e-07 1.19527883e-08 9.95990774e-07 1.19527878e-08 9.96090774e-07 1.19527885e-08 9.96190774e-07 1.19527878e-08 9.96290774e-07 1.19527885e-08 9.96390774e-07 1.19527878e-08
+ 9.96490774e-07 1.19527885e-08 9.96590774e-07 1.1952788e-08 9.96690774e-07 1.19527888e-08 9.96790774e-07 1.1952788e-08 9.96890774e-07 1.19527886e-08 9.96990774e-07 1.19527881e-08 9.97090774e-07 1.19527886e-08 9.97190774e-07 1.19527882e-08
+ 9.97290774e-07 1.19527883e-08 9.97390774e-07 1.1952788e-08 9.97490774e-07 1.19527883e-08 9.97590774e-07 1.1952788e-08 9.97690774e-07 1.19527881e-08 9.97790774e-07 1.19527881e-08 9.97890774e-07 1.19527881e-08 9.97990774e-07 1.19527882e-08
+ 9.98090774e-07 1.19527882e-08 9.98190774e-07 1.19527881e-08 9.98290774e-07 1.19527882e-08 9.98390774e-07 1.19527881e-08 9.98490774e-07 1.19527881e-08 9.98590774e-07 1.19527881e-08 9.98690774e-07 1.19527883e-08 9.98790774e-07 1.19527881e-08
+ 9.98890774e-07 1.19527883e-08 9.98990774e-07 1.19527883e-08 9.99090774e-07 1.19527881e-08 9.99190774e-07 1.19527882e-08 9.99290774e-07 1.1952788e-08 9.99390774e-07 1.19527883e-08 9.99490774e-07 1.1952788e-08 9.99590774e-07 1.19527883e-08
+ 9.99690774e-07 1.19527881e-08 9.99790774e-07 1.19527881e-08 9.99890774e-07 1.19527882e-08 9.99990774e-07 1.19527881e-08 1e-06 1.19527879e-08 )
* Beban sederhana: hanya resistor biar ada arus
Rload in 0 1k

* Simulasi transient
.tran 0.1n 1u
.control
* Plot hasil
run
plot v(in) v(in2)+5 v(in4)+10
.endc
.end
