* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__pfet_20v0__toxe_mult = 0.948
+ sky130_fd_pr__pfet_20v0__rshn_mult = 1.0
+ sky130_fd_pr__pfet_20v0__overlap_mult = 0.10
+ sky130_fd_pr__pfet_20v0__ajunction_mult = 9.3222e-1
+ sky130_fd_pr__pfet_20v0__pjunction_mult = 9.4436e-1
+ sky130_fd_pr__pfet_20v0__lint_diff = 1.7325e-8
+ sky130_fd_pr__pfet_20v0__wint_diff = -3.2175e-8
+ sky130_fd_pr__pfet_20v0__dlc_diff = 8.7000e-8
+ sky130_fd_pr__pfet_20v0__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__pfet_20v0, Bin 000, W = 30.0, L = 1.0
* -----------------------------------
.param
+ sky130_fd_pr__pfet_20v0__rdrift_mult = 7.4899e-1
+ sky130_fd_pr__pfet_20v0__vth0_diff = 2.2906e-1
+ sky130_fd_pr__pfet_20v0__u0_diff = 1.1548e-2
+ sky130_fd_pr__pfet_20v0__k2_diff = 0.0
+ sky130_fd_pr__pfet_20v0__agidl_diff = 0.0
.include "sky130_fd_pr__pfet_20v0__subcircuit.pm3.spice"
