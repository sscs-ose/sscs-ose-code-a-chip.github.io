magic
tech sky130A
magscale 1 2
timestamp 1762074413
<< pwell >>
rect -276 -610 276 610
<< nmos >>
rect -80 -400 80 400
<< ndiff >>
rect -138 388 -80 400
rect -138 -388 -126 388
rect -92 -388 -80 388
rect -138 -400 -80 -388
rect 80 388 138 400
rect 80 -388 92 388
rect 126 -388 138 388
rect 80 -400 138 -388
<< ndiffc >>
rect -126 -388 -92 388
rect 92 -388 126 388
<< psubdiff >>
rect -240 540 -144 574
rect 144 540 240 574
rect -240 478 -206 540
rect 206 478 240 540
rect -240 -540 -206 -478
rect 206 -540 240 -478
rect -240 -574 -144 -540
rect 144 -574 240 -540
<< psubdiffcont >>
rect -144 540 144 574
rect -240 -478 -206 478
rect 206 -478 240 478
rect -144 -574 144 -540
<< poly >>
rect -80 472 80 488
rect -80 438 -64 472
rect 64 438 80 472
rect -80 400 80 438
rect -80 -438 80 -400
rect -80 -472 -64 -438
rect 64 -472 80 -438
rect -80 -488 80 -472
<< polycont >>
rect -64 438 64 472
rect -64 -472 64 -438
<< locali >>
rect -240 540 -144 574
rect 144 540 240 574
rect -240 478 -206 540
rect 206 478 240 540
rect -80 438 -64 472
rect 64 438 80 472
rect -126 388 -92 404
rect -126 -404 -92 -388
rect 92 388 126 404
rect 92 -404 126 -388
rect -80 -472 -64 -438
rect 64 -472 80 -438
rect -240 -540 -206 -478
rect 206 -540 240 -478
rect -240 -574 -144 -540
rect 144 -574 240 -540
<< viali >>
rect -64 438 64 472
rect -126 -388 -92 388
rect 92 -388 126 388
rect -64 -472 64 -438
<< metal1 >>
rect -76 472 76 478
rect -76 438 -64 472
rect 64 438 76 472
rect -76 432 76 438
rect -132 388 -86 400
rect -132 -388 -126 388
rect -92 -388 -86 388
rect -132 -400 -86 -388
rect 86 388 132 400
rect 86 -388 92 388
rect 126 -388 132 388
rect 86 -400 132 -388
rect -76 -438 76 -432
rect -76 -472 -64 -438
rect 64 -472 76 -438
rect -76 -478 76 -472
<< labels >>
rlabel psubdiffcont 0 -557 0 -557 0 B
port 1 nsew
rlabel ndiffc -109 0 -109 0 0 D
port 2 nsew
rlabel ndiffc 109 0 109 0 0 S
port 3 nsew
rlabel polycont 0 455 0 455 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -223 -557 223 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
