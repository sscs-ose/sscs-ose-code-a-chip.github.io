.subckt avsd_cmp vcc gnd en vout inn inp net4

XM2 VDIFF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 
XM1 net1 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 
XM12 VOUT2 VOUT1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
XM10 VOUT1 VDIFF VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=6 

XM16 VOUT VOUT2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
XM22 VOUT2 EN VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
XM20 VOUT VOUT2 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 
XM17 net5 EN GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 
XM13 VOUT2 VOUT1 net5 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 
XM11 VOUT1 VCC GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 
XM7 net3 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 
XM18 net4 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 
XM6 net1 VOUT2 net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 
XM8 VDIFF VOUT1 net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 
XM5 net2 VCC GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 
XM3 net1 INN net2 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 
XM4 VDIFF INP net2 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 

xR1 vdd ref gnd sky130_fd_pr__res_high_po_0p69 l=100

.ends
