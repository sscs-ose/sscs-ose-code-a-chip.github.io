* SKY130 Spice File.
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope=2.0e-3
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope=0.0255
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope1=2.0e-3
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope1=0.028
