** sch_path: /foss/designs/clockdiv_try.sch
**.subckt clockdiv_try
Vinp4 net72 net68 DC 1.5 PWL(0 -0.5u 0.008 5.85u 0.016 5.06u 0.024 -4.9u 0.032 -4.6u 0.04 6.71u 0.048 11.2u 0.056 -1.3u 0.064
+ -10.4u 0.072 -27.5u 0.08 -24.0u 0.088 -22.5u 0.096 -16.1u 0.104 -12.5u 0.112 -16.1u 0.12 -12.5u 0.128 -7.8u 0.136 -12.6u 0.144 -0.9u
+ 0.152 20.7u 0.16 20.7u 0.168 34.7u 0.176 23.7u 0.184 20.7u 0.192 23.7u 0.2 20.7u 0.208 35.3u 0.216 24.6u 0.224 8.00u 0.232 8u 0.24
+ 6.43u 0.248 -0.2u 0.256 -4.5u 0.264 -1.7u 0.272 -1.6u 0.28 -6.5u 0.288 -11.6u 0.296 -14.5u 0.304 -6.3u 0.312 -14.5u 0.32 -6.3u 0.328
+ -0.8u 0.336 6.53u 0.344 3.69u 0.352 -12.4u 0.36 -17.6u 0.368 -10.4u 0.376 -9.5u 0.384 -6.9u 0.392 -9.5u 0.4 -6.9u)
R1 net72 Vin1p 50k m=1
Vinn4 net68 GND 1.0
R2 net68 Vin1n 50k m=1
Vinp5 net73 net69 DC 1.5 PWL(0 1.30u 0.008 3.10u 0.016 0.21u 0.024 -14.u 0.032 -8.9u 0.04 2.00u 0.048 10.0u 0.056 -0.3u 0.064
+ -27.9u 0.072 -36.3u 0.08 -34.7u 0.088 -41.3u 0.096 -27.6u 0.104 -16.1u 0.112 -27.6u 0.12 -16.1u 0.128 -5.7u 0.136 -2.6u 0.144 9.37u
+ 0.152 36.5u 0.16 48.6u 0.168 50.1u 0.176 32.8u 0.184 30.5u 0.192 32.8u 0.2 30.5u 0.208 32.3u 0.216 20.9u 0.224 18.7u 0.232 18.7u 0.24
+ 15.3u 0.248 3.39u 0.256 3.14u 0.264 1.34u 0.272 -2.8u 0.28 -9.9u 0.288 -17.0u 0.296 -20.0u 0.304 -17.3u 0.312 -20.0u 0.32 -17.3u 0.328
+ -2.6u 0.336 -4.5u 0.344 -6.4u 0.352 -17.3u 0.36 -35.2u 0.368 -32.8u 0.376 -32.1u 0.384 -34.7u 0.392 -32.1u 0.4 -34.7u)
R7 net73 Vin2p 50k m=1
Vinn5 net69 GND 1.0
R12 net69 Vin2n 50k m=1
Vinp6 net74 net70 DC 1.5 PWL(0 -1.2u 0.008 2.51u 0.016 1.86u 0.024 -9.7u 0.032 -5.4u 0.04 -0.8u 0.048 5.06u 0.056 2.51u 0.064
+ -15.4u 0.072 -19.0u 0.08 -18.4u 0.088 -25.4u 0.096 -17.7u 0.104 -11.4u 0.112 17.7u 0.12 -11.4u 0.128 -5.98u 0.136 0.34u 0.144 5.98u
+ 0.152 19.3u 0.16 30.2u 0.168 29.2u 0.176 13.7u 0.184 17.8u 0.192 13.7u 0.2 17.8u 0.208 15.7u 0.216 8.20u 0.224 13.4u 0.232 13.4u 0.24
+ 14.7u 0.248 5.86u 0.256 1.73u 0.264 4.34u 0.272 -3.7u 0.28 -8.3u 0.288 -13.u 0.296 -15.u 0.304 -9.2u 0.312 -15.4u 0.32 -9.2u 0.328
+ 1.98u 0.336 -2.9u 0.344 -2.6u 0.352 -9.7u 0.36 -27.4u 0.368 -29.0u 0.376 -23.9u 0.384 -28.1u 0.392 -23.9u 0.4 -28.1u)
R13 net74 Vin3p 50k m=1
Vinn6 net70 GND 1.0
R14 net70 Vin3n 50k m=1
Vinp7 net75 net71 DC 1.5 PWL(0 -5.2u 0.008 -2.1u 0.016 4.16u 0.024 -7.5u 0.032 -5.6u 0.04 -1.2u 0.048 4.29u 0.056 5.27u 0.064
+ -12.0u 0.072 -16.4u 0.08 -14.9u 0.088 -22.7u 0.096 -11.1u 0.104 -2.1u 0.112 -11.1u 0.12 -2.1u 0.128 -1.2u 0.136 8.03u 0.144 7.09u 0.152
+ 14.1u 0.16 23.2u 0.168 20.9u 0.176 11.2u 0.184 12.6u 0.192 11.2u 0.2 12.6u 0.208 7.04u 0.216 -2.2u 0.224 8.14u 0.232 8.14u 0.24 13.9u
+ 0.248 0.46u 0.256 0.23u 0.264 4.14u 0.272 -3.7u 0.28 -5.4u 0.288 -10.1u 0.296 -10.5u 0.304 -5.9u 0.312 -10.5u 0.32 -5.9u 0.328 0.59u
+ 0.336 -2.7u 0.344 -3.02u 0.352 -8.3u 0.36 -29.9u 0.368 -33.6u 0.376 -23.0u 0.384 -24.1u 0.392 -23.0u 0.4 -24.1u)
R15 net75 Vin4p 50k m=1
Vinn7 net71 GND 1.0
R16 net71 Vin4n 50k m=1
VDD net77 GND DC 3.3
R3 net77 net4 150m m=1
Vclkin net78 GND PULSE(0 3.3 0 10n 10n 0.5m 1m)
R4 net78 net5 50 m=1
VDD1 net79 GND DC 3.3
R5 net79 VDD 150m m=1
Vclkin1 net80 GND PULSE(0 3.3 0 10n 10n 125u 250u)
R6 net80 net1 50 m=1
VDD2 net81 GND DC 3.3
R8 net81 net3 150m m=1
Vclkin2 net82 GND PULSE(0 3.3 0 10n 10n 250u 500u)
R9 net82 net2 50 m=1
* noconn _CLKA
* noconn CLKA
* noconn _CLKB
* noconn CLKB
* noconn _CLKC
* noconn CLKC
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn VDD
* noconn VDD
* noconn VDD
* noconn _CLKB
* noconn CLKB
* noconn VDD
* noconn _CLKB
* noconn CLKB
* noconn VDD
* noconn VDD
* noconn _CLKC
* noconn CLKC
* noconn VDD
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn _CLKA
* noconn CLKA
* noconn VDD
* noconn VDD
* noconn VDD
* noconn _CLKB
* noconn CLKB
* noconn VDD
* noconn _CLKB
* noconn CLKB
* noconn VDD
* noconn VDD
* noconn _CLKC
* noconn CLKC
* noconn VDD
V19 net59 GND 1.5
V20 net60 GND 3.3
R10 net60 VDD 150m m=1
R11 net59 VBIAS 150m m=1
V2 net61 GND 1
R17 net61 VCM 150m m=1
* noconn VDD
* noconn VBIAS
* noconn VCM
* noconn VDD
* noconn OUTCH1PFIN
* noconn OUTCH1NFIN
* noconn OUTCH2PFIN
* noconn OUTCH2NFIN
* noconn OUTCH3PFIN
* noconn OUTCH3NFIN
* noconn OUTCH4PFIN
* noconn OUTCH4NFIN
* noconn VDD
* noconn VDD
* noconn VDD
* noconn VDD
x24 VDD VBIAS net51 net62 net52 net76 net45 net53 net46 net54 net55 net47 net48 net56 net57 net49 net50 net58 GND VCM FULL_INA_TB
x25 _CLKA CLKA Vin1p net6 net7 Vin1n VDD GND switch_A
x1 _CLKA CLKA Vin2p net8 net9 Vin2n VDD GND switch_A
x2 _CLKA CLKA Vin3p net10 net11 Vin3n VDD GND switch_A
x3 _CLKA CLKA Vin4p net12 net13 Vin4n VDD GND switch_A
x4 _CLKA CLKA net37 net22 net63 net38 VDD GND switch_A
x5 _CLKA CLKA net39 net23 net24 net40 VDD GND switch_A
x6 _CLKA CLKA net41 net25 net26 net42 VDD GND switch_A
x7 _CLKA CLKA net43 net27 net28 net44 VDD GND switch_A
x8 _CLKB CLKB net7 net14 net16 net9 net15 net6 net17 net8 GND VDD switch_B
x9 _CLKB CLKB net11 net18 net20 net13 net19 net10 net21 net12 GND VDD switch_B
x10 _CLKB CLKB net29 net37 net39 net31 net38 net30 net40 net32 GND VDD switch_B
x11 _CLKB CLKB net33 net41 net43 net35 net42 net34 net44 net36 GND VDD switch_B
x12 CLKC _CLKC net62 net14 net18 net47 net45 net16 net49 net20 net76 net15 net48 net19 net17 net46 net50 net21 GND VDD switch_C
x13 CLKC _CLKC net29 net51 net55 net33 net31 net53 net35 net57 net30 net52 net34 net56 net54 net32 net36 net58 GND VDD switch_C
x14 net64 net67 GND net63 OUTCH1NFIN VDD net66 net65 OUTCH1PFIN net22 lpf
x15 net64 net67 GND net24 OUTCH2NFIN VDD net66 net65 OUTCH2PFIN net23 lpf
x16 net64 net67 GND net26 OUTCH3NFIN VDD net66 net65 OUTCH3PFIN net25 lpf
x17 net64 net67 GND net28 OUTCH4NFIN VDD net66 net65 OUTCH4PFIN net27 lpf
x18 VDD net64 net65 GND net1 net66 net67 clk_lpf
x19 VDD _CLKA GND net1 CLKA clk
x20 net3 _CLKB GND net2 CLKB clk
x21 net4 _CLKC GND net5 CLKC clk
**** begin user architecture code


.tran 100u 0.4 0 100u
.options method=gear
.options plotwinsize=0
.control
run
plot v(OUTCH1PFIN)-V(OUTCH1NFIN) v(OUTCH2PFIN)-V(OUTCH2NFIN) v(OUTCH3PFIN)-V(OUTCH3NFIN) v(OUTCH4PFIN)-V(OUTCH4NFIN)
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical
* .lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_statistical

**** end user architecture code
**.ends

* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/INA/FULL_INA_TB.sym # of pins=40
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/INA/FULL_INA_TB.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/INA/FULL_INA_TB.sch
.subckt FULL_INA_TB VDD VBIAS ch1_out+ ch1_in+ ch1_out- ch1_in- ch2_in+ ch2_out+ ch2_in- ch2_out- ch3_out+ ch3_in+ ch3_in-
+ ch3_out- ch4_out+ ch4_in+ ch4_in- ch4_out- VSS VCM
*.opin ch1_out-
*.opin ch1_out+
*.ipin ch1_in+
*.ipin ch1_in-
*.iopin VCM
*.iopin VBIAS
*.iopin VDD
*.opin ch2_out-
*.ipin ch2_in+
*.ipin ch2_in-
*.opin ch3_out+
*.ipin ch3_in+
*.ipin ch3_in-
*.opin ch4_out-
*.opin ch4_out+
*.ipin ch4_in+
*.ipin ch4_in-
*.iopin VSS
*.opin ch3_out-
*.opin ch2_out+
x1 VCM VDD VBIAS ch1_out- ch1_out+ ch1_in+ ch1_in- VSS INA_STAGE_FIXED
x2 VCM VDD VBIAS ch2_out- ch2_out+ ch2_in+ ch2_in- VSS INA_STAGE_FIXED
x3 VCM VDD VBIAS ch3_out- ch3_out+ ch3_in+ ch3_in- VSS INA_STAGE_FIXED
x4 VCM VDD VBIAS ch4_out- ch4_out+ ch4_in+ ch4_in- VSS INA_STAGE_FIXED
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_A.sym # of pins=8
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_A.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_A.sch
.subckt switch_A CLK _CLK Vin1 Vout2 Vout1 Vin2 VDD VSS
*.ipin Vin1
*.opin Vout2
*.ipin Vin2
*.opin Vout1
*.ipin CLK
*.ipin _CLK
*.ipin VDD
*.ipin VSS
XM1 Vout1 CLK Vin1 VSS nfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 Vout1 _CLK Vin1 VDD pfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 Vout2 _CLK Vin1 VSS nfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 Vout2 CLK Vin1 VDD pfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 Vin2 CLK Vout2 VSS nfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 Vin2 _CLK Vout2 VDD pfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 Vin2 _CLK Vout1 VSS nfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 Vin2 CLK Vout1 VDD pfet_03v3 L=0.5u W=15u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_B.sym # of pins=12
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_B.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_B.sch
.subckt switch_B CLK _CLK Vin1p Vout1p Vout2p Vin2p Vout1n Vin1n Vout2n Vin2n VSS VDD
*.ipin Vin1p
*.ipin Vin2p
*.ipin Vin1n
*.ipin Vin2n
*.opin Vout1p
*.opin Vout2p
*.opin Vout1n
*.opin Vout2n
*.ipin CLK
*.ipin _CLK
*.ipin VDD
*.ipin VSS
x1 CLK _CLK Vin1p Vout2p Vout1p Vin2p VDD VSS switch_A
x2 CLK _CLK Vin1n Vout2n Vout1n Vin2n VDD VSS switch_A
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_C.sym # of pins=20
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_C.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/switch_C.sch
.subckt switch_C CLK _CLK Vout1p Vin1p Vin3p Vout3p Vout2p Vin2p Vout4p Vin4p Vout1n Vin1n Vout3n Vin3n Vin2n Vout2n Vout4n Vin4n
+ VSS VDD
*.ipin Vin1p
*.ipin Vin2p
*.opin Vout1p
*.opin Vout2p
*.ipin Vin4n
*.opin Vout4n
*.ipin Vin2n
*.opin Vout2n
*.ipin Vin3n
*.opin Vout3n
*.ipin Vin1n
*.opin Vout1n
*.ipin Vin4p
*.opin Vout4p
*.ipin Vin3p
*.opin Vout3p
*.ipin CLK
*.ipin _CLK
*.ipin VDD
*.ipin VSS
x1 CLK _CLK Vin1p Vout1p Vout3p Vin3p VDD VSS switch_A
x2 CLK _CLK Vin2p Vout2p Vout4p Vin4p VDD VSS switch_A
x3 CLK _CLK Vin1n Vout1n Vout3n Vin3n VDD VSS switch_A
x4 CLK _CLK Vin2n Vout2n Vout4n Vin4n VDD VSS switch_A
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/LPF/lpf.sym # of pins=10
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/LPF/lpf.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/LPF/lpf.sch
.subckt lpf _CLK CLK1 VSS Vin1 Vout1 VDD CLK _CLK1 Vout2 Vin2
*.ipin VSS
*.ipin VDD
*.ipin _CLK
*.ipin CLK
*.ipin Vin1
*.ipin Vin2
*.ipin CLK1
*.ipin _CLK1
*.opin Vout1
*.opin Vout2
XM3 net1 _CLK Vin1 VSS nfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net1 CLK Vin1 VDD pfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 Vin2 _CLK net2 VSS nfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 Vin2 CLK net2 VDD pfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM19 Vout1 CLK1 net1 VSS nfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM20 Vout1 _CLK1 net1 VDD pfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM23 net2 CLK1 Vout2 VSS nfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM24 net2 _CLK1 Vout2 VDD pfet_03v3 L=0.3u W=5u nf=3 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XC1 net1 net2 cap_mim_2f0fF c_width=10e-6 c_length=10e-6 m=3
XC2 net1 net2 cap_mim_2f0fF c_width=10e-6 c_length=10e-6 m=3
XC3 Vout1 Vout2 cap_mim_2f0fF c_width=10e-6 c_length=10e-6 m=3
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/LPF/Complementary Clk for LPF/clk_lpf.sym # of pins=7
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/LPF/Complementary Clk for LPF/clk_lpf.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/LPF/Complementary Clk for LPF/clk_lpf.sch
.subckt clk_lpf VDD _CLK _CLK1 VSS CLK_IN CLK CLK1
*.opin _CLK1
*.ipin CLK_IN
*.opin CLK1
*.ipin VDD
*.ipin VSS
*.opin _CLK
*.opin CLK
XM9 net1 VDD CLK_IN VSS nfet_03v3 L=0.5u W=3u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM10 CLK_IN VSS net1 VDD pfet_03v3 L=0.5u W=3u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM11 _CLK net1 VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM12 _CLK net1 VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM14 net2 CLK_IN VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM15 net2 CLK_IN VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM16 CLK net2 VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM17 CLK net2 VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
* noconn _CLK
* noconn CLK
XM1 net3 CLK VDD VDD pfet_03v3 L=0.5u W=1u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net3 CLK VSS VSS nfet_03v3 L=0.5u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 CLK1 net3 VDD VDD pfet_03v3 L=0.5u W=1u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 CLK1 net3 VSS VSS nfet_03v3 L=0.5u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
* noconn _CLK
XM13 net4 _CLK VDD VDD pfet_03v3 L=0.5u W=1u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM18 net4 _CLK VSS VSS nfet_03v3 L=0.5u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM21 _CLK1 net4 VDD VDD pfet_03v3 L=0.5u W=1u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM22 _CLK1 net4 VSS VSS nfet_03v3 L=0.5u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/Complementary_CLK_CS/clk.sym # of pins=5
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/Complementary_CLK_CS/clk.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/CHOPPER SWITCHES/Complementary_CLK_CS/clk.sch
.subckt clk VDD _CLK VSS CLK_IN CLK
*.opin CLK
*.opin _CLK
*.ipin VSS
*.ipin VDD
*.ipin CLK_IN
XM1 net1 VDD CLK_IN VSS nfet_03v3 L=0.5u W=3u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 CLK_IN VSS net1 VDD pfet_03v3 L=0.5u W=3u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 _CLK net1 VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 _CLK net1 VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net2 CLK_IN VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net2 CLK_IN VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 CLK net2 VDD VDD pfet_03v3 L=0.3u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 CLK net2 VSS VSS nfet_03v3 L=0.3u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  DESIGN_ONLY/FULL_SCH_FILE/INA/INA_STAGE_FIXED.sym # of pins=8
** sym_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/INA/INA_STAGE_FIXED.sym
** sch_path: /foss/designs/DESIGN_ONLY/FULL_SCH_FILE/INA/INA_STAGE_FIXED.sch
.subckt INA_STAGE_FIXED VCM VDD VB out2 out1 in1 in2 VSS
*.opin out1
*.opin out2
*.ipin in1
*.ipin in2
*.iopin VDD
*.iopin VB
*.iopin VSS
*.iopin VCM
XM10 net1 VB VDD VDD pfet_03v3 L=3u W=0.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM11 out1 in1 net1 net1 pfet_03v3 L=3u W=6u nf=6 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM12 out2 in2 net1 net1 pfet_03v3 L=3u W=6u nf=6 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM13 out1 in1 net2 net2 nfet_03v3 L=3u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM14 out2 in2 net2 net2 nfet_03v3 L=3u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM15 net2 out1 VSS VSS nfet_03v3 L=3u W=0.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM16 net2 out2 VSS VSS nfet_03v3 L=3u W=0.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM17 VCM VCM in1 in1 pfet_03v3 L=3u W=0.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM18 VCM VCM in2 in2 pfet_03v3 L=3u W=0.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
