# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_20v0_nvt_withptap_iso
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_20v0_nvt_withptap_iso ;
  ORIGIN  15.29000  9.910000 ;
  SIZE  32.08000 BY  49.82500 ;
  OBS
    LAYER li1 ;
      RECT -15.290000 -9.910000  16.790000 -9.500000 ;
      RECT -15.290000 -9.500000 -14.880000 39.505000 ;
      RECT -15.290000 39.505000  16.790000 39.915000 ;
      RECT  -5.340000  0.045000  -4.670000 29.955000 ;
      RECT  -4.150000  0.045000  -3.480000 29.955000 ;
      RECT  -1.045000 -3.285000   2.775000 -2.215000 ;
      RECT   0.075000  0.215000   1.425000 29.785000 ;
      RECT   4.980000  0.045000   5.650000 29.955000 ;
      RECT   6.170000  0.045000   6.840000 29.955000 ;
      RECT  16.380000 -9.500000  16.790000 39.505000 ;
    LAYER mcon ;
      RECT -15.170000 -9.385000 -15.000000 -9.215000 ;
      RECT -15.170000 -9.025000 -15.000000 -8.855000 ;
      RECT -15.170000 -8.665000 -15.000000 -8.495000 ;
      RECT -15.170000 -8.305000 -15.000000 -8.135000 ;
      RECT -15.170000 -7.945000 -15.000000 -7.775000 ;
      RECT -15.170000 -7.585000 -15.000000 -7.415000 ;
      RECT -15.170000 -7.225000 -15.000000 -7.055000 ;
      RECT -15.170000 -6.865000 -15.000000 -6.695000 ;
      RECT -15.170000 -6.505000 -15.000000 -6.335000 ;
      RECT -15.170000 -6.145000 -15.000000 -5.975000 ;
      RECT -15.170000 -5.785000 -15.000000 -5.615000 ;
      RECT -15.170000 -5.425000 -15.000000 -5.255000 ;
      RECT -15.170000 -5.065000 -15.000000 -4.895000 ;
      RECT -15.170000 -4.705000 -15.000000 -4.535000 ;
      RECT -15.170000 -4.345000 -15.000000 -4.175000 ;
      RECT -15.170000 -3.985000 -15.000000 -3.815000 ;
      RECT -15.170000 -3.625000 -15.000000 -3.455000 ;
      RECT -15.170000 -3.265000 -15.000000 -3.095000 ;
      RECT -15.170000 -2.905000 -15.000000 -2.735000 ;
      RECT -15.170000 -2.545000 -15.000000 -2.375000 ;
      RECT -15.170000 -2.185000 -15.000000 -2.015000 ;
      RECT -15.170000 -1.825000 -15.000000 -1.655000 ;
      RECT -15.170000 -1.465000 -15.000000 -1.295000 ;
      RECT -15.170000 -1.105000 -15.000000 -0.935000 ;
      RECT -15.170000 -0.745000 -15.000000 -0.575000 ;
      RECT -15.170000 -0.385000 -15.000000 -0.215000 ;
      RECT -15.170000 -0.025000 -15.000000  0.145000 ;
      RECT -15.170000  0.335000 -15.000000  0.505000 ;
      RECT -15.170000  0.695000 -15.000000  0.865000 ;
      RECT -15.170000  1.055000 -15.000000  1.225000 ;
      RECT -15.170000  1.415000 -15.000000  1.585000 ;
      RECT -15.170000  1.775000 -15.000000  1.945000 ;
      RECT -15.170000  2.135000 -15.000000  2.305000 ;
      RECT -15.170000  2.495000 -15.000000  2.665000 ;
      RECT -15.170000  2.855000 -15.000000  3.025000 ;
      RECT -15.170000  3.215000 -15.000000  3.385000 ;
      RECT -15.170000  3.575000 -15.000000  3.745000 ;
      RECT -15.170000  3.935000 -15.000000  4.105000 ;
      RECT -15.170000  4.295000 -15.000000  4.465000 ;
      RECT -15.170000  4.655000 -15.000000  4.825000 ;
      RECT -15.170000  5.015000 -15.000000  5.185000 ;
      RECT -15.170000  5.375000 -15.000000  5.545000 ;
      RECT -15.170000  5.735000 -15.000000  5.905000 ;
      RECT -15.170000  6.095000 -15.000000  6.265000 ;
      RECT -15.170000  6.455000 -15.000000  6.625000 ;
      RECT -15.170000  6.815000 -15.000000  6.985000 ;
      RECT -15.170000  7.175000 -15.000000  7.345000 ;
      RECT -15.170000  7.535000 -15.000000  7.705000 ;
      RECT -15.170000  7.895000 -15.000000  8.065000 ;
      RECT -15.170000  8.255000 -15.000000  8.425000 ;
      RECT -15.170000  8.615000 -15.000000  8.785000 ;
      RECT -15.170000  8.975000 -15.000000  9.145000 ;
      RECT -15.170000  9.335000 -15.000000  9.505000 ;
      RECT -15.170000  9.695000 -15.000000  9.865000 ;
      RECT -15.170000 10.055000 -15.000000 10.225000 ;
      RECT -15.170000 10.415000 -15.000000 10.585000 ;
      RECT -15.170000 10.775000 -15.000000 10.945000 ;
      RECT -15.170000 11.135000 -15.000000 11.305000 ;
      RECT -15.170000 11.495000 -15.000000 11.665000 ;
      RECT -15.170000 11.855000 -15.000000 12.025000 ;
      RECT -15.170000 12.215000 -15.000000 12.385000 ;
      RECT -15.170000 12.575000 -15.000000 12.745000 ;
      RECT -15.170000 12.935000 -15.000000 13.105000 ;
      RECT -15.170000 13.295000 -15.000000 13.465000 ;
      RECT -15.170000 13.655000 -15.000000 13.825000 ;
      RECT -15.170000 14.015000 -15.000000 14.185000 ;
      RECT -15.170000 14.375000 -15.000000 14.545000 ;
      RECT -15.170000 14.735000 -15.000000 14.905000 ;
      RECT -15.170000 15.095000 -15.000000 15.265000 ;
      RECT -15.170000 15.455000 -15.000000 15.625000 ;
      RECT -15.170000 15.815000 -15.000000 15.985000 ;
      RECT -15.170000 16.175000 -15.000000 16.345000 ;
      RECT -15.170000 16.535000 -15.000000 16.705000 ;
      RECT -15.170000 16.895000 -15.000000 17.065000 ;
      RECT -15.170000 17.255000 -15.000000 17.425000 ;
      RECT -15.170000 17.615000 -15.000000 17.785000 ;
      RECT -15.170000 17.975000 -15.000000 18.145000 ;
      RECT -15.170000 18.335000 -15.000000 18.505000 ;
      RECT -15.170000 18.695000 -15.000000 18.865000 ;
      RECT -15.170000 19.055000 -15.000000 19.225000 ;
      RECT -15.170000 19.415000 -15.000000 19.585000 ;
      RECT -15.170000 19.775000 -15.000000 19.945000 ;
      RECT -15.170000 20.135000 -15.000000 20.305000 ;
      RECT -15.170000 20.495000 -15.000000 20.665000 ;
      RECT -15.170000 20.855000 -15.000000 21.025000 ;
      RECT -15.170000 21.215000 -15.000000 21.385000 ;
      RECT -15.170000 21.575000 -15.000000 21.745000 ;
      RECT -15.170000 21.935000 -15.000000 22.105000 ;
      RECT -15.170000 22.295000 -15.000000 22.465000 ;
      RECT -15.170000 22.655000 -15.000000 22.825000 ;
      RECT -15.170000 23.015000 -15.000000 23.185000 ;
      RECT -15.170000 23.375000 -15.000000 23.545000 ;
      RECT -15.170000 23.735000 -15.000000 23.905000 ;
      RECT -15.170000 24.095000 -15.000000 24.265000 ;
      RECT -15.170000 24.455000 -15.000000 24.625000 ;
      RECT -15.170000 24.815000 -15.000000 24.985000 ;
      RECT -15.170000 25.175000 -15.000000 25.345000 ;
      RECT -15.170000 25.535000 -15.000000 25.705000 ;
      RECT -15.170000 25.895000 -15.000000 26.065000 ;
      RECT -15.170000 26.255000 -15.000000 26.425000 ;
      RECT -15.170000 26.615000 -15.000000 26.785000 ;
      RECT -15.170000 26.975000 -15.000000 27.145000 ;
      RECT -15.170000 27.335000 -15.000000 27.505000 ;
      RECT -15.170000 27.695000 -15.000000 27.865000 ;
      RECT -15.170000 28.055000 -15.000000 28.225000 ;
      RECT -15.170000 28.415000 -15.000000 28.585000 ;
      RECT -15.170000 28.775000 -15.000000 28.945000 ;
      RECT -15.170000 29.135000 -15.000000 29.305000 ;
      RECT -15.170000 29.495000 -15.000000 29.665000 ;
      RECT -15.170000 29.855000 -15.000000 30.025000 ;
      RECT -15.170000 30.215000 -15.000000 30.385000 ;
      RECT -15.170000 30.575000 -15.000000 30.745000 ;
      RECT -15.170000 30.935000 -15.000000 31.105000 ;
      RECT -15.170000 31.295000 -15.000000 31.465000 ;
      RECT -15.170000 31.655000 -15.000000 31.825000 ;
      RECT -15.170000 32.015000 -15.000000 32.185000 ;
      RECT -15.170000 32.375000 -15.000000 32.545000 ;
      RECT -15.170000 32.735000 -15.000000 32.905000 ;
      RECT -15.170000 33.095000 -15.000000 33.265000 ;
      RECT -15.170000 33.455000 -15.000000 33.625000 ;
      RECT -15.170000 33.815000 -15.000000 33.985000 ;
      RECT -15.170000 34.175000 -15.000000 34.345000 ;
      RECT -15.170000 34.535000 -15.000000 34.705000 ;
      RECT -15.170000 34.895000 -15.000000 35.065000 ;
      RECT -15.170000 35.255000 -15.000000 35.425000 ;
      RECT -15.170000 35.615000 -15.000000 35.785000 ;
      RECT -15.170000 35.975000 -15.000000 36.145000 ;
      RECT -15.170000 36.335000 -15.000000 36.505000 ;
      RECT -15.170000 36.695000 -15.000000 36.865000 ;
      RECT -15.170000 37.055000 -15.000000 37.225000 ;
      RECT -15.170000 37.415000 -15.000000 37.585000 ;
      RECT -15.170000 37.775000 -15.000000 37.945000 ;
      RECT -15.170000 38.135000 -15.000000 38.305000 ;
      RECT -15.170000 38.495000 -15.000000 38.665000 ;
      RECT -15.170000 38.855000 -15.000000 39.025000 ;
      RECT -15.170000 39.215000 -15.000000 39.385000 ;
      RECT -14.635000 -9.790000 -14.465000 -9.620000 ;
      RECT -14.635000 39.625000 -14.465000 39.795000 ;
      RECT -14.275000 -9.790000 -14.105000 -9.620000 ;
      RECT -14.275000 39.625000 -14.105000 39.795000 ;
      RECT -13.915000 -9.790000 -13.745000 -9.620000 ;
      RECT -13.915000 39.625000 -13.745000 39.795000 ;
      RECT -13.555000 -9.790000 -13.385000 -9.620000 ;
      RECT -13.555000 39.625000 -13.385000 39.795000 ;
      RECT -13.195000 -9.790000 -13.025000 -9.620000 ;
      RECT -13.195000 39.625000 -13.025000 39.795000 ;
      RECT -12.835000 -9.790000 -12.665000 -9.620000 ;
      RECT -12.835000 39.625000 -12.665000 39.795000 ;
      RECT -12.475000 -9.790000 -12.305000 -9.620000 ;
      RECT -12.475000 39.625000 -12.305000 39.795000 ;
      RECT -12.115000 -9.790000 -11.945000 -9.620000 ;
      RECT -12.115000 39.625000 -11.945000 39.795000 ;
      RECT -11.755000 -9.790000 -11.585000 -9.620000 ;
      RECT -11.755000 39.625000 -11.585000 39.795000 ;
      RECT -11.395000 -9.790000 -11.225000 -9.620000 ;
      RECT -11.395000 39.625000 -11.225000 39.795000 ;
      RECT -11.035000 -9.790000 -10.865000 -9.620000 ;
      RECT -11.035000 39.625000 -10.865000 39.795000 ;
      RECT -10.675000 -9.790000 -10.505000 -9.620000 ;
      RECT -10.675000 39.625000 -10.505000 39.795000 ;
      RECT -10.315000 -9.790000 -10.145000 -9.620000 ;
      RECT -10.315000 39.625000 -10.145000 39.795000 ;
      RECT  -9.955000 -9.790000  -9.785000 -9.620000 ;
      RECT  -9.955000 39.625000  -9.785000 39.795000 ;
      RECT  -9.595000 -9.790000  -9.425000 -9.620000 ;
      RECT  -9.595000 39.625000  -9.425000 39.795000 ;
      RECT  -9.235000 -9.790000  -9.065000 -9.620000 ;
      RECT  -9.235000 39.625000  -9.065000 39.795000 ;
      RECT  -8.875000 -9.790000  -8.705000 -9.620000 ;
      RECT  -8.875000 39.625000  -8.705000 39.795000 ;
      RECT  -8.515000 -9.790000  -8.345000 -9.620000 ;
      RECT  -8.515000 39.625000  -8.345000 39.795000 ;
      RECT  -8.155000 -9.790000  -7.985000 -9.620000 ;
      RECT  -8.155000 39.625000  -7.985000 39.795000 ;
      RECT  -7.795000 -9.790000  -7.625000 -9.620000 ;
      RECT  -7.795000 39.625000  -7.625000 39.795000 ;
      RECT  -7.435000 -9.790000  -7.265000 -9.620000 ;
      RECT  -7.435000 39.625000  -7.265000 39.795000 ;
      RECT  -7.075000 -9.790000  -6.905000 -9.620000 ;
      RECT  -7.075000 39.625000  -6.905000 39.795000 ;
      RECT  -6.715000 -9.790000  -6.545000 -9.620000 ;
      RECT  -6.715000 39.625000  -6.545000 39.795000 ;
      RECT  -6.355000 -9.790000  -6.185000 -9.620000 ;
      RECT  -6.355000 39.625000  -6.185000 39.795000 ;
      RECT  -5.995000 -9.790000  -5.825000 -9.620000 ;
      RECT  -5.995000 39.625000  -5.825000 39.795000 ;
      RECT  -5.635000 -9.790000  -5.465000 -9.620000 ;
      RECT  -5.635000 39.625000  -5.465000 39.795000 ;
      RECT  -5.275000 -9.790000  -5.105000 -9.620000 ;
      RECT  -5.275000 39.625000  -5.105000 39.795000 ;
      RECT  -5.270000  0.155000  -4.740000 29.845000 ;
      RECT  -4.915000 -9.790000  -4.745000 -9.620000 ;
      RECT  -4.915000 39.625000  -4.745000 39.795000 ;
      RECT  -4.555000 -9.790000  -4.385000 -9.620000 ;
      RECT  -4.555000 39.625000  -4.385000 39.795000 ;
      RECT  -4.195000 -9.790000  -4.025000 -9.620000 ;
      RECT  -4.195000 39.625000  -4.025000 39.795000 ;
      RECT  -4.080000  0.155000  -3.550000 29.845000 ;
      RECT  -3.835000 -9.790000  -3.665000 -9.620000 ;
      RECT  -3.835000 39.625000  -3.665000 39.795000 ;
      RECT  -3.475000 -9.790000  -3.305000 -9.620000 ;
      RECT  -3.475000 39.625000  -3.305000 39.795000 ;
      RECT  -3.115000 -9.790000  -2.945000 -9.620000 ;
      RECT  -3.115000 39.625000  -2.945000 39.795000 ;
      RECT  -2.755000 -9.790000  -2.585000 -9.620000 ;
      RECT  -2.755000 39.625000  -2.585000 39.795000 ;
      RECT  -2.395000 -9.790000  -2.225000 -9.620000 ;
      RECT  -2.395000 39.625000  -2.225000 39.795000 ;
      RECT  -2.035000 -9.790000  -1.865000 -9.620000 ;
      RECT  -2.035000 39.625000  -1.865000 39.795000 ;
      RECT  -1.675000 -9.790000  -1.505000 -9.620000 ;
      RECT  -1.675000 39.625000  -1.505000 39.795000 ;
      RECT  -1.315000 -9.790000  -1.145000 -9.620000 ;
      RECT  -1.315000 39.625000  -1.145000 39.795000 ;
      RECT  -0.955000 -9.790000  -0.785000 -9.620000 ;
      RECT  -0.955000 39.625000  -0.785000 39.795000 ;
      RECT  -0.900000 -3.205000  -0.730000 -3.035000 ;
      RECT  -0.900000 -2.835000  -0.730000 -2.665000 ;
      RECT  -0.900000 -2.465000  -0.730000 -2.295000 ;
      RECT  -0.595000 -9.790000  -0.425000 -9.620000 ;
      RECT  -0.595000 39.625000  -0.425000 39.795000 ;
      RECT  -0.530000 -3.205000  -0.360000 -3.035000 ;
      RECT  -0.530000 -2.835000  -0.360000 -2.665000 ;
      RECT  -0.530000 -2.465000  -0.360000 -2.295000 ;
      RECT  -0.235000 -9.790000  -0.065000 -9.620000 ;
      RECT  -0.235000 39.625000  -0.065000 39.795000 ;
      RECT  -0.160000 -3.205000   0.010000 -3.035000 ;
      RECT  -0.160000 -2.835000   0.010000 -2.665000 ;
      RECT  -0.160000 -2.465000   0.010000 -2.295000 ;
      RECT   0.125000 -9.790000   0.295000 -9.620000 ;
      RECT   0.125000  0.335000   1.375000 29.665000 ;
      RECT   0.125000 39.625000   0.295000 39.795000 ;
      RECT   0.210000 -3.205000   0.380000 -3.035000 ;
      RECT   0.210000 -2.835000   0.380000 -2.665000 ;
      RECT   0.210000 -2.465000   0.380000 -2.295000 ;
      RECT   0.485000 -9.790000   0.655000 -9.620000 ;
      RECT   0.485000 39.625000   0.655000 39.795000 ;
      RECT   0.580000 -3.205000   0.750000 -3.035000 ;
      RECT   0.580000 -2.835000   0.750000 -2.665000 ;
      RECT   0.580000 -2.465000   0.750000 -2.295000 ;
      RECT   0.845000 -9.790000   1.015000 -9.620000 ;
      RECT   0.845000 39.625000   1.015000 39.795000 ;
      RECT   0.950000 -3.205000   1.120000 -3.035000 ;
      RECT   0.950000 -2.835000   1.120000 -2.665000 ;
      RECT   0.950000 -2.465000   1.120000 -2.295000 ;
      RECT   1.205000 -9.790000   1.375000 -9.620000 ;
      RECT   1.205000 39.625000   1.375000 39.795000 ;
      RECT   1.320000 -3.205000   1.490000 -3.035000 ;
      RECT   1.320000 -2.835000   1.490000 -2.665000 ;
      RECT   1.320000 -2.465000   1.490000 -2.295000 ;
      RECT   1.565000 -9.790000   1.735000 -9.620000 ;
      RECT   1.565000 39.625000   1.735000 39.795000 ;
      RECT   1.690000 -3.205000   1.860000 -3.035000 ;
      RECT   1.690000 -2.835000   1.860000 -2.665000 ;
      RECT   1.690000 -2.465000   1.860000 -2.295000 ;
      RECT   1.925000 -9.790000   2.095000 -9.620000 ;
      RECT   1.925000 39.625000   2.095000 39.795000 ;
      RECT   2.060000 -3.205000   2.230000 -3.035000 ;
      RECT   2.060000 -2.835000   2.230000 -2.665000 ;
      RECT   2.060000 -2.465000   2.230000 -2.295000 ;
      RECT   2.285000 -9.790000   2.455000 -9.620000 ;
      RECT   2.285000 39.625000   2.455000 39.795000 ;
      RECT   2.430000 -3.205000   2.600000 -3.035000 ;
      RECT   2.430000 -2.835000   2.600000 -2.665000 ;
      RECT   2.430000 -2.465000   2.600000 -2.295000 ;
      RECT   2.645000 -9.790000   2.815000 -9.620000 ;
      RECT   2.645000 39.625000   2.815000 39.795000 ;
      RECT   3.005000 -9.790000   3.175000 -9.620000 ;
      RECT   3.005000 39.625000   3.175000 39.795000 ;
      RECT   3.365000 -9.790000   3.535000 -9.620000 ;
      RECT   3.365000 39.625000   3.535000 39.795000 ;
      RECT   3.725000 -9.790000   3.895000 -9.620000 ;
      RECT   3.725000 39.625000   3.895000 39.795000 ;
      RECT   4.085000 -9.790000   4.255000 -9.620000 ;
      RECT   4.085000 39.625000   4.255000 39.795000 ;
      RECT   4.445000 -9.790000   4.615000 -9.620000 ;
      RECT   4.445000 39.625000   4.615000 39.795000 ;
      RECT   4.805000 -9.790000   4.975000 -9.620000 ;
      RECT   4.805000 39.625000   4.975000 39.795000 ;
      RECT   5.050000  0.155000   5.580000 29.845000 ;
      RECT   5.165000 -9.790000   5.335000 -9.620000 ;
      RECT   5.165000 39.625000   5.335000 39.795000 ;
      RECT   5.525000 -9.790000   5.695000 -9.620000 ;
      RECT   5.525000 39.625000   5.695000 39.795000 ;
      RECT   5.885000 -9.790000   6.055000 -9.620000 ;
      RECT   5.885000 39.625000   6.055000 39.795000 ;
      RECT   6.240000  0.155000   6.770000 29.845000 ;
      RECT   6.245000 -9.790000   6.415000 -9.620000 ;
      RECT   6.245000 39.625000   6.415000 39.795000 ;
      RECT   6.605000 -9.790000   6.775000 -9.620000 ;
      RECT   6.605000 39.625000   6.775000 39.795000 ;
      RECT   6.965000 -9.790000   7.135000 -9.620000 ;
      RECT   6.965000 39.625000   7.135000 39.795000 ;
      RECT   7.325000 -9.790000   7.495000 -9.620000 ;
      RECT   7.325000 39.625000   7.495000 39.795000 ;
      RECT   7.685000 -9.790000   7.855000 -9.620000 ;
      RECT   7.685000 39.625000   7.855000 39.795000 ;
      RECT   8.045000 -9.790000   8.215000 -9.620000 ;
      RECT   8.045000 39.625000   8.215000 39.795000 ;
      RECT   8.405000 -9.790000   8.575000 -9.620000 ;
      RECT   8.405000 39.625000   8.575000 39.795000 ;
      RECT   8.765000 -9.790000   8.935000 -9.620000 ;
      RECT   8.765000 39.625000   8.935000 39.795000 ;
      RECT   9.125000 -9.790000   9.295000 -9.620000 ;
      RECT   9.125000 39.625000   9.295000 39.795000 ;
      RECT   9.485000 -9.790000   9.655000 -9.620000 ;
      RECT   9.485000 39.625000   9.655000 39.795000 ;
      RECT   9.845000 -9.790000  10.015000 -9.620000 ;
      RECT   9.845000 39.625000  10.015000 39.795000 ;
      RECT  10.205000 -9.790000  10.375000 -9.620000 ;
      RECT  10.205000 39.625000  10.375000 39.795000 ;
      RECT  10.565000 -9.790000  10.735000 -9.620000 ;
      RECT  10.565000 39.625000  10.735000 39.795000 ;
      RECT  10.925000 -9.790000  11.095000 -9.620000 ;
      RECT  10.925000 39.625000  11.095000 39.795000 ;
      RECT  11.285000 -9.790000  11.455000 -9.620000 ;
      RECT  11.285000 39.625000  11.455000 39.795000 ;
      RECT  11.645000 -9.790000  11.815000 -9.620000 ;
      RECT  11.645000 39.625000  11.815000 39.795000 ;
      RECT  12.005000 -9.790000  12.175000 -9.620000 ;
      RECT  12.005000 39.625000  12.175000 39.795000 ;
      RECT  12.365000 -9.790000  12.535000 -9.620000 ;
      RECT  12.365000 39.625000  12.535000 39.795000 ;
      RECT  12.725000 -9.790000  12.895000 -9.620000 ;
      RECT  12.725000 39.625000  12.895000 39.795000 ;
      RECT  13.085000 -9.790000  13.255000 -9.620000 ;
      RECT  13.085000 39.625000  13.255000 39.795000 ;
      RECT  13.445000 -9.790000  13.615000 -9.620000 ;
      RECT  13.445000 39.625000  13.615000 39.795000 ;
      RECT  13.805000 -9.790000  13.975000 -9.620000 ;
      RECT  13.805000 39.625000  13.975000 39.795000 ;
      RECT  14.165000 -9.790000  14.335000 -9.620000 ;
      RECT  14.165000 39.625000  14.335000 39.795000 ;
      RECT  14.525000 -9.790000  14.695000 -9.620000 ;
      RECT  14.525000 39.625000  14.695000 39.795000 ;
      RECT  14.885000 -9.790000  15.055000 -9.620000 ;
      RECT  14.885000 39.625000  15.055000 39.795000 ;
      RECT  15.245000 -9.790000  15.415000 -9.620000 ;
      RECT  15.245000 39.625000  15.415000 39.795000 ;
      RECT  15.605000 -9.790000  15.775000 -9.620000 ;
      RECT  15.605000 39.625000  15.775000 39.795000 ;
      RECT  15.965000 -9.790000  16.135000 -9.620000 ;
      RECT  15.965000 39.625000  16.135000 39.795000 ;
      RECT  16.500000 -9.385000  16.670000 -9.215000 ;
      RECT  16.500000 -9.025000  16.670000 -8.855000 ;
      RECT  16.500000 -8.665000  16.670000 -8.495000 ;
      RECT  16.500000 -8.305000  16.670000 -8.135000 ;
      RECT  16.500000 -7.945000  16.670000 -7.775000 ;
      RECT  16.500000 -7.585000  16.670000 -7.415000 ;
      RECT  16.500000 -7.225000  16.670000 -7.055000 ;
      RECT  16.500000 -6.865000  16.670000 -6.695000 ;
      RECT  16.500000 -6.505000  16.670000 -6.335000 ;
      RECT  16.500000 -6.145000  16.670000 -5.975000 ;
      RECT  16.500000 -5.785000  16.670000 -5.615000 ;
      RECT  16.500000 -5.425000  16.670000 -5.255000 ;
      RECT  16.500000 -5.065000  16.670000 -4.895000 ;
      RECT  16.500000 -4.705000  16.670000 -4.535000 ;
      RECT  16.500000 -4.345000  16.670000 -4.175000 ;
      RECT  16.500000 -3.985000  16.670000 -3.815000 ;
      RECT  16.500000 -3.625000  16.670000 -3.455000 ;
      RECT  16.500000 -3.265000  16.670000 -3.095000 ;
      RECT  16.500000 -2.905000  16.670000 -2.735000 ;
      RECT  16.500000 -2.545000  16.670000 -2.375000 ;
      RECT  16.500000 -2.185000  16.670000 -2.015000 ;
      RECT  16.500000 -1.825000  16.670000 -1.655000 ;
      RECT  16.500000 -1.465000  16.670000 -1.295000 ;
      RECT  16.500000 -1.105000  16.670000 -0.935000 ;
      RECT  16.500000 -0.745000  16.670000 -0.575000 ;
      RECT  16.500000 -0.385000  16.670000 -0.215000 ;
      RECT  16.500000 -0.025000  16.670000  0.145000 ;
      RECT  16.500000  0.335000  16.670000  0.505000 ;
      RECT  16.500000  0.695000  16.670000  0.865000 ;
      RECT  16.500000  1.055000  16.670000  1.225000 ;
      RECT  16.500000  1.415000  16.670000  1.585000 ;
      RECT  16.500000  1.775000  16.670000  1.945000 ;
      RECT  16.500000  2.135000  16.670000  2.305000 ;
      RECT  16.500000  2.495000  16.670000  2.665000 ;
      RECT  16.500000  2.855000  16.670000  3.025000 ;
      RECT  16.500000  3.215000  16.670000  3.385000 ;
      RECT  16.500000  3.575000  16.670000  3.745000 ;
      RECT  16.500000  3.935000  16.670000  4.105000 ;
      RECT  16.500000  4.295000  16.670000  4.465000 ;
      RECT  16.500000  4.655000  16.670000  4.825000 ;
      RECT  16.500000  5.015000  16.670000  5.185000 ;
      RECT  16.500000  5.375000  16.670000  5.545000 ;
      RECT  16.500000  5.735000  16.670000  5.905000 ;
      RECT  16.500000  6.095000  16.670000  6.265000 ;
      RECT  16.500000  6.455000  16.670000  6.625000 ;
      RECT  16.500000  6.815000  16.670000  6.985000 ;
      RECT  16.500000  7.175000  16.670000  7.345000 ;
      RECT  16.500000  7.535000  16.670000  7.705000 ;
      RECT  16.500000  7.895000  16.670000  8.065000 ;
      RECT  16.500000  8.255000  16.670000  8.425000 ;
      RECT  16.500000  8.615000  16.670000  8.785000 ;
      RECT  16.500000  8.975000  16.670000  9.145000 ;
      RECT  16.500000  9.335000  16.670000  9.505000 ;
      RECT  16.500000  9.695000  16.670000  9.865000 ;
      RECT  16.500000 10.055000  16.670000 10.225000 ;
      RECT  16.500000 10.415000  16.670000 10.585000 ;
      RECT  16.500000 10.775000  16.670000 10.945000 ;
      RECT  16.500000 11.135000  16.670000 11.305000 ;
      RECT  16.500000 11.495000  16.670000 11.665000 ;
      RECT  16.500000 11.855000  16.670000 12.025000 ;
      RECT  16.500000 12.215000  16.670000 12.385000 ;
      RECT  16.500000 12.575000  16.670000 12.745000 ;
      RECT  16.500000 12.935000  16.670000 13.105000 ;
      RECT  16.500000 13.295000  16.670000 13.465000 ;
      RECT  16.500000 13.655000  16.670000 13.825000 ;
      RECT  16.500000 14.015000  16.670000 14.185000 ;
      RECT  16.500000 14.375000  16.670000 14.545000 ;
      RECT  16.500000 14.735000  16.670000 14.905000 ;
      RECT  16.500000 15.095000  16.670000 15.265000 ;
      RECT  16.500000 15.455000  16.670000 15.625000 ;
      RECT  16.500000 15.815000  16.670000 15.985000 ;
      RECT  16.500000 16.175000  16.670000 16.345000 ;
      RECT  16.500000 16.535000  16.670000 16.705000 ;
      RECT  16.500000 16.895000  16.670000 17.065000 ;
      RECT  16.500000 17.255000  16.670000 17.425000 ;
      RECT  16.500000 17.615000  16.670000 17.785000 ;
      RECT  16.500000 17.975000  16.670000 18.145000 ;
      RECT  16.500000 18.335000  16.670000 18.505000 ;
      RECT  16.500000 18.695000  16.670000 18.865000 ;
      RECT  16.500000 19.055000  16.670000 19.225000 ;
      RECT  16.500000 19.415000  16.670000 19.585000 ;
      RECT  16.500000 19.775000  16.670000 19.945000 ;
      RECT  16.500000 20.135000  16.670000 20.305000 ;
      RECT  16.500000 20.495000  16.670000 20.665000 ;
      RECT  16.500000 20.855000  16.670000 21.025000 ;
      RECT  16.500000 21.215000  16.670000 21.385000 ;
      RECT  16.500000 21.575000  16.670000 21.745000 ;
      RECT  16.500000 21.935000  16.670000 22.105000 ;
      RECT  16.500000 22.295000  16.670000 22.465000 ;
      RECT  16.500000 22.655000  16.670000 22.825000 ;
      RECT  16.500000 23.015000  16.670000 23.185000 ;
      RECT  16.500000 23.375000  16.670000 23.545000 ;
      RECT  16.500000 23.735000  16.670000 23.905000 ;
      RECT  16.500000 24.095000  16.670000 24.265000 ;
      RECT  16.500000 24.455000  16.670000 24.625000 ;
      RECT  16.500000 24.815000  16.670000 24.985000 ;
      RECT  16.500000 25.175000  16.670000 25.345000 ;
      RECT  16.500000 25.535000  16.670000 25.705000 ;
      RECT  16.500000 25.895000  16.670000 26.065000 ;
      RECT  16.500000 26.255000  16.670000 26.425000 ;
      RECT  16.500000 26.615000  16.670000 26.785000 ;
      RECT  16.500000 26.975000  16.670000 27.145000 ;
      RECT  16.500000 27.335000  16.670000 27.505000 ;
      RECT  16.500000 27.695000  16.670000 27.865000 ;
      RECT  16.500000 28.055000  16.670000 28.225000 ;
      RECT  16.500000 28.415000  16.670000 28.585000 ;
      RECT  16.500000 28.775000  16.670000 28.945000 ;
      RECT  16.500000 29.135000  16.670000 29.305000 ;
      RECT  16.500000 29.495000  16.670000 29.665000 ;
      RECT  16.500000 29.855000  16.670000 30.025000 ;
      RECT  16.500000 30.215000  16.670000 30.385000 ;
      RECT  16.500000 30.575000  16.670000 30.745000 ;
      RECT  16.500000 30.935000  16.670000 31.105000 ;
      RECT  16.500000 31.295000  16.670000 31.465000 ;
      RECT  16.500000 31.655000  16.670000 31.825000 ;
      RECT  16.500000 32.015000  16.670000 32.185000 ;
      RECT  16.500000 32.375000  16.670000 32.545000 ;
      RECT  16.500000 32.735000  16.670000 32.905000 ;
      RECT  16.500000 33.095000  16.670000 33.265000 ;
      RECT  16.500000 33.455000  16.670000 33.625000 ;
      RECT  16.500000 33.815000  16.670000 33.985000 ;
      RECT  16.500000 34.175000  16.670000 34.345000 ;
      RECT  16.500000 34.535000  16.670000 34.705000 ;
      RECT  16.500000 34.895000  16.670000 35.065000 ;
      RECT  16.500000 35.255000  16.670000 35.425000 ;
      RECT  16.500000 35.615000  16.670000 35.785000 ;
      RECT  16.500000 35.975000  16.670000 36.145000 ;
      RECT  16.500000 36.335000  16.670000 36.505000 ;
      RECT  16.500000 36.695000  16.670000 36.865000 ;
      RECT  16.500000 37.055000  16.670000 37.225000 ;
      RECT  16.500000 37.415000  16.670000 37.585000 ;
      RECT  16.500000 37.775000  16.670000 37.945000 ;
      RECT  16.500000 38.135000  16.670000 38.305000 ;
      RECT  16.500000 38.495000  16.670000 38.665000 ;
      RECT  16.500000 38.855000  16.670000 39.025000 ;
      RECT  16.500000 39.215000  16.670000 39.385000 ;
    LAYER met1 ;
      RECT -15.290000 -9.910000  16.790000 -9.500000 ;
      RECT -15.290000 -9.500000 -14.880000 39.505000 ;
      RECT -15.290000 39.505000  16.790000 39.915000 ;
      RECT  -5.330000  0.095000  -4.680000 29.905000 ;
      RECT  -4.140000  0.095000  -3.490000 29.905000 ;
      RECT  -1.045000 -3.285000   2.775000 -2.215000 ;
      RECT   0.065000  0.275000   1.435000 29.725000 ;
      RECT   4.990000  0.095000   5.640000 29.905000 ;
      RECT   6.180000  0.095000   6.830000 29.905000 ;
      RECT  16.380000 -9.500000  16.790000 39.505000 ;
    LAYER met2 ;
      RECT -1.045000 -3.285000 2.775000 -2.215000 ;
      RECT  0.110000  0.285000 1.390000 29.725000 ;
    LAYER via ;
      RECT -0.945000 -3.250000 -0.685000 -2.990000 ;
      RECT -0.945000 -2.880000 -0.685000 -2.620000 ;
      RECT -0.945000 -2.510000 -0.685000 -2.250000 ;
      RECT -0.575000 -3.250000 -0.315000 -2.990000 ;
      RECT -0.575000 -2.880000 -0.315000 -2.620000 ;
      RECT -0.575000 -2.510000 -0.315000 -2.250000 ;
      RECT -0.205000 -3.250000  0.055000 -2.990000 ;
      RECT -0.205000 -2.880000  0.055000 -2.620000 ;
      RECT -0.205000 -2.510000  0.055000 -2.250000 ;
      RECT  0.140000  0.315000  1.360000 29.695000 ;
      RECT  0.165000 -3.250000  0.425000 -2.990000 ;
      RECT  0.165000 -2.880000  0.425000 -2.620000 ;
      RECT  0.165000 -2.510000  0.425000 -2.250000 ;
      RECT  0.535000 -3.250000  0.795000 -2.990000 ;
      RECT  0.535000 -2.880000  0.795000 -2.620000 ;
      RECT  0.535000 -2.510000  0.795000 -2.250000 ;
      RECT  0.905000 -3.250000  1.165000 -2.990000 ;
      RECT  0.905000 -2.880000  1.165000 -2.620000 ;
      RECT  0.905000 -2.510000  1.165000 -2.250000 ;
      RECT  1.275000 -3.250000  1.535000 -2.990000 ;
      RECT  1.275000 -2.880000  1.535000 -2.620000 ;
      RECT  1.275000 -2.510000  1.535000 -2.250000 ;
      RECT  1.645000 -3.250000  1.905000 -2.990000 ;
      RECT  1.645000 -2.880000  1.905000 -2.620000 ;
      RECT  1.645000 -2.510000  1.905000 -2.250000 ;
      RECT  2.015000 -3.250000  2.275000 -2.990000 ;
      RECT  2.015000 -2.880000  2.275000 -2.620000 ;
      RECT  2.015000 -2.510000  2.275000 -2.250000 ;
      RECT  2.385000 -3.250000  2.645000 -2.990000 ;
      RECT  2.385000 -2.880000  2.645000 -2.620000 ;
      RECT  2.385000 -2.510000  2.645000 -2.250000 ;
  END
END sky130_fd_pr__rf_nfet_20v0_nvt_withptap_iso
END LIBRARY
