# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__pnp_05v5_W3p40L3p40
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pnp_05v5_W3p40L3p40 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  3.720000 BY  3.845000 ;
  OBS
    LAYER li1 ;
      RECT 0.130000 0.130000 3.850000 0.635000 ;
      RECT 0.130000 0.635000 0.635000 3.345000 ;
      RECT 0.130000 3.345000 3.850000 3.850000 ;
      RECT 0.945000 0.945000 3.035000 1.305000 ;
      RECT 0.945000 1.305000 1.305000 2.675000 ;
      RECT 0.945000 2.675000 3.035000 3.035000 ;
      RECT 1.595000 1.595000 2.385000 2.385000 ;
      RECT 2.675000 1.305000 3.035000 2.675000 ;
      RECT 3.345000 0.635000 3.850000 3.345000 ;
    LAYER mcon ;
      RECT 1.665000 1.665000 1.835000 1.835000 ;
      RECT 1.665000 2.145000 1.835000 2.315000 ;
      RECT 2.145000 1.665000 2.315000 1.835000 ;
      RECT 2.145000 2.145000 2.315000 2.315000 ;
    LAYER met1 ;
      RECT 1.575000 1.575000 2.405000 2.405000 ;
  END
END sky130_fd_pr__pnp_05v5_W3p40L3p40
END LIBRARY
