# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o2subcell
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o2subcell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.580000 BY  7.840000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.320000 0.270000 0.460000 ;
      RECT 0.000000 0.460000 8.140000 0.630000 ;
      RECT 0.000000 0.630000 0.270000 1.160000 ;
      RECT 0.000000 1.160000 8.140000 1.330000 ;
      RECT 0.000000 1.330000 0.270000 1.860000 ;
      RECT 0.000000 1.860000 8.140000 2.030000 ;
      RECT 0.000000 2.030000 0.270000 2.560000 ;
      RECT 0.000000 2.560000 8.140000 2.730000 ;
      RECT 0.000000 2.730000 0.270000 3.260000 ;
      RECT 0.000000 3.260000 8.140000 3.430000 ;
      RECT 0.000000 3.430000 0.270000 3.960000 ;
      RECT 0.000000 3.960000 8.140000 4.130000 ;
      RECT 0.000000 4.130000 0.270000 4.660000 ;
      RECT 0.000000 4.660000 8.140000 4.830000 ;
      RECT 0.000000 4.830000 0.270000 5.360000 ;
      RECT 0.000000 5.360000 8.140000 5.530000 ;
      RECT 0.000000 5.530000 0.270000 6.060000 ;
      RECT 0.000000 6.060000 8.140000 6.230000 ;
      RECT 0.000000 6.230000 0.270000 6.760000 ;
      RECT 0.000000 6.760000 8.140000 6.930000 ;
      RECT 0.000000 6.930000 0.270000 7.380000 ;
      RECT 0.440000 0.810000 8.580000 0.980000 ;
      RECT 0.440000 1.510000 8.580000 1.680000 ;
      RECT 0.440000 2.210000 8.580000 2.380000 ;
      RECT 0.440000 2.910000 8.580000 3.080000 ;
      RECT 0.440000 3.610000 8.580000 3.780000 ;
      RECT 0.440000 4.310000 8.580000 4.480000 ;
      RECT 0.440000 5.010000 8.580000 5.180000 ;
      RECT 0.440000 5.710000 8.580000 5.880000 ;
      RECT 0.440000 6.410000 8.580000 6.580000 ;
      RECT 0.440000 7.110000 8.580000 7.280000 ;
      RECT 8.310000 0.460000 8.580000 0.810000 ;
      RECT 8.310000 0.980000 8.580000 1.510000 ;
      RECT 8.310000 1.680000 8.580000 2.210000 ;
      RECT 8.310000 2.380000 8.580000 2.910000 ;
      RECT 8.310000 3.080000 8.580000 3.610000 ;
      RECT 8.310000 3.780000 8.580000 4.310000 ;
      RECT 8.310000 4.480000 8.580000 5.010000 ;
      RECT 8.310000 5.180000 8.580000 5.710000 ;
      RECT 8.310000 5.880000 8.580000 6.410000 ;
      RECT 8.310000 6.580000 8.580000 7.110000 ;
      RECT 8.310000 7.280000 8.580000 7.520000 ;
    LAYER mcon ;
      RECT 0.050000 0.450000 0.220000 0.620000 ;
      RECT 0.050000 0.810000 0.220000 0.980000 ;
      RECT 0.050000 1.170000 0.220000 1.340000 ;
      RECT 0.050000 1.530000 0.220000 1.700000 ;
      RECT 0.050000 1.890000 0.220000 2.060000 ;
      RECT 0.050000 2.250000 0.220000 2.420000 ;
      RECT 0.050000 2.610000 0.220000 2.780000 ;
      RECT 0.050000 2.970000 0.220000 3.140000 ;
      RECT 0.050000 3.330000 0.220000 3.500000 ;
      RECT 0.050000 3.690000 0.220000 3.860000 ;
      RECT 0.050000 4.050000 0.220000 4.220000 ;
      RECT 0.050000 4.410000 0.220000 4.580000 ;
      RECT 0.050000 4.770000 0.220000 4.940000 ;
      RECT 0.050000 5.130000 0.220000 5.300000 ;
      RECT 0.050000 5.490000 0.220000 5.660000 ;
      RECT 0.050000 5.850000 0.220000 6.020000 ;
      RECT 0.050000 6.210000 0.220000 6.380000 ;
      RECT 0.050000 6.570000 0.220000 6.740000 ;
      RECT 0.050000 6.930000 0.220000 7.100000 ;
      RECT 8.360000 0.575000 8.530000 0.745000 ;
      RECT 8.360000 0.935000 8.530000 1.105000 ;
      RECT 8.360000 1.295000 8.530000 1.465000 ;
      RECT 8.360000 1.655000 8.530000 1.825000 ;
      RECT 8.360000 2.015000 8.530000 2.185000 ;
      RECT 8.360000 2.375000 8.530000 2.545000 ;
      RECT 8.360000 2.735000 8.530000 2.905000 ;
      RECT 8.360000 3.095000 8.530000 3.265000 ;
      RECT 8.360000 3.455000 8.530000 3.625000 ;
      RECT 8.360000 3.815000 8.530000 3.985000 ;
      RECT 8.360000 4.175000 8.530000 4.345000 ;
      RECT 8.360000 4.535000 8.530000 4.705000 ;
      RECT 8.360000 4.895000 8.530000 5.065000 ;
      RECT 8.360000 5.255000 8.530000 5.425000 ;
      RECT 8.360000 5.615000 8.530000 5.785000 ;
      RECT 8.360000 5.975000 8.530000 6.145000 ;
      RECT 8.360000 6.335000 8.530000 6.505000 ;
      RECT 8.360000 6.695000 8.530000 6.865000 ;
      RECT 8.360000 7.055000 8.530000 7.225000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 8.580000 0.320000 ;
      RECT 0.000000 0.320000 0.270000 7.380000 ;
      RECT 0.000000 7.520000 8.580000 7.840000 ;
      RECT 0.440000 0.320000 0.580000 7.380000 ;
      RECT 0.720000 0.460000 0.860000 7.520000 ;
      RECT 1.000000 0.320000 1.140000 7.380000 ;
      RECT 1.280000 0.460000 1.420000 7.520000 ;
      RECT 1.560000 0.320000 1.700000 7.380000 ;
      RECT 1.840000 0.460000 1.980000 7.520000 ;
      RECT 2.120000 0.320000 2.260000 7.380000 ;
      RECT 2.400000 0.460000 2.540000 7.520000 ;
      RECT 2.680000 0.320000 2.820000 7.380000 ;
      RECT 2.960000 0.460000 3.100000 7.520000 ;
      RECT 3.240000 0.320000 3.380000 7.380000 ;
      RECT 3.520000 0.460000 3.660000 7.520000 ;
      RECT 3.800000 0.320000 3.940000 7.380000 ;
      RECT 4.080000 0.460000 4.220000 7.520000 ;
      RECT 4.360000 0.320000 4.500000 7.380000 ;
      RECT 4.640000 0.460000 4.780000 7.520000 ;
      RECT 4.920000 0.320000 5.060000 7.380000 ;
      RECT 5.200000 0.460000 5.340000 7.520000 ;
      RECT 5.480000 0.320000 5.620000 7.380000 ;
      RECT 5.760000 0.460000 5.900000 7.520000 ;
      RECT 6.040000 0.320000 6.180000 7.380000 ;
      RECT 6.320000 0.460000 6.460000 7.520000 ;
      RECT 6.600000 0.320000 6.740000 7.380000 ;
      RECT 6.880000 0.460000 7.020000 7.520000 ;
      RECT 7.160000 0.320000 7.300000 7.380000 ;
      RECT 7.440000 0.460000 7.580000 7.520000 ;
      RECT 7.720000 0.320000 7.860000 7.380000 ;
      RECT 8.000000 0.460000 8.140000 7.520000 ;
      RECT 8.310000 0.460000 8.580000 7.520000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 8.580000 0.320000 ;
      RECT 0.000000 0.320000 0.270000 7.380000 ;
      RECT 0.000000 7.520000 8.580000 7.840000 ;
      RECT 0.440000 0.460000 0.580000 7.520000 ;
      RECT 0.720000 0.320000 0.860000 7.380000 ;
      RECT 1.000000 0.460000 1.140000 7.520000 ;
      RECT 1.280000 0.320000 1.420000 7.380000 ;
      RECT 1.560000 0.460000 1.700000 7.520000 ;
      RECT 1.840000 0.320000 1.980000 7.380000 ;
      RECT 2.120000 0.460000 2.260000 7.520000 ;
      RECT 2.400000 0.320000 2.540000 7.380000 ;
      RECT 2.680000 0.460000 2.820000 7.520000 ;
      RECT 2.960000 0.320000 3.100000 7.380000 ;
      RECT 3.240000 0.460000 3.380000 7.520000 ;
      RECT 3.520000 0.320000 3.660000 7.380000 ;
      RECT 3.800000 0.460000 3.940000 7.520000 ;
      RECT 4.080000 0.320000 4.220000 7.380000 ;
      RECT 4.360000 0.460000 4.500000 7.520000 ;
      RECT 4.640000 0.320000 4.780000 7.380000 ;
      RECT 4.920000 0.460000 5.060000 7.520000 ;
      RECT 5.200000 0.320000 5.340000 7.380000 ;
      RECT 5.480000 0.460000 5.620000 7.520000 ;
      RECT 5.760000 0.320000 5.900000 7.380000 ;
      RECT 6.040000 0.460000 6.180000 7.520000 ;
      RECT 6.320000 0.320000 6.460000 7.380000 ;
      RECT 6.600000 0.460000 6.740000 7.520000 ;
      RECT 6.880000 0.320000 7.020000 7.380000 ;
      RECT 7.160000 0.460000 7.300000 7.520000 ;
      RECT 7.440000 0.320000 7.580000 7.380000 ;
      RECT 7.720000 0.460000 7.860000 7.520000 ;
      RECT 8.000000 0.320000 8.140000 7.380000 ;
      RECT 8.310000 0.460000 8.580000 7.520000 ;
    LAYER via ;
      RECT 0.005000 0.265000 0.265000 0.525000 ;
      RECT 0.005000 0.585000 0.265000 0.845000 ;
      RECT 0.005000 0.905000 0.265000 1.165000 ;
      RECT 0.005000 1.225000 0.265000 1.485000 ;
      RECT 0.005000 1.545000 0.265000 1.805000 ;
      RECT 0.005000 1.865000 0.265000 2.125000 ;
      RECT 0.005000 2.185000 0.265000 2.445000 ;
      RECT 0.005000 2.505000 0.265000 2.765000 ;
      RECT 0.005000 2.825000 0.265000 3.085000 ;
      RECT 0.005000 3.145000 0.265000 3.405000 ;
      RECT 0.005000 3.465000 0.265000 3.725000 ;
      RECT 0.005000 3.785000 0.265000 4.045000 ;
      RECT 0.005000 4.105000 0.265000 4.365000 ;
      RECT 0.005000 4.425000 0.265000 4.685000 ;
      RECT 0.005000 4.745000 0.265000 5.005000 ;
      RECT 0.005000 5.065000 0.265000 5.325000 ;
      RECT 0.005000 5.385000 0.265000 5.645000 ;
      RECT 0.005000 5.705000 0.265000 5.965000 ;
      RECT 0.005000 6.025000 0.265000 6.285000 ;
      RECT 0.005000 6.345000 0.265000 6.605000 ;
      RECT 0.005000 6.665000 0.265000 6.925000 ;
      RECT 0.005000 6.985000 0.265000 7.245000 ;
      RECT 0.380000 0.030000 0.640000 0.290000 ;
      RECT 0.380000 7.550000 0.640000 7.810000 ;
      RECT 0.700000 0.030000 0.960000 0.290000 ;
      RECT 0.700000 7.550000 0.960000 7.810000 ;
      RECT 1.020000 0.030000 1.280000 0.290000 ;
      RECT 1.020000 7.550000 1.280000 7.810000 ;
      RECT 1.340000 0.030000 1.600000 0.290000 ;
      RECT 1.340000 7.550000 1.600000 7.810000 ;
      RECT 1.660000 0.030000 1.920000 0.290000 ;
      RECT 1.660000 7.550000 1.920000 7.810000 ;
      RECT 1.980000 0.030000 2.240000 0.290000 ;
      RECT 1.980000 7.550000 2.240000 7.810000 ;
      RECT 2.300000 0.030000 2.560000 0.290000 ;
      RECT 2.300000 7.550000 2.560000 7.810000 ;
      RECT 2.620000 0.030000 2.880000 0.290000 ;
      RECT 2.620000 7.550000 2.880000 7.810000 ;
      RECT 2.940000 0.030000 3.200000 0.290000 ;
      RECT 2.940000 7.550000 3.200000 7.810000 ;
      RECT 3.260000 0.030000 3.520000 0.290000 ;
      RECT 3.260000 7.550000 3.520000 7.810000 ;
      RECT 3.580000 0.030000 3.840000 0.290000 ;
      RECT 3.580000 7.550000 3.840000 7.810000 ;
      RECT 3.900000 0.030000 4.160000 0.290000 ;
      RECT 3.900000 7.550000 4.160000 7.810000 ;
      RECT 4.220000 0.030000 4.480000 0.290000 ;
      RECT 4.220000 7.550000 4.480000 7.810000 ;
      RECT 4.540000 0.030000 4.800000 0.290000 ;
      RECT 4.540000 7.550000 4.800000 7.810000 ;
      RECT 4.860000 0.030000 5.120000 0.290000 ;
      RECT 4.860000 7.550000 5.120000 7.810000 ;
      RECT 5.180000 0.030000 5.440000 0.290000 ;
      RECT 5.180000 7.550000 5.440000 7.810000 ;
      RECT 5.500000 0.030000 5.760000 0.290000 ;
      RECT 5.500000 7.550000 5.760000 7.810000 ;
      RECT 5.820000 0.030000 6.080000 0.290000 ;
      RECT 5.820000 7.550000 6.080000 7.810000 ;
      RECT 6.140000 0.030000 6.400000 0.290000 ;
      RECT 6.140000 7.550000 6.400000 7.810000 ;
      RECT 6.460000 0.030000 6.720000 0.290000 ;
      RECT 6.460000 7.550000 6.720000 7.810000 ;
      RECT 6.780000 0.030000 7.040000 0.290000 ;
      RECT 6.780000 7.550000 7.040000 7.810000 ;
      RECT 7.100000 0.030000 7.360000 0.290000 ;
      RECT 7.100000 7.550000 7.360000 7.810000 ;
      RECT 7.420000 0.030000 7.680000 0.290000 ;
      RECT 7.420000 7.550000 7.680000 7.810000 ;
      RECT 7.740000 0.030000 8.000000 0.290000 ;
      RECT 7.740000 7.550000 8.000000 7.810000 ;
      RECT 8.060000 0.030000 8.320000 0.290000 ;
      RECT 8.060000 7.550000 8.320000 7.810000 ;
      RECT 8.315000 0.490000 8.575000 0.750000 ;
      RECT 8.315000 0.810000 8.575000 1.070000 ;
      RECT 8.315000 1.130000 8.575000 1.390000 ;
      RECT 8.315000 1.450000 8.575000 1.710000 ;
      RECT 8.315000 1.770000 8.575000 2.030000 ;
      RECT 8.315000 2.090000 8.575000 2.350000 ;
      RECT 8.315000 2.410000 8.575000 2.670000 ;
      RECT 8.315000 2.730000 8.575000 2.990000 ;
      RECT 8.315000 3.050000 8.575000 3.310000 ;
      RECT 8.315000 3.370000 8.575000 3.630000 ;
      RECT 8.315000 3.690000 8.575000 3.950000 ;
      RECT 8.315000 4.010000 8.575000 4.270000 ;
      RECT 8.315000 4.330000 8.575000 4.590000 ;
      RECT 8.315000 4.650000 8.575000 4.910000 ;
      RECT 8.315000 4.970000 8.575000 5.230000 ;
      RECT 8.315000 5.290000 8.575000 5.550000 ;
      RECT 8.315000 5.610000 8.575000 5.870000 ;
      RECT 8.315000 5.930000 8.575000 6.190000 ;
      RECT 8.315000 6.250000 8.575000 6.510000 ;
      RECT 8.315000 6.570000 8.575000 6.830000 ;
      RECT 8.315000 6.890000 8.575000 7.150000 ;
      RECT 8.315000 7.210000 8.575000 7.470000 ;
  END
END sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o2subcell
END LIBRARY
