# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_test_coil1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_test_coil1 ;
  ORIGIN  72.52000  72.52000 ;
  SIZE  150.0200 BY  145.0400 ;
  OBS
    LAYER met2 ;
      POLYGON  -6.555000  55.010000  3.455000  55.010000  3.455000  45.000000 ;
      POLYGON  -3.445000 -65.020000  4.055000 -65.020000 -3.445000 -72.520000 ;
      POLYGON  -3.445000  62.510000  4.055000  55.010000 -3.445000  55.010000 ;
      POLYGON   3.455000 -55.010000  3.455000 -65.020000 -6.555000 -65.020000 ;
      POLYGON   4.055000 -62.510000  6.565000 -62.510000  4.055000 -65.020000 ;
      POLYGON   4.055000  55.010000  6.565000  52.500000  4.055000  52.500000 ;
      RECT -20.615000 -72.520000 -3.445000 -65.020000 ;
      RECT -20.395000  55.010000 -3.445000  62.510000 ;
      RECT   3.455000 -65.020000  4.055000 -62.510000 ;
      RECT   3.455000 -62.510000 19.625000 -55.010000 ;
      RECT   3.455000  45.000000 20.120000  52.500000 ;
      RECT   3.455000  52.500000  4.055000  55.010000 ;
      RECT  32.040000  -3.750000 77.500000   3.750000 ;
    LAYER met3 ;
      POLYGON -72.520000 -30.045000 -66.055000 -30.045000 -66.055000 -36.510000 ;
      POLYGON -66.055000 -36.510000 -55.445000 -36.510000 -55.445000 -47.120000 ;
      POLYGON -65.020000 -26.935000 -62.510000 -29.445000 -65.020000 -29.445000 ;
      POLYGON -65.020000  30.045000 -61.910000  30.045000 -65.020000  26.935000 ;
      POLYGON -62.510000 -29.445000 -58.990000 -32.965000 -62.510000 -32.965000 ;
      POLYGON -62.510000 -25.900000 -61.475000 -25.900000 -61.475000 -26.935000 ;
      POLYGON -61.910000  30.680000 -61.275000  30.680000 -61.910000  30.045000 ;
      POLYGON -61.910000  40.655000 -61.910000  30.045000 -72.520000  30.045000 ;
      POLYGON -61.475000 -26.935000 -58.965000 -26.935000 -58.965000 -29.445000 ;
      POLYGON -61.475000  26.935000 -61.475000  25.900000 -62.510000  25.900000 ;
      POLYGON -61.275000  34.225000 -57.730000  34.225000 -61.275000  30.680000 ;
      POLYGON -58.990000 -32.965000 -55.445000 -36.510000 -58.990000 -36.510000 ;
      POLYGON -58.965000 -29.445000 -55.445000 -29.445000 -55.445000 -32.965000 ;
      POLYGON -58.965000  29.445000 -58.965000  26.935000 -61.475000  26.935000 ;
      POLYGON -58.365000  30.045000 -58.365000  29.445000 -58.965000  29.445000 ;
      POLYGON -57.730000  30.680000 -57.730000  30.045000 -58.365000  30.045000 ;
      POLYGON -57.730000  37.110000 -54.845000  37.110000 -57.730000  34.225000 ;
      POLYGON -55.695000  46.870000 -55.695000  40.655000 -61.910000  40.655000 ;
      POLYGON -55.445000 -47.120000 -44.835000 -47.120000 -44.835000 -57.730000 ;
      POLYGON -55.445000 -36.510000 -51.900000 -40.055000 -55.445000 -40.055000 ;
      POLYGON -55.445000 -32.965000 -51.900000 -32.965000 -51.900000 -36.510000 ;
      POLYGON -55.010000 -22.790000 -52.500000 -25.300000 -55.010000 -25.300000 ;
      POLYGON -55.010000  25.300000 -52.500000  25.300000 -55.010000  22.790000 ;
      POLYGON -54.845000  40.655000 -51.300000  40.655000 -54.845000  37.110000 ;
      POLYGON -54.415000  48.150000 -54.415000  46.870000 -55.695000  46.870000 ;
      POLYGON -54.185000  34.225000 -54.185000  30.680000 -57.730000  30.680000 ;
      POLYGON -52.500000 -25.300000 -50.865000 -26.935000 -52.500000 -26.935000 ;
      POLYGON -52.500000 -21.755000 -51.465000 -21.755000 -51.465000 -22.790000 ;
      POLYGON -52.500000  26.935000 -50.865000  26.935000 -52.500000  25.300000 ;
      POLYGON -51.900000 -40.055000 -48.380000 -43.575000 -51.900000 -43.575000 ;
      POLYGON -51.900000 -36.510000 -48.355000 -36.510000 -48.355000 -40.055000 ;
      POLYGON -51.465000 -22.790000 -48.955000 -22.790000 -48.955000 -25.300000 ;
      POLYGON -51.465000  22.790000 -51.465000  21.755000 -52.500000  21.755000 ;
      POLYGON -51.300000  37.110000 -51.300000  34.225000 -54.185000  34.225000 ;
      POLYGON -51.300000  41.290000 -50.665000  41.290000 -51.300000  40.655000 ;
      POLYGON -50.865000 -26.935000 -47.720000 -30.080000 -50.865000 -30.080000 ;
      POLYGON -50.865000  30.045000 -47.755000  30.045000 -50.865000  26.935000 ;
      POLYGON -50.665000  44.835000 -47.120000  44.835000 -50.665000  41.290000 ;
      POLYGON -48.955000 -25.300000 -47.320000 -25.300000 -47.320000 -26.935000 ;
      POLYGON -48.955000  25.300000 -48.955000  22.790000 -51.465000  22.790000 ;
      POLYGON -48.380000 -43.575000 -44.835000 -47.120000 -48.380000 -47.120000 ;
      POLYGON -48.355000 -40.055000 -44.835000 -40.055000 -44.835000 -43.575000 ;
      POLYGON -47.755000  31.280000 -46.520000  31.280000 -47.755000  30.045000 ;
      POLYGON -47.755000  40.655000 -47.755000  37.110000 -51.300000  37.110000 ;
      POLYGON -47.720000 -30.080000 -45.435000 -32.365000 -47.720000 -32.365000 ;
      POLYGON -47.320000 -26.935000 -44.175000 -26.935000 -44.175000 -30.080000 ;
      POLYGON -47.320000  26.935000 -47.320000  25.300000 -48.955000  25.300000 ;
      POLYGON -47.120000  41.290000 -47.120000  40.655000 -47.755000  40.655000 ;
      POLYGON -47.120000  46.870000 -45.085000  46.870000 -47.120000  44.835000 ;
      POLYGON -46.520000  34.825000 -42.975000  34.825000 -46.520000  31.280000 ;
      POLYGON -45.680000  56.885000 -45.680000  48.150000 -54.415000  48.150000 ;
      POLYGON -45.435000 -32.365000 -41.890000 -35.910000 -45.435000 -35.910000 ;
      POLYGON -45.085000  49.340000 -42.615000  49.340000 -45.085000  46.870000 ;
      POLYGON -45.000000 -18.645000 -36.710000 -26.935000 -45.000000 -26.935000 ;
      POLYGON -45.000000  26.935000 -36.710000  26.935000 -45.000000  18.645000 ;
      POLYGON -44.835000 -57.730000 -40.055000 -57.730000 -40.055000 -62.510000 ;
      POLYGON -44.835000 -47.120000 -41.290000 -50.665000 -44.835000 -50.665000 ;
      POLYGON -44.835000 -43.575000 -41.290000 -43.575000 -41.290000 -47.120000 ;
      POLYGON -44.210000  30.045000 -44.210000  26.935000 -47.320000  26.935000 ;
      POLYGON -44.175000 -30.080000 -41.890000 -30.080000 -41.890000 -32.365000 ;
      POLYGON -43.575000  44.835000 -43.575000  41.290000 -47.120000  41.290000 ;
      POLYGON -43.210000  59.355000 -43.210000  56.885000 -45.680000  56.885000 ;
      POLYGON -42.975000  31.280000 -42.975000  30.045000 -44.210000  30.045000 ;
      POLYGON -42.975000  37.110000 -40.690000  37.110000 -42.975000  34.825000 ;
      POLYGON -42.615000  51.900000 -40.055000  51.900000 -42.615000  49.340000 ;
      POLYGON -41.890000 -35.910000 -40.690000 -37.110000 -41.890000 -37.110000 ;
      POLYGON -41.890000 -32.365000 -38.345000 -32.365000 -38.345000 -35.910000 ;
      POLYGON -41.540000  46.870000 -41.540000  44.835000 -43.575000  44.835000 ;
      POLYGON -41.290000 -50.665000 -40.480000 -51.475000 -41.290000 -51.475000 ;
      POLYGON -41.290000 -47.120000 -37.745000 -47.120000 -37.745000 -50.665000 ;
      POLYGON -40.690000 -37.110000 -37.145000 -40.655000 -40.690000 -40.655000 ;
      POLYGON -40.690000  40.655000 -37.145000  40.655000 -40.690000  37.110000 ;
      POLYGON -40.480000 -51.475000 -36.935000 -55.020000 -40.480000 -55.020000 ;
      POLYGON -40.055000 -62.510000 -30.045000 -62.510000 -30.045000 -72.520000 ;
      POLYGON -40.055000  55.445000 -36.510000  55.445000 -40.055000  51.900000 ;
      POLYGON -39.430000  34.825000 -39.430000  31.280000 -42.975000  31.280000 ;
      POLYGON -39.070000  49.340000 -39.070000  46.870000 -41.540000  46.870000 ;
      POLYGON -38.345000 -35.910000 -37.145000 -35.910000 -37.145000 -37.110000 ;
      POLYGON -37.745000 -50.665000 -36.935000 -50.665000 -36.935000 -51.475000 ;
      POLYGON -37.545000  65.020000 -37.545000  59.355000 -43.210000  59.355000 ;
      POLYGON -37.145000 -40.655000 -34.825000 -42.975000 -37.145000 -42.975000 ;
      POLYGON -37.145000 -37.110000 -33.600000 -37.110000 -33.600000 -40.655000 ;
      POLYGON -37.145000  37.110000 -37.145000  34.825000 -39.430000  34.825000 ;
      POLYGON -37.145000  41.890000 -35.910000  41.890000 -37.145000  40.655000 ;
      POLYGON -36.935000 -55.020000 -33.790000 -58.165000 -36.935000 -58.165000 ;
      POLYGON -36.935000 -51.475000 -33.390000 -51.475000 -33.390000 -55.020000 ;
      POLYGON -36.710000 -26.935000 -27.135000 -36.510000 -36.710000 -36.510000 ;
      POLYGON -36.710000  36.510000 -27.135000  36.510000 -36.710000  26.935000 ;
      POLYGON -36.510000  51.900000 -36.510000  49.340000 -39.070000  49.340000 ;
      POLYGON -36.510000  58.330000 -33.625000  58.330000 -36.510000  55.445000 ;
      POLYGON -35.910000  45.000000 -32.800000  45.000000 -35.910000  41.890000 ;
      POLYGON -34.825000 -42.975000 -31.280000 -46.520000 -34.825000 -46.520000 ;
      POLYGON -33.790000 -58.165000 -30.680000 -61.275000 -33.790000 -61.275000 ;
      POLYGON -33.625000  61.875000 -30.080000  61.875000 -33.625000  58.330000 ;
      POLYGON -33.600000 -40.655000 -31.280000 -40.655000 -31.280000 -42.975000 ;
      POLYGON -33.600000  40.655000 -33.600000  37.110000 -37.145000  37.110000 ;
      POLYGON -33.390000 -55.020000 -30.245000 -55.020000 -30.245000 -58.165000 ;
      POLYGON -32.965000  55.445000 -32.965000  51.900000 -36.510000  51.900000 ;
      POLYGON -32.800000  48.355000 -29.445000  48.355000 -32.800000  45.000000 ;
      POLYGON -32.365000  41.890000 -32.365000  40.655000 -33.600000  40.655000 ;
      POLYGON -31.525000  56.885000 -31.525000  55.445000 -32.965000  55.445000 ;
      POLYGON -31.280000 -46.520000 -30.080000 -47.720000 -31.280000 -47.720000 ;
      POLYGON -31.280000 -42.975000 -27.735000 -42.975000 -27.735000 -46.520000 ;
      POLYGON -30.680000 -61.275000 -29.445000 -62.510000 -30.680000 -62.510000 ;
      POLYGON -30.245000 -58.165000 -27.135000 -58.165000 -27.135000 -61.275000 ;
      POLYGON -30.080000 -47.720000 -26.535000 -51.265000 -30.080000 -51.265000 ;
      POLYGON -30.080000  58.330000 -30.080000  56.885000 -31.525000  56.885000 ;
      POLYGON -30.080000  65.020000 -26.935000  65.020000 -30.080000  61.875000 ;
      POLYGON -30.045000  72.520000 -30.045000  65.020000 -37.545000  65.020000 ;
      POLYGON -29.445000 -62.510000 -26.935000 -65.020000 -29.445000 -65.020000 ;
      POLYGON -29.445000  51.900000 -25.900000  51.900000 -29.445000  48.355000 ;
      POLYGON -29.255000  45.000000 -29.255000  41.890000 -32.365000  41.890000 ;
      POLYGON -27.735000 -46.520000 -26.535000 -46.520000 -26.535000 -47.720000 ;
      POLYGON -27.135000 -61.275000 -25.900000 -61.275000 -25.900000 -62.510000 ;
      POLYGON -27.135000 -36.510000 -18.645000 -45.000000 -27.135000 -45.000000 ;
      POLYGON -27.135000  45.000000 -18.645000  45.000000 -27.135000  36.510000 ;
      POLYGON -26.535000 -51.265000 -25.300000 -52.500000 -26.535000 -52.500000 ;
      POLYGON -26.535000 -47.720000 -22.990000 -47.720000 -22.990000 -51.265000 ;
      POLYGON -26.535000  61.875000 -26.535000  58.330000 -30.080000  58.330000 ;
      POLYGON -25.900000  48.355000 -25.900000  45.000000 -29.255000  45.000000 ;
      POLYGON -25.900000  55.010000 -22.790000  55.010000 -25.900000  51.900000 ;
      POLYGON -25.900000  62.510000 -25.900000  61.875000 -26.535000  61.875000 ;
      POLYGON -25.300000 -52.500000 -22.780000 -55.020000 -25.300000 -55.020000 ;
      POLYGON -22.990000 -51.265000 -21.755000 -51.265000 -21.755000 -52.500000 ;
      POLYGON -22.355000  51.900000 -22.355000  48.355000 -25.900000  48.355000 ;
      POLYGON -21.755000  52.500000 -21.755000  51.900000 -22.355000  51.900000 ;
      POLYGON  -8.915000 -71.150000  -7.545000 -71.150000  -8.915000 -72.520000 ;
      POLYGON  -8.915000 -65.020000  -7.545000 -66.390000  -8.915000 -66.390000 ;
      POLYGON  -8.695000  56.380000  -7.325000  56.380000  -8.695000  55.010000 ;
      POLYGON  -8.695000  62.510000  -7.325000  61.140000  -8.695000  61.140000 ;
      POLYGON  -6.565000 -62.510000  -4.055000 -62.510000  -4.055000 -65.020000 ;
      POLYGON  -4.055000 -65.020000   3.445000 -65.020000   3.445000 -72.520000 ;
      POLYGON  -4.055000  55.010000  -4.055000  52.500000  -6.565000  52.500000 ;
      POLYGON  -3.455000  50.620000   2.165000  50.620000  -3.455000  45.000000 ;
      POLYGON  -3.445000 -55.020000   6.555000 -65.020000  -3.445000 -65.020000 ;
      POLYGON  -2.685000  56.380000  -2.685000  55.010000  -4.055000  55.010000 ;
      POLYGON   2.075000  61.140000   2.075000  56.380000  -2.685000  56.380000 ;
      POLYGON   2.165000  55.010000   6.555000  55.010000   2.165000  50.620000 ;
      POLYGON   2.810000  61.875000   2.810000  61.140000   2.075000  61.140000 ;
      POLYGON   3.445000  62.510000   3.445000  61.875000   2.810000  61.875000 ;
      POLYGON   6.555000 -61.140000   7.925000 -61.140000   7.925000 -62.510000 ;
      POLYGON   7.050000  46.370000   8.420000  46.370000   8.420000  45.000000 ;
      POLYGON   7.915000 -55.020000   7.915000 -56.380000   6.555000 -56.380000 ;
      POLYGON   7.925000 -55.010000   7.925000 -55.020000   7.915000 -55.020000 ;
      POLYGON   8.420000  52.500000   8.420000  51.130000   7.050000  51.130000 ;
      POLYGON  18.645000  45.000000  27.135000  45.000000  27.135000  36.510000 ;
      POLYGON  21.755000 -51.265000  22.990000 -51.265000  21.755000 -52.500000 ;
      POLYGON  21.755000  52.500000  22.990000  51.265000  21.755000  51.265000 ;
      POLYGON  22.790000  55.010000  25.300000  55.010000  25.300000  52.500000 ;
      POLYGON  22.990000 -47.720000  26.535000 -47.720000  22.990000 -51.265000 ;
      POLYGON  22.990000  51.265000  26.535000  47.720000  22.990000  47.720000 ;
      POLYGON  25.300000 -52.500000  25.300000 -55.010000  22.790000 -55.010000 ;
      POLYGON  25.300000  52.500000  26.535000  52.500000  26.535000  51.265000 ;
      POLYGON  25.900000 -61.910000  26.500000 -61.910000  25.900000 -62.510000 ;
      POLYGON  25.900000  62.510000  26.535000  61.875000  25.900000  61.875000 ;
      POLYGON  26.500000 -58.365000  30.045000 -58.365000  26.500000 -61.910000 ;
      POLYGON  26.535000 -51.265000  26.535000 -52.500000  25.300000 -52.500000 ;
      POLYGON  26.535000 -45.435000  28.820000 -45.435000  26.535000 -47.720000 ;
      POLYGON  26.535000  47.720000  29.255000  45.000000  26.535000  45.000000 ;
      POLYGON  26.535000  51.265000  30.080000  51.265000  30.080000  47.720000 ;
      POLYGON  26.535000  61.875000  27.135000  61.275000  26.535000  61.275000 ;
      POLYGON  26.935000  65.020000  29.445000  65.020000  29.445000  62.510000 ;
      POLYGON  27.135000 -36.510000  27.135000 -45.000000  18.645000 -45.000000 ;
      POLYGON  27.135000  36.510000  36.710000  36.510000  36.710000  26.935000 ;
      POLYGON  27.135000  61.275000  30.680000  57.730000  27.135000  57.730000 ;
      POLYGON  28.820000 -41.890000  32.365000 -41.890000  28.820000 -45.435000 ;
      POLYGON  29.255000  45.000000  31.280000  42.975000  29.255000  42.975000 ;
      POLYGON  29.445000 -62.510000  29.445000 -65.020000  26.935000 -65.020000 ;
      POLYGON  29.445000  62.510000  30.080000  62.510000  30.080000  61.875000 ;
      POLYGON  30.045000 -61.910000  30.045000 -62.510000  29.445000 -62.510000 ;
      POLYGON  30.045000 -61.910000  40.655000 -61.910000  30.045000 -72.520000 ;
      POLYGON  30.045000 -55.445000  32.965000 -55.445000  30.045000 -58.365000 ;
      POLYGON  30.045000  72.520000  37.545000  65.020000  30.045000  65.020000 ;
      POLYGON  30.080000 -47.720000  30.080000 -51.265000  26.535000 -51.265000 ;
      POLYGON  30.080000  47.720000  32.800000  47.720000  32.800000  45.000000 ;
      POLYGON  30.080000  61.875000  30.680000  61.875000  30.680000  61.275000 ;
      POLYGON  30.680000  57.730000  34.225000  54.185000  30.680000  54.185000 ;
      POLYGON  30.680000  61.275000  34.225000  61.275000  34.225000  57.730000 ;
      POLYGON  31.280000 -32.365000  31.280000 -36.510000  27.135000 -36.510000 ;
      POLYGON  31.280000  42.975000  33.600000  40.655000  31.280000  40.655000 ;
      POLYGON  32.365000 -45.435000  32.365000 -47.720000  30.080000 -47.720000 ;
      POLYGON  32.365000 -40.655000  33.600000 -40.655000  32.365000 -41.890000 ;
      POLYGON  32.365000 -31.280000  32.365000 -32.365000  31.280000 -32.365000 ;
      POLYGON  32.800000  45.000000  34.825000  45.000000  34.825000  42.975000 ;
      POLYGON  32.965000 -51.900000  36.510000 -51.900000  32.965000 -55.445000 ;
      POLYGON  33.590000 -58.365000  33.590000 -61.910000  30.045000 -61.910000 ;
      POLYGON  33.600000 -37.110000  37.145000 -37.110000  33.600000 -40.655000 ;
      POLYGON  33.600000  40.655000  37.145000  37.110000  33.600000  37.110000 ;
      POLYGON  34.225000  54.185000  37.745000  50.665000  34.225000  50.665000 ;
      POLYGON  34.225000  57.730000  37.770000  57.730000  37.770000  54.185000 ;
      POLYGON  34.825000  42.975000  37.145000  42.975000  37.145000  40.655000 ;
      POLYGON  35.910000 -41.890000  35.910000 -45.435000  32.365000 -45.435000 ;
      POLYGON  36.510000 -55.445000  36.510000 -58.365000  33.590000 -58.365000 ;
      POLYGON  36.510000 -51.300000  37.110000 -51.300000  36.510000 -51.900000 ;
      POLYGON  36.710000 -26.935000  36.710000 -31.280000  32.365000 -31.280000 ;
      POLYGON  36.710000  26.935000  45.000000  26.935000  45.000000  18.645000 ;
      POLYGON  37.110000 -47.755000  40.655000 -47.755000  37.110000 -51.300000 ;
      POLYGON  37.145000 -40.655000  37.145000 -41.890000  35.910000 -41.890000 ;
      POLYGON  37.145000 -34.825000  39.430000 -34.825000  37.145000 -37.110000 ;
      POLYGON  37.145000  37.110000  38.345000  35.910000  37.145000  35.910000 ;
      POLYGON  37.145000  40.655000  40.690000  40.655000  40.690000  37.110000 ;
      POLYGON  37.545000  65.020000  44.835000  57.730000  37.545000  57.730000 ;
      POLYGON  37.745000  50.665000  41.290000  47.120000  37.745000  47.120000 ;
      POLYGON  37.770000  54.185000  41.290000  54.185000  41.290000  50.665000 ;
      POLYGON  38.345000  35.910000  41.890000  32.365000  38.345000  32.365000 ;
      POLYGON  39.430000 -31.280000  42.975000 -31.280000  39.430000 -34.825000 ;
      POLYGON  40.055000 -51.900000  40.055000 -55.445000  36.510000 -55.445000 ;
      POLYGON  40.655000 -51.300000  40.655000 -51.900000  40.055000 -51.900000 ;
      POLYGON  40.655000 -51.300000  51.265000 -51.300000  40.655000 -61.910000 ;
      POLYGON  40.655000 -44.835000  43.575000 -44.835000  40.655000 -47.755000 ;
      POLYGON  40.690000 -37.110000  40.690000 -40.655000  37.145000 -40.655000 ;
      POLYGON  40.690000  37.110000  41.890000  37.110000  41.890000  35.910000 ;
      POLYGON  40.855000 -22.790000  40.855000 -26.935000  36.710000 -26.935000 ;
      POLYGON  41.290000  47.120000  44.835000  43.575000  41.290000  43.575000 ;
      POLYGON  41.290000  50.665000  44.835000  50.665000  44.835000  47.120000 ;
      POLYGON  41.890000  32.365000  44.210000  30.045000  41.890000  30.045000 ;
      POLYGON  41.890000  35.910000  45.435000  35.910000  45.435000  32.365000 ;
      POLYGON  42.975000 -34.825000  42.975000 -37.110000  40.690000 -37.110000 ;
      POLYGON  42.975000 -30.080000  44.175000 -30.080000  42.975000 -31.280000 ;
      POLYGON  43.575000 -41.290000  47.120000 -41.290000  43.575000 -44.835000 ;
      POLYGON  44.175000 -26.935000  47.320000 -26.935000  44.175000 -30.080000 ;
      POLYGON  44.200000 -47.755000  44.200000 -51.300000  40.655000 -51.300000 ;
      POLYGON  44.210000  30.045000  47.320000  26.935000  44.210000  26.935000 ;
      POLYGON  44.835000  43.575000  48.355000  40.055000  44.835000  40.055000 ;
      POLYGON  44.835000  47.120000  48.380000  47.120000  48.380000  43.575000 ;
      POLYGON  44.835000  57.730000  55.445000  47.120000  44.835000  47.120000 ;
      POLYGON  45.000000 -18.645000  45.000000 -22.790000  40.855000 -22.790000 ;
      POLYGON  45.435000  32.365000  47.755000  32.365000  47.755000  30.045000 ;
      POLYGON  46.520000 -31.280000  46.520000 -34.825000  42.975000 -34.825000 ;
      POLYGON  47.120000 -44.835000  47.120000 -47.755000  44.200000 -47.755000 ;
      POLYGON  47.120000 -40.690000  47.720000 -40.690000  47.120000 -41.290000 ;
      POLYGON  47.320000 -25.300000  48.955000 -25.300000  47.320000 -26.935000 ;
      POLYGON  47.320000  26.935000  48.955000  25.300000  47.320000  25.300000 ;
      POLYGON  47.720000 -37.145000  51.265000 -37.145000  47.720000 -40.690000 ;
      POLYGON  47.720000 -30.080000  47.720000 -31.280000  46.520000 -31.280000 ;
      POLYGON  47.755000  30.045000  50.865000  30.045000  50.865000  26.935000 ;
      POLYGON  48.355000  40.055000  51.900000  36.510000  48.355000  36.510000 ;
      POLYGON  48.380000  43.575000  51.900000  43.575000  51.900000  40.055000 ;
      POLYGON  48.955000 -21.755000  52.500000 -21.755000  48.955000 -25.300000 ;
      POLYGON  48.955000  25.300000  52.500000  21.755000  48.955000  21.755000 ;
      POLYGON  50.665000 -41.290000  50.665000 -44.835000  47.120000 -44.835000 ;
      POLYGON  50.865000 -26.935000  50.865000 -30.080000  47.720000 -30.080000 ;
      POLYGON  50.865000  26.935000  52.500000  26.935000  52.500000  25.300000 ;
      POLYGON  51.265000 -41.290000  61.275000 -41.290000  51.265000 -51.300000 ;
      POLYGON  51.265000 -40.690000  51.265000 -41.290000  50.665000 -41.290000 ;
      POLYGON  51.265000 -34.225000  54.185000 -34.225000  51.265000 -37.145000 ;
      POLYGON  51.900000  36.510000  55.445000  32.965000  51.900000  32.965000 ;
      POLYGON  51.900000  40.055000  55.445000  40.055000  55.445000  36.510000 ;
      POLYGON  52.500000 -25.300000  52.500000 -26.935000  50.865000 -26.935000 ;
      POLYGON  52.500000  25.300000  55.010000  25.300000  55.010000  22.790000 ;
      POLYGON  54.185000 -30.680000  57.730000 -30.680000  54.185000 -34.225000 ;
      POLYGON  54.810000 -37.145000  54.810000 -40.690000  51.265000 -40.690000 ;
      POLYGON  55.010000 -22.790000  55.010000 -25.300000  52.500000 -25.300000 ;
      POLYGON  55.445000  32.965000  58.965000  29.445000  55.445000  29.445000 ;
      POLYGON  55.445000  36.510000  58.990000  36.510000  58.990000  32.965000 ;
      POLYGON  55.445000  47.120000  66.055000  36.510000  55.445000  36.510000 ;
      POLYGON  57.730000 -34.225000  57.730000 -37.145000  54.810000 -37.145000 ;
      POLYGON  57.730000 -29.445000  58.965000 -29.445000  57.730000 -30.680000 ;
      POLYGON  58.965000 -25.900000  62.510000 -25.900000  58.965000 -29.445000 ;
      POLYGON  58.965000  29.445000  62.510000  25.900000  58.965000  25.900000 ;
      POLYGON  58.990000  32.965000  62.510000  32.965000  62.510000  29.445000 ;
      POLYGON  61.275000 -30.680000  61.275000 -34.225000  57.730000 -34.225000 ;
      POLYGON  61.275000 -30.680000  71.885000 -30.680000  61.275000 -41.290000 ;
      POLYGON  62.510000 -29.445000  62.510000 -30.680000  61.275000 -30.680000 ;
      POLYGON  62.510000  29.445000  65.020000  29.445000  65.020000  26.935000 ;
      POLYGON  65.020000 -26.935000  65.020000 -29.445000  62.510000 -29.445000 ;
      POLYGON  66.055000  36.510000  72.520000  30.045000  66.055000  30.045000 ;
      POLYGON  71.885000 -30.045000  72.520000 -30.045000  71.885000 -30.680000 ;
      RECT -72.520000 -30.045000 -62.510000 -29.445000 ;
      RECT -72.520000 -29.445000 -65.020000  30.045000 ;
      RECT -66.055000 -36.510000 -58.990000 -32.965000 ;
      RECT -66.055000 -32.965000 -62.510000 -30.045000 ;
      RECT -62.510000 -25.900000 -52.500000 -25.300000 ;
      RECT -62.510000 -25.300000 -55.010000  25.300000 ;
      RECT -62.510000  25.300000 -52.500000  25.900000 ;
      RECT -61.910000  30.680000 -61.275000  34.225000 ;
      RECT -61.910000  34.225000 -57.730000  37.110000 ;
      RECT -61.910000  37.110000 -54.845000  40.655000 ;
      RECT -61.475000 -26.935000 -52.500000 -25.900000 ;
      RECT -61.475000  25.900000 -52.500000  26.935000 ;
      RECT -58.965000 -29.445000 -50.865000 -26.935000 ;
      RECT -58.965000  26.935000 -50.865000  29.445000 ;
      RECT -58.365000  29.445000 -50.865000  30.045000 ;
      RECT -57.730000  30.045000 -47.755000  30.680000 ;
      RECT -55.695000  40.655000 -51.300000  41.290000 ;
      RECT -55.695000  41.290000 -50.665000  44.835000 ;
      RECT -55.695000  44.835000 -47.120000  46.870000 ;
      RECT -55.445000 -47.120000 -48.380000 -43.575000 ;
      RECT -55.445000 -43.575000 -51.900000 -40.055000 ;
      RECT -55.445000 -32.965000 -45.435000 -32.365000 ;
      RECT -55.445000 -32.365000 -47.720000 -30.080000 ;
      RECT -55.445000 -30.080000 -50.865000 -29.445000 ;
      RECT -54.415000  46.870000 -45.085000  48.150000 ;
      RECT -54.185000  30.680000 -47.755000  31.280000 ;
      RECT -54.185000  31.280000 -46.520000  34.225000 ;
      RECT -52.500000 -21.755000 -45.000000  -3.750000 ;
      RECT -52.500000  -3.750000  40.000000   3.750000 ;
      RECT -52.500000   3.750000 -45.000000  21.755000 ;
      RECT -51.900000 -36.510000 -41.890000 -35.910000 ;
      RECT -51.900000 -35.910000 -45.435000 -32.965000 ;
      RECT -51.465000 -22.790000 -45.000000 -21.755000 ;
      RECT -51.465000  21.755000 -45.000000  22.790000 ;
      RECT -51.300000  34.225000 -46.520000  34.825000 ;
      RECT -51.300000  34.825000 -42.975000  37.110000 ;
      RECT -48.955000 -25.300000 -45.000000 -22.790000 ;
      RECT -48.955000  22.790000 -45.000000  25.300000 ;
      RECT -48.355000 -40.055000 -40.690000 -37.110000 ;
      RECT -48.355000 -37.110000 -41.890000 -36.510000 ;
      RECT -47.755000  37.110000 -40.690000  40.655000 ;
      RECT -47.320000 -26.935000 -45.000000 -25.300000 ;
      RECT -47.320000  25.300000 -45.000000  26.935000 ;
      RECT -47.120000  40.655000 -37.145000  41.290000 ;
      RECT -45.680000  48.150000 -45.085000  49.340000 ;
      RECT -45.680000  49.340000 -42.615000  51.900000 ;
      RECT -45.680000  51.900000 -40.055000  55.445000 ;
      RECT -45.680000  55.445000 -36.510000  56.885000 ;
      RECT -44.835000 -57.730000 -36.935000 -55.020000 ;
      RECT -44.835000 -55.020000 -40.480000 -51.475000 ;
      RECT -44.835000 -51.475000 -41.290000 -50.665000 ;
      RECT -44.835000 -43.575000 -34.825000 -42.975000 ;
      RECT -44.835000 -42.975000 -37.145000 -40.655000 ;
      RECT -44.835000 -40.655000 -40.690000 -40.055000 ;
      RECT -44.210000  26.935000 -36.710000  30.045000 ;
      RECT -44.175000 -30.080000 -36.710000 -26.935000 ;
      RECT -43.575000  41.290000 -37.145000  41.890000 ;
      RECT -43.575000  41.890000 -35.910000  44.835000 ;
      RECT -43.210000  56.885000 -36.510000  58.330000 ;
      RECT -43.210000  58.330000 -33.625000  59.355000 ;
      RECT -42.975000  30.045000 -36.710000  31.280000 ;
      RECT -41.890000 -32.365000 -36.710000 -30.080000 ;
      RECT -41.540000  44.835000 -35.910000  45.000000 ;
      RECT -41.540000  45.000000 -32.800000  46.870000 ;
      RECT -41.290000 -47.120000 -31.280000 -46.520000 ;
      RECT -41.290000 -46.520000 -34.825000 -43.575000 ;
      RECT -40.055000 -62.510000 -30.680000 -61.275000 ;
      RECT -40.055000 -61.275000 -33.790000 -58.165000 ;
      RECT -40.055000 -58.165000 -36.935000 -57.730000 ;
      RECT -39.430000  31.280000 -36.710000  34.825000 ;
      RECT -39.070000  46.870000 -32.800000  48.355000 ;
      RECT -39.070000  48.355000 -29.445000  49.340000 ;
      RECT -38.345000 -35.910000 -36.710000 -32.365000 ;
      RECT -37.745000 -50.665000 -30.080000 -47.720000 ;
      RECT -37.745000 -47.720000 -31.280000 -47.120000 ;
      RECT -37.545000  59.355000 -33.625000  61.875000 ;
      RECT -37.545000  61.875000 -30.080000  65.020000 ;
      RECT -37.145000 -37.110000 -27.135000 -36.510000 ;
      RECT -37.145000 -36.510000 -36.710000 -35.910000 ;
      RECT -37.145000  34.825000 -36.710000  36.510000 ;
      RECT -37.145000  36.510000 -27.135000  37.110000 ;
      RECT -36.935000 -51.475000 -26.535000 -51.265000 ;
      RECT -36.935000 -51.265000 -30.080000 -50.665000 ;
      RECT -36.510000  49.340000 -29.445000  51.900000 ;
      RECT -33.600000 -40.655000 -27.135000 -37.110000 ;
      RECT -33.600000  37.110000 -27.135000  40.655000 ;
      RECT -33.390000 -55.020000 -25.300000 -52.500000 ;
      RECT -33.390000 -52.500000 -26.535000 -51.475000 ;
      RECT -32.965000  51.900000 -25.900000  55.010000 ;
      RECT -32.965000  55.010000  -8.695000  55.445000 ;
      RECT -32.365000  40.655000 -27.135000  41.890000 ;
      RECT -31.525000  55.445000  -8.695000  56.380000 ;
      RECT -31.525000  56.380000  -7.265000  56.885000 ;
      RECT -31.280000 -42.975000 -27.135000 -40.655000 ;
      RECT -30.245000 -58.165000  -3.445000 -55.020000 ;
      RECT -30.080000  56.885000  -7.265000  58.330000 ;
      RECT -30.045000 -72.520000  -8.915000 -71.150000 ;
      RECT -30.045000 -71.150000  -7.545000 -66.390000 ;
      RECT -30.045000 -66.390000  -8.915000 -65.020000 ;
      RECT -30.045000 -65.020000 -29.445000 -62.510000 ;
      RECT -30.045000  65.020000  30.045000  72.520000 ;
      RECT -29.255000  41.890000 -27.135000  45.000000 ;
      RECT -27.735000 -46.520000  26.535000 -45.435000 ;
      RECT -27.735000 -45.435000  28.820000 -45.000000 ;
      RECT -27.735000 -45.000000 -27.135000 -42.975000 ;
      RECT -27.135000 -61.275000  -3.445000 -58.165000 ;
      RECT -26.535000 -47.720000  26.535000 -46.520000 ;
      RECT -26.535000  58.330000  -7.265000  61.140000 ;
      RECT -26.535000  61.140000  -8.695000  61.875000 ;
      RECT -25.900000 -62.510000  -3.445000 -61.275000 ;
      RECT -25.900000  45.000000  -3.455000  48.355000 ;
      RECT -25.900000  61.875000  -8.695000  62.510000 ;
      RECT -22.990000 -51.265000  22.990000 -47.720000 ;
      RECT -22.355000  48.355000  -3.455000  50.620000 ;
      RECT -22.355000  50.620000   2.165000  51.900000 ;
      RECT -21.755000 -52.500000  21.755000 -51.265000 ;
      RECT -21.755000  51.900000   2.165000  52.500000 ;
      RECT  -4.055000 -65.020000  -3.445000 -62.510000 ;
      RECT  -4.055000  52.500000   2.165000  55.010000 ;
      RECT  -2.685000  55.010000  30.680000  56.380000 ;
      RECT   2.075000  56.380000  30.680000  57.730000 ;
      RECT   2.075000  57.730000  27.135000  61.140000 ;
      RECT   2.810000  61.140000  27.135000  61.275000 ;
      RECT   2.810000  61.275000  26.535000  61.875000 ;
      RECT   3.445000 -72.520000  30.045000 -65.020000 ;
      RECT   3.445000  61.875000  25.900000  62.510000 ;
      RECT   6.555000 -61.140000  26.500000 -58.365000 ;
      RECT   6.555000 -58.365000  30.045000 -56.380000 ;
      RECT   7.050000  46.370000  26.535000  47.720000 ;
      RECT   7.050000  47.720000  22.990000  51.130000 ;
      RECT   7.915000 -56.380000  30.045000 -55.445000 ;
      RECT   7.915000 -55.445000  32.965000 -55.020000 ;
      RECT   7.925000 -62.510000  25.900000 -61.910000 ;
      RECT   7.925000 -61.910000  26.500000 -61.140000 ;
      RECT   7.925000 -55.020000  32.965000 -55.010000 ;
      RECT   8.420000  45.000000  26.535000  46.370000 ;
      RECT   8.420000  51.130000  22.990000  51.265000 ;
      RECT   8.420000  51.265000  21.755000  52.500000 ;
      RECT  25.300000 -55.010000  32.965000 -52.500000 ;
      RECT  25.300000  52.500000  34.225000  54.185000 ;
      RECT  25.300000  54.185000  30.680000  55.010000 ;
      RECT  26.535000 -52.500000  32.965000 -51.900000 ;
      RECT  26.535000 -51.900000  36.510000 -51.300000 ;
      RECT  26.535000 -51.300000  37.110000 -51.265000 ;
      RECT  26.535000  51.265000  34.225000  52.500000 ;
      RECT  27.135000 -45.000000  28.820000 -41.890000 ;
      RECT  27.135000 -41.890000  32.365000 -40.655000 ;
      RECT  27.135000 -40.655000  33.600000 -37.110000 ;
      RECT  27.135000 -37.110000  37.145000 -36.510000 ;
      RECT  27.135000  36.510000  37.145000  37.110000 ;
      RECT  27.135000  37.110000  33.600000  40.655000 ;
      RECT  27.135000  40.655000  31.280000  42.975000 ;
      RECT  27.135000  42.975000  29.255000  45.000000 ;
      RECT  29.445000 -65.020000  30.045000 -62.510000 ;
      RECT  29.445000  62.510000  37.545000  65.020000 ;
      RECT  30.080000 -51.265000  37.110000 -47.755000 ;
      RECT  30.080000 -47.755000  40.655000 -47.720000 ;
      RECT  30.080000  47.720000  37.745000  50.665000 ;
      RECT  30.080000  50.665000  34.225000  51.265000 ;
      RECT  30.080000  61.875000  37.545000  62.510000 ;
      RECT  30.680000  61.275000  37.545000  61.875000 ;
      RECT  31.280000 -36.510000  37.145000 -34.825000 ;
      RECT  31.280000 -34.825000  39.430000 -32.365000 ;
      RECT  32.365000 -47.720000  40.655000 -45.435000 ;
      RECT  32.365000 -32.365000  39.430000 -31.280000 ;
      RECT  32.800000  45.000000  41.290000  47.120000 ;
      RECT  32.800000  47.120000  37.745000  47.720000 ;
      RECT  33.590000 -61.910000  40.655000 -58.365000 ;
      RECT  34.225000  57.730000  37.545000  61.275000 ;
      RECT  34.825000  42.975000  44.835000  43.575000 ;
      RECT  34.825000  43.575000  41.290000  45.000000 ;
      RECT  35.910000 -45.435000  40.655000 -44.835000 ;
      RECT  35.910000 -44.835000  43.575000 -41.890000 ;
      RECT  36.510000 -58.365000  40.655000 -55.445000 ;
      RECT  36.710000 -31.280000  42.975000 -30.080000 ;
      RECT  36.710000 -30.080000  44.175000 -26.935000 ;
      RECT  36.710000  26.935000  44.210000  30.045000 ;
      RECT  36.710000  30.045000  41.890000  32.365000 ;
      RECT  36.710000  32.365000  38.345000  35.910000 ;
      RECT  36.710000  35.910000  37.145000  36.510000 ;
      RECT  37.145000 -41.890000  43.575000 -41.290000 ;
      RECT  37.145000 -41.290000  47.120000 -40.690000 ;
      RECT  37.145000 -40.690000  47.720000 -40.655000 ;
      RECT  37.145000  40.655000  44.835000  42.975000 ;
      RECT  37.770000  54.185000  44.835000  57.730000 ;
      RECT  40.055000 -55.445000  40.655000 -51.900000 ;
      RECT  40.690000 -40.655000  47.720000 -37.145000 ;
      RECT  40.690000 -37.145000  51.265000 -37.110000 ;
      RECT  40.690000  37.110000  48.355000  40.055000 ;
      RECT  40.690000  40.055000  44.835000  40.655000 ;
      RECT  40.855000 -26.935000  47.320000 -25.300000 ;
      RECT  40.855000 -25.300000  48.955000 -22.790000 ;
      RECT  41.290000  50.665000  44.835000  54.185000 ;
      RECT  41.890000  35.910000  51.900000  36.510000 ;
      RECT  41.890000  36.510000  48.355000  37.110000 ;
      RECT  42.975000 -37.110000  51.265000 -34.825000 ;
      RECT  44.200000 -51.300000  51.265000 -47.755000 ;
      RECT  45.000000 -22.790000  48.955000 -21.755000 ;
      RECT  45.000000 -21.755000  52.500000  21.755000 ;
      RECT  45.000000  21.755000  48.955000  25.300000 ;
      RECT  45.000000  25.300000  47.320000  26.935000 ;
      RECT  45.435000  32.365000  55.445000  32.965000 ;
      RECT  45.435000  32.965000  51.900000  35.910000 ;
      RECT  46.520000 -34.825000  51.265000 -34.225000 ;
      RECT  46.520000 -34.225000  54.185000 -31.280000 ;
      RECT  47.120000 -47.755000  51.265000 -44.835000 ;
      RECT  47.720000 -31.280000  54.185000 -30.680000 ;
      RECT  47.720000 -30.680000  57.730000 -30.080000 ;
      RECT  47.755000  30.045000  55.445000  32.365000 ;
      RECT  48.380000  43.575000  55.445000  47.120000 ;
      RECT  50.665000 -44.835000  51.265000 -41.290000 ;
      RECT  50.865000 -30.080000  57.730000 -29.445000 ;
      RECT  50.865000 -29.445000  58.965000 -26.935000 ;
      RECT  50.865000  26.935000  58.965000  29.445000 ;
      RECT  50.865000  29.445000  55.445000  30.045000 ;
      RECT  51.265000 -41.290000  61.275000 -40.690000 ;
      RECT  51.900000  40.055000  55.445000  43.575000 ;
      RECT  52.500000 -26.935000  58.965000 -25.900000 ;
      RECT  52.500000 -25.900000  62.510000 -25.300000 ;
      RECT  52.500000  25.300000  62.510000  25.900000 ;
      RECT  52.500000  25.900000  58.965000  26.935000 ;
      RECT  54.810000 -40.690000  61.275000 -37.145000 ;
      RECT  55.010000 -25.300000  62.510000  25.300000 ;
      RECT  57.730000 -37.145000  61.275000 -34.225000 ;
      RECT  58.990000  32.965000  66.055000  36.510000 ;
      RECT  62.510000 -30.680000  71.885000 -30.045000 ;
      RECT  62.510000 -30.045000  72.520000 -29.445000 ;
      RECT  62.510000  29.445000  72.520000  30.045000 ;
      RECT  62.510000  30.045000  66.055000  32.965000 ;
      RECT  65.020000 -29.445000  72.520000 -16.250000 ;
      RECT  65.020000 -16.250000  77.500000  -8.750000 ;
      RECT  65.020000   8.750000  77.500000  16.250000 ;
      RECT  65.020000  16.250000  72.520000  29.445000 ;
    LAYER via2 ;
      RECT -20.120000 -70.635000 -18.840000 -69.355000 ;
      RECT -20.120000 -68.165000 -18.840000 -66.885000 ;
      RECT -19.830000  56.885000 -18.550000  58.165000 ;
      RECT -19.830000  59.355000 -18.550000  60.635000 ;
      RECT -17.500000 -70.635000 -16.220000 -69.355000 ;
      RECT -17.500000 -68.165000 -16.220000 -66.885000 ;
      RECT -17.210000  56.885000 -15.930000  58.165000 ;
      RECT -17.210000  59.355000 -15.930000  60.635000 ;
      RECT -14.730000 -70.635000 -13.450000 -69.355000 ;
      RECT -14.730000 -68.165000 -13.450000 -66.885000 ;
      RECT -14.440000  56.885000 -13.160000  58.165000 ;
      RECT -14.440000  59.355000 -13.160000  60.635000 ;
      RECT -11.960000 -70.635000 -10.680000 -69.355000 ;
      RECT -11.960000 -68.165000 -10.680000 -66.885000 ;
      RECT -11.670000  56.885000 -10.390000  58.165000 ;
      RECT -11.670000  59.355000 -10.390000  60.635000 ;
      RECT  -9.340000 -70.635000  -8.060000 -69.355000 ;
      RECT  -9.340000 -68.165000  -8.060000 -66.885000 ;
      RECT  -9.050000  56.885000  -7.770000  58.165000 ;
      RECT  -9.050000  59.355000  -7.770000  60.635000 ;
      RECT   7.050000 -60.635000   8.330000 -59.355000 ;
      RECT   7.050000 -58.165000   8.330000 -56.885000 ;
      RECT   7.555000  46.870000   8.835000  48.150000 ;
      RECT   7.555000  49.340000   8.835000  50.620000 ;
      RECT   9.670000 -60.635000  10.950000 -59.355000 ;
      RECT   9.670000 -58.165000  10.950000 -56.885000 ;
      RECT  10.175000  46.870000  11.455000  48.150000 ;
      RECT  10.175000  49.340000  11.455000  50.620000 ;
      RECT  12.440000 -60.635000  13.720000 -59.355000 ;
      RECT  12.440000 -58.165000  13.720000 -56.885000 ;
      RECT  12.945000  46.870000  14.225000  48.150000 ;
      RECT  12.945000  49.340000  14.225000  50.620000 ;
      RECT  15.210000 -60.635000  16.490000 -59.355000 ;
      RECT  15.210000 -58.165000  16.490000 -56.885000 ;
      RECT  15.715000  46.870000  16.995000  48.150000 ;
      RECT  15.715000  49.340000  16.995000  50.620000 ;
      RECT  17.830000 -60.635000  19.110000 -59.355000 ;
      RECT  17.830000 -58.165000  19.110000 -56.885000 ;
      RECT  18.335000  46.870000  19.615000  48.150000 ;
      RECT  18.335000  49.340000  19.615000  50.620000 ;
      RECT  32.760000  -1.875000  34.040000  -0.595000 ;
      RECT  32.760000   0.595000  34.040000   1.875000 ;
      RECT  35.380000  -1.875000  36.660000  -0.595000 ;
      RECT  35.380000   0.595000  36.660000   1.875000 ;
      RECT  38.150000  -1.875000  39.430000  -0.595000 ;
      RECT  38.150000   0.595000  39.430000   1.875000 ;
  END
END sky130_fd_pr__rf_test_coil1
END LIBRARY
