# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4_top
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4_top ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.27000 BY  11.85000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT  0.000000  0.000000 13.270000  0.330000 ;
        RECT  0.000000  0.330000  0.330000  5.760000 ;
        RECT  0.000000  5.760000 13.270000  6.090000 ;
        RECT  0.000000  6.090000  0.330000 11.520000 ;
        RECT  0.000000 11.520000 13.270000 11.850000 ;
        RECT  1.270000  0.330000  1.610000  2.580000 ;
        RECT  1.270000  3.510000  1.610000  5.760000 ;
        RECT  1.270000  6.090000  1.610000  8.340000 ;
        RECT  1.270000  9.270000  1.610000 11.520000 ;
        RECT  2.550000  0.330000  2.890000  2.580000 ;
        RECT  2.550000  3.510000  2.890000  5.760000 ;
        RECT  2.550000  6.090000  2.890000  8.340000 ;
        RECT  2.550000  9.270000  2.890000 11.520000 ;
        RECT  3.910000  0.330000  4.250000  2.580000 ;
        RECT  3.910000  3.510000  4.250000  5.760000 ;
        RECT  3.910000  6.090000  4.250000  8.340000 ;
        RECT  3.910000  9.270000  4.250000 11.520000 ;
        RECT  5.190000  0.330000  5.530000  2.580000 ;
        RECT  5.190000  3.510000  5.530000  5.760000 ;
        RECT  5.190000  6.090000  5.530000  8.340000 ;
        RECT  5.190000  9.270000  5.530000 11.520000 ;
        RECT  6.470000  0.330000  6.800000  5.760000 ;
        RECT  6.470000  6.090000  6.800000 11.520000 ;
        RECT  7.740000  0.330000  8.080000  2.580000 ;
        RECT  7.740000  3.510000  8.080000  5.760000 ;
        RECT  7.740000  6.090000  8.080000  8.340000 ;
        RECT  7.740000  9.270000  8.080000 11.520000 ;
        RECT  9.020000  0.330000  9.360000  2.580000 ;
        RECT  9.020000  3.510000  9.360000  5.760000 ;
        RECT  9.020000  6.090000  9.360000  8.340000 ;
        RECT  9.020000  9.270000  9.360000 11.520000 ;
        RECT 10.380000  0.330000 10.720000  2.580000 ;
        RECT 10.380000  3.510000 10.720000  5.760000 ;
        RECT 10.380000  6.090000 10.720000  8.340000 ;
        RECT 10.380000  9.270000 10.720000 11.520000 ;
        RECT 11.660000  0.330000 12.000000  2.580000 ;
        RECT 11.660000  3.510000 12.000000  5.760000 ;
        RECT 11.660000  6.090000 12.000000  8.340000 ;
        RECT 11.660000  9.270000 12.000000 11.520000 ;
        RECT 12.940000  0.330000 13.270000  5.760000 ;
        RECT 12.940000  6.090000 13.270000 11.520000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT  0.630000 0.630000  0.970000  2.880000 ;
        RECT  0.630000 2.880000  6.170000  3.210000 ;
        RECT  0.630000 3.210000  0.970000  5.460000 ;
        RECT  0.630000 6.390000  0.970000  8.640000 ;
        RECT  0.630000 8.640000  6.170000  8.970000 ;
        RECT  0.630000 8.970000  0.970000 11.220000 ;
        RECT  1.910000 0.630000  2.250000  2.880000 ;
        RECT  1.910000 3.210000  2.250000  5.460000 ;
        RECT  1.910000 6.390000  2.250000  8.640000 ;
        RECT  1.910000 8.970000  2.250000 11.220000 ;
        RECT  3.190000 0.630000  3.610000  2.880000 ;
        RECT  3.190000 3.210000  3.610000  5.460000 ;
        RECT  3.190000 6.390000  3.610000  8.640000 ;
        RECT  3.190000 8.970000  3.610000 11.220000 ;
        RECT  4.550000 0.630000  4.890000  2.880000 ;
        RECT  4.550000 3.210000  4.890000  5.460000 ;
        RECT  4.550000 6.390000  4.890000  8.640000 ;
        RECT  4.550000 8.970000  4.890000 11.220000 ;
        RECT  5.830000 0.630000  6.170000  2.880000 ;
        RECT  5.830000 3.210000  6.170000  5.460000 ;
        RECT  5.830000 6.390000  6.170000  8.640000 ;
        RECT  5.830000 8.970000  6.170000 11.220000 ;
        RECT  7.100000 0.630000  7.440000  2.880000 ;
        RECT  7.100000 2.880000 12.640000  3.210000 ;
        RECT  7.100000 3.210000  7.440000  5.460000 ;
        RECT  7.100000 6.390000  7.440000  8.640000 ;
        RECT  7.100000 8.640000 12.640000  8.970000 ;
        RECT  7.100000 8.970000  7.440000 11.220000 ;
        RECT  8.380000 0.630000  8.720000  2.880000 ;
        RECT  8.380000 3.210000  8.720000  5.460000 ;
        RECT  8.380000 6.390000  8.720000  8.640000 ;
        RECT  8.380000 8.970000  8.720000 11.220000 ;
        RECT  9.660000 0.630000 10.080000  2.880000 ;
        RECT  9.660000 3.210000 10.080000  5.460000 ;
        RECT  9.660000 6.390000 10.080000  8.640000 ;
        RECT  9.660000 8.970000 10.080000 11.220000 ;
        RECT 11.020000 0.630000 11.360000  2.880000 ;
        RECT 11.020000 3.210000 11.360000  5.460000 ;
        RECT 11.020000 6.390000 11.360000  8.640000 ;
        RECT 11.020000 8.970000 11.360000 11.220000 ;
        RECT 12.300000 0.630000 12.640000  2.880000 ;
        RECT 12.300000 3.210000 12.640000  5.460000 ;
        RECT 12.300000 6.390000 12.640000  8.640000 ;
        RECT 12.300000 8.970000 12.640000 11.220000 ;
    END
  END C1
  PIN M4
    PORT
      LAYER met4 ;
        RECT 0.000000 0.000000 13.270000 11.850000 ;
    END
  END M4
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 5.895000 6.345000 5.945000 6.395000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT  0.000000  0.000000 13.270000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.860000 ;
      RECT  0.000000  0.860000  3.055000  1.030000 ;
      RECT  0.000000  1.030000  0.330000  1.560000 ;
      RECT  0.000000  1.560000  3.055000  1.730000 ;
      RECT  0.000000  1.730000  0.330000  2.260000 ;
      RECT  0.000000  2.260000  3.055000  2.430000 ;
      RECT  0.000000  2.430000  0.330000  2.960000 ;
      RECT  0.000000  2.960000  3.055000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.660000 ;
      RECT  0.000000  3.660000  3.055000  3.830000 ;
      RECT  0.000000  3.830000  0.330000  4.360000 ;
      RECT  0.000000  4.360000  3.055000  4.530000 ;
      RECT  0.000000  4.530000  0.330000  5.060000 ;
      RECT  0.000000  5.060000  3.055000  5.230000 ;
      RECT  0.000000  5.230000  0.330000  5.760000 ;
      RECT  0.000000  5.760000 13.270000  6.090000 ;
      RECT  0.000000  6.090000  0.330000  6.620000 ;
      RECT  0.000000  6.620000  3.055000  6.790000 ;
      RECT  0.000000  6.790000  0.330000  7.320000 ;
      RECT  0.000000  7.320000  3.055000  7.490000 ;
      RECT  0.000000  7.490000  0.330000  8.020000 ;
      RECT  0.000000  8.020000  3.055000  8.190000 ;
      RECT  0.000000  8.190000  0.330000  8.720000 ;
      RECT  0.000000  8.720000  3.055000  8.890000 ;
      RECT  0.000000  8.890000  0.330000  9.420000 ;
      RECT  0.000000  9.420000  3.055000  9.590000 ;
      RECT  0.000000  9.590000  0.330000 10.120000 ;
      RECT  0.000000 10.120000  3.055000 10.290000 ;
      RECT  0.000000 10.290000  0.330000 10.820000 ;
      RECT  0.000000 10.820000  3.055000 10.990000 ;
      RECT  0.000000 10.990000  0.330000 11.520000 ;
      RECT  0.000000 11.520000 13.270000 11.850000 ;
      RECT  0.500000  0.500000  6.300000  0.690000 ;
      RECT  0.500000  1.200000  6.300000  1.390000 ;
      RECT  0.500000  1.900000  6.300000  2.090000 ;
      RECT  0.500000  2.600000  6.300000  2.790000 ;
      RECT  0.500000  3.300000  6.300000  3.490000 ;
      RECT  0.500000  4.000000  6.300000  4.190000 ;
      RECT  0.500000  4.700000  6.300000  4.890000 ;
      RECT  0.500000  5.400000  6.300000  5.590000 ;
      RECT  0.500000  6.260000  6.300000  6.450000 ;
      RECT  0.500000  6.960000  6.300000  7.150000 ;
      RECT  0.500000  7.660000  6.300000  7.850000 ;
      RECT  0.500000  8.360000  6.300000  8.550000 ;
      RECT  0.500000  9.060000  6.300000  9.250000 ;
      RECT  0.500000  9.760000  6.300000  9.950000 ;
      RECT  0.500000 10.460000  6.300000 10.650000 ;
      RECT  0.500000 11.160000  6.300000 11.350000 ;
      RECT  3.240000  0.690000  3.560000  1.200000 ;
      RECT  3.240000  1.390000  3.560000  1.900000 ;
      RECT  3.240000  2.090000  3.560000  2.600000 ;
      RECT  3.240000  2.790000  3.560000  3.300000 ;
      RECT  3.240000  3.490000  3.560000  4.000000 ;
      RECT  3.240000  4.190000  3.560000  4.700000 ;
      RECT  3.240000  4.890000  3.560000  5.400000 ;
      RECT  3.240000  6.450000  3.560000  6.960000 ;
      RECT  3.240000  7.150000  3.560000  7.660000 ;
      RECT  3.240000  7.850000  3.560000  8.360000 ;
      RECT  3.240000  8.550000  3.560000  9.060000 ;
      RECT  3.240000  9.250000  3.560000  9.760000 ;
      RECT  3.240000  9.950000  3.560000 10.460000 ;
      RECT  3.240000 10.650000  3.560000 11.160000 ;
      RECT  3.730000  0.860000  9.525000  1.030000 ;
      RECT  3.730000  1.560000  9.525000  1.730000 ;
      RECT  3.730000  2.260000  9.525000  2.430000 ;
      RECT  3.730000  2.960000  9.525000  3.130000 ;
      RECT  3.730000  3.660000  9.525000  3.830000 ;
      RECT  3.730000  4.360000  9.525000  4.530000 ;
      RECT  3.730000  5.060000  9.525000  5.230000 ;
      RECT  3.730000  6.620000  9.525000  6.790000 ;
      RECT  3.730000  7.320000  9.525000  7.490000 ;
      RECT  3.730000  8.020000  9.525000  8.190000 ;
      RECT  3.730000  8.720000  9.525000  8.890000 ;
      RECT  3.730000  9.420000  9.525000  9.590000 ;
      RECT  3.730000 10.120000  9.525000 10.290000 ;
      RECT  3.730000 10.820000  9.525000 10.990000 ;
      RECT  6.470000  0.330000  6.800000  0.860000 ;
      RECT  6.470000  1.030000  6.800000  1.560000 ;
      RECT  6.470000  1.730000  6.800000  2.260000 ;
      RECT  6.470000  2.430000  6.800000  2.960000 ;
      RECT  6.470000  3.130000  6.800000  3.660000 ;
      RECT  6.470000  3.830000  6.800000  4.360000 ;
      RECT  6.470000  4.530000  6.800000  5.060000 ;
      RECT  6.470000  5.230000  6.800000  5.760000 ;
      RECT  6.470000  6.090000  6.800000  6.620000 ;
      RECT  6.470000  6.790000  6.800000  7.320000 ;
      RECT  6.470000  7.490000  6.800000  8.020000 ;
      RECT  6.470000  8.190000  6.800000  8.720000 ;
      RECT  6.470000  8.890000  6.800000  9.420000 ;
      RECT  6.470000  9.590000  6.800000 10.120000 ;
      RECT  6.470000 10.290000  6.800000 10.820000 ;
      RECT  6.470000 10.990000  6.800000 11.520000 ;
      RECT  6.970000  0.500000 12.770000  0.690000 ;
      RECT  6.970000  1.200000 12.770000  1.390000 ;
      RECT  6.970000  1.900000 12.770000  2.090000 ;
      RECT  6.970000  2.600000 12.770000  2.790000 ;
      RECT  6.970000  3.300000 12.770000  3.490000 ;
      RECT  6.970000  4.000000 12.770000  4.190000 ;
      RECT  6.970000  4.700000 12.770000  4.890000 ;
      RECT  6.970000  5.400000 12.770000  5.590000 ;
      RECT  6.970000  6.260000 12.770000  6.450000 ;
      RECT  6.970000  6.960000 12.770000  7.150000 ;
      RECT  6.970000  7.660000 12.770000  7.850000 ;
      RECT  6.970000  8.360000 12.770000  8.550000 ;
      RECT  6.970000  9.060000 12.770000  9.250000 ;
      RECT  6.970000  9.760000 12.770000  9.950000 ;
      RECT  6.970000 10.460000 12.770000 10.650000 ;
      RECT  6.970000 11.160000 12.770000 11.350000 ;
      RECT  9.710000  0.690000 10.030000  1.200000 ;
      RECT  9.710000  1.390000 10.030000  1.900000 ;
      RECT  9.710000  2.090000 10.030000  2.600000 ;
      RECT  9.710000  2.790000 10.030000  3.300000 ;
      RECT  9.710000  3.490000 10.030000  4.000000 ;
      RECT  9.710000  4.190000 10.030000  4.700000 ;
      RECT  9.710000  4.890000 10.030000  5.400000 ;
      RECT  9.710000  6.450000 10.030000  6.960000 ;
      RECT  9.710000  7.150000 10.030000  7.660000 ;
      RECT  9.710000  7.850000 10.030000  8.360000 ;
      RECT  9.710000  8.550000 10.030000  9.060000 ;
      RECT  9.710000  9.250000 10.030000  9.760000 ;
      RECT  9.710000  9.950000 10.030000 10.460000 ;
      RECT  9.710000 10.650000 10.030000 11.160000 ;
      RECT 10.200000  0.860000 13.270000  1.030000 ;
      RECT 10.200000  1.560000 13.270000  1.730000 ;
      RECT 10.200000  2.260000 13.270000  2.430000 ;
      RECT 10.200000  2.960000 13.270000  3.130000 ;
      RECT 10.200000  3.660000 13.270000  3.830000 ;
      RECT 10.200000  4.360000 13.270000  4.530000 ;
      RECT 10.200000  5.060000 13.270000  5.230000 ;
      RECT 10.200000  6.620000 13.270000  6.790000 ;
      RECT 10.200000  7.320000 13.270000  7.490000 ;
      RECT 10.200000  8.020000 13.270000  8.190000 ;
      RECT 10.200000  8.720000 13.270000  8.890000 ;
      RECT 10.200000  9.420000 13.270000  9.590000 ;
      RECT 10.200000 10.120000 13.270000 10.290000 ;
      RECT 10.200000 10.820000 13.270000 10.990000 ;
      RECT 12.940000  0.330000 13.270000  0.860000 ;
      RECT 12.940000  1.030000 13.270000  1.560000 ;
      RECT 12.940000  1.730000 13.270000  2.260000 ;
      RECT 12.940000  2.430000 13.270000  2.960000 ;
      RECT 12.940000  3.130000 13.270000  3.660000 ;
      RECT 12.940000  3.830000 13.270000  4.360000 ;
      RECT 12.940000  4.530000 13.270000  5.060000 ;
      RECT 12.940000  5.230000 13.270000  5.760000 ;
      RECT 12.940000  6.090000 13.270000  6.620000 ;
      RECT 12.940000  6.790000 13.270000  7.320000 ;
      RECT 12.940000  7.490000 13.270000  8.020000 ;
      RECT 12.940000  8.190000 13.270000  8.720000 ;
      RECT 12.940000  8.890000 13.270000  9.420000 ;
      RECT 12.940000  9.590000 13.270000 10.120000 ;
      RECT 12.940000 10.290000 13.270000 10.820000 ;
      RECT 12.940000 10.990000 13.270000 11.520000 ;
    LAYER mcon ;
      RECT  0.080000  0.440000  0.250000  0.610000 ;
      RECT  0.080000  0.800000  0.250000  0.970000 ;
      RECT  0.080000  1.160000  0.250000  1.330000 ;
      RECT  0.080000  1.520000  0.250000  1.690000 ;
      RECT  0.080000  1.880000  0.250000  2.050000 ;
      RECT  0.080000  2.240000  0.250000  2.410000 ;
      RECT  0.080000  2.600000  0.250000  2.770000 ;
      RECT  0.080000  2.960000  0.250000  3.130000 ;
      RECT  0.080000  3.320000  0.250000  3.490000 ;
      RECT  0.080000  3.680000  0.250000  3.850000 ;
      RECT  0.080000  4.040000  0.250000  4.210000 ;
      RECT  0.080000  4.400000  0.250000  4.570000 ;
      RECT  0.080000  4.760000  0.250000  4.930000 ;
      RECT  0.080000  5.120000  0.250000  5.290000 ;
      RECT  0.080000  5.480000  0.250000  5.650000 ;
      RECT  0.080000  6.200000  0.250000  6.370000 ;
      RECT  0.080000  6.560000  0.250000  6.730000 ;
      RECT  0.080000  6.920000  0.250000  7.090000 ;
      RECT  0.080000  7.280000  0.250000  7.450000 ;
      RECT  0.080000  7.640000  0.250000  7.810000 ;
      RECT  0.080000  8.000000  0.250000  8.170000 ;
      RECT  0.080000  8.360000  0.250000  8.530000 ;
      RECT  0.080000  8.720000  0.250000  8.890000 ;
      RECT  0.080000  9.080000  0.250000  9.250000 ;
      RECT  0.080000  9.440000  0.250000  9.610000 ;
      RECT  0.080000  9.800000  0.250000  9.970000 ;
      RECT  0.080000 10.160000  0.250000 10.330000 ;
      RECT  0.080000 10.520000  0.250000 10.690000 ;
      RECT  0.080000 10.880000  0.250000 11.050000 ;
      RECT  0.080000 11.240000  0.250000 11.410000 ;
      RECT  0.410000  0.080000  0.580000  0.250000 ;
      RECT  0.410000  5.840000  0.580000  6.010000 ;
      RECT  0.410000 11.600000  0.580000 11.770000 ;
      RECT  0.770000  0.080000  0.940000  0.250000 ;
      RECT  0.770000  5.840000  0.940000  6.010000 ;
      RECT  0.770000 11.600000  0.940000 11.770000 ;
      RECT  1.130000  0.080000  1.300000  0.250000 ;
      RECT  1.130000  5.840000  1.300000  6.010000 ;
      RECT  1.130000 11.600000  1.300000 11.770000 ;
      RECT  1.490000  0.080000  1.660000  0.250000 ;
      RECT  1.490000  5.840000  1.660000  6.010000 ;
      RECT  1.490000 11.600000  1.660000 11.770000 ;
      RECT  1.850000  0.080000  2.020000  0.250000 ;
      RECT  1.850000  5.840000  2.020000  6.010000 ;
      RECT  1.850000 11.600000  2.020000 11.770000 ;
      RECT  2.210000  0.080000  2.380000  0.250000 ;
      RECT  2.210000  5.840000  2.380000  6.010000 ;
      RECT  2.210000 11.600000  2.380000 11.770000 ;
      RECT  2.570000  0.080000  2.740000  0.250000 ;
      RECT  2.570000  5.840000  2.740000  6.010000 ;
      RECT  2.570000 11.600000  2.740000 11.770000 ;
      RECT  2.930000  0.080000  3.100000  0.250000 ;
      RECT  2.930000  5.840000  3.100000  6.010000 ;
      RECT  2.930000 11.600000  3.100000 11.770000 ;
      RECT  3.315000  0.080000  3.485000  0.250000 ;
      RECT  3.315000  0.800000  3.485000  0.970000 ;
      RECT  3.315000  1.160000  3.485000  1.330000 ;
      RECT  3.315000  1.520000  3.485000  1.690000 ;
      RECT  3.315000  1.880000  3.485000  2.050000 ;
      RECT  3.315000  2.240000  3.485000  2.410000 ;
      RECT  3.315000  2.600000  3.485000  2.770000 ;
      RECT  3.315000  2.960000  3.485000  3.130000 ;
      RECT  3.315000  3.320000  3.485000  3.490000 ;
      RECT  3.315000  3.680000  3.485000  3.850000 ;
      RECT  3.315000  4.040000  3.485000  4.210000 ;
      RECT  3.315000  4.400000  3.485000  4.570000 ;
      RECT  3.315000  4.760000  3.485000  4.930000 ;
      RECT  3.315000  5.120000  3.485000  5.290000 ;
      RECT  3.315000  5.840000  3.485000  6.010000 ;
      RECT  3.315000  6.560000  3.485000  6.730000 ;
      RECT  3.315000  6.920000  3.485000  7.090000 ;
      RECT  3.315000  7.280000  3.485000  7.450000 ;
      RECT  3.315000  7.640000  3.485000  7.810000 ;
      RECT  3.315000  8.000000  3.485000  8.170000 ;
      RECT  3.315000  8.360000  3.485000  8.530000 ;
      RECT  3.315000  8.720000  3.485000  8.890000 ;
      RECT  3.315000  9.080000  3.485000  9.250000 ;
      RECT  3.315000  9.440000  3.485000  9.610000 ;
      RECT  3.315000  9.800000  3.485000  9.970000 ;
      RECT  3.315000 10.160000  3.485000 10.330000 ;
      RECT  3.315000 10.520000  3.485000 10.690000 ;
      RECT  3.315000 10.880000  3.485000 11.050000 ;
      RECT  3.315000 11.600000  3.485000 11.770000 ;
      RECT  3.700000  0.080000  3.870000  0.250000 ;
      RECT  3.700000  5.840000  3.870000  6.010000 ;
      RECT  3.700000 11.600000  3.870000 11.770000 ;
      RECT  4.060000  0.080000  4.230000  0.250000 ;
      RECT  4.060000  5.840000  4.230000  6.010000 ;
      RECT  4.060000 11.600000  4.230000 11.770000 ;
      RECT  4.420000  0.080000  4.590000  0.250000 ;
      RECT  4.420000  5.840000  4.590000  6.010000 ;
      RECT  4.420000 11.600000  4.590000 11.770000 ;
      RECT  4.780000  0.080000  4.950000  0.250000 ;
      RECT  4.780000  5.840000  4.950000  6.010000 ;
      RECT  4.780000 11.600000  4.950000 11.770000 ;
      RECT  5.140000  0.080000  5.310000  0.250000 ;
      RECT  5.140000  5.840000  5.310000  6.010000 ;
      RECT  5.140000 11.600000  5.310000 11.770000 ;
      RECT  5.500000  0.080000  5.670000  0.250000 ;
      RECT  5.500000  5.840000  5.670000  6.010000 ;
      RECT  5.500000 11.600000  5.670000 11.770000 ;
      RECT  5.860000  0.080000  6.030000  0.250000 ;
      RECT  5.860000  5.840000  6.030000  6.010000 ;
      RECT  5.860000 11.600000  6.030000 11.770000 ;
      RECT  6.220000  0.080000  6.390000  0.250000 ;
      RECT  6.220000  5.840000  6.390000  6.010000 ;
      RECT  6.220000 11.600000  6.390000 11.770000 ;
      RECT  6.550000  0.440000  6.720000  0.610000 ;
      RECT  6.550000  0.800000  6.720000  0.970000 ;
      RECT  6.550000  1.160000  6.720000  1.330000 ;
      RECT  6.550000  1.520000  6.720000  1.690000 ;
      RECT  6.550000  1.880000  6.720000  2.050000 ;
      RECT  6.550000  2.240000  6.720000  2.410000 ;
      RECT  6.550000  2.600000  6.720000  2.770000 ;
      RECT  6.550000  2.960000  6.720000  3.130000 ;
      RECT  6.550000  3.320000  6.720000  3.490000 ;
      RECT  6.550000  3.680000  6.720000  3.850000 ;
      RECT  6.550000  4.040000  6.720000  4.210000 ;
      RECT  6.550000  4.400000  6.720000  4.570000 ;
      RECT  6.550000  4.760000  6.720000  4.930000 ;
      RECT  6.550000  5.120000  6.720000  5.290000 ;
      RECT  6.550000  5.480000  6.720000  5.650000 ;
      RECT  6.550000  6.200000  6.720000  6.370000 ;
      RECT  6.550000  6.560000  6.720000  6.730000 ;
      RECT  6.550000  6.920000  6.720000  7.090000 ;
      RECT  6.550000  7.280000  6.720000  7.450000 ;
      RECT  6.550000  7.640000  6.720000  7.810000 ;
      RECT  6.550000  8.000000  6.720000  8.170000 ;
      RECT  6.550000  8.360000  6.720000  8.530000 ;
      RECT  6.550000  8.720000  6.720000  8.890000 ;
      RECT  6.550000  9.080000  6.720000  9.250000 ;
      RECT  6.550000  9.440000  6.720000  9.610000 ;
      RECT  6.550000  9.800000  6.720000  9.970000 ;
      RECT  6.550000 10.160000  6.720000 10.330000 ;
      RECT  6.550000 10.520000  6.720000 10.690000 ;
      RECT  6.550000 10.880000  6.720000 11.050000 ;
      RECT  6.550000 11.240000  6.720000 11.410000 ;
      RECT  6.880000  0.080000  7.050000  0.250000 ;
      RECT  6.880000  5.840000  7.050000  6.010000 ;
      RECT  6.880000 11.600000  7.050000 11.770000 ;
      RECT  7.240000  0.080000  7.410000  0.250000 ;
      RECT  7.240000  5.840000  7.410000  6.010000 ;
      RECT  7.240000 11.600000  7.410000 11.770000 ;
      RECT  7.600000  0.080000  7.770000  0.250000 ;
      RECT  7.600000  5.840000  7.770000  6.010000 ;
      RECT  7.600000 11.600000  7.770000 11.770000 ;
      RECT  7.960000  0.080000  8.130000  0.250000 ;
      RECT  7.960000  5.840000  8.130000  6.010000 ;
      RECT  7.960000 11.600000  8.130000 11.770000 ;
      RECT  8.320000  0.080000  8.490000  0.250000 ;
      RECT  8.320000  5.840000  8.490000  6.010000 ;
      RECT  8.320000 11.600000  8.490000 11.770000 ;
      RECT  8.680000  0.080000  8.850000  0.250000 ;
      RECT  8.680000  5.840000  8.850000  6.010000 ;
      RECT  8.680000 11.600000  8.850000 11.770000 ;
      RECT  9.040000  0.080000  9.210000  0.250000 ;
      RECT  9.040000  5.840000  9.210000  6.010000 ;
      RECT  9.040000 11.600000  9.210000 11.770000 ;
      RECT  9.400000  0.080000  9.570000  0.250000 ;
      RECT  9.400000  5.840000  9.570000  6.010000 ;
      RECT  9.400000 11.600000  9.570000 11.770000 ;
      RECT  9.785000  0.080000  9.955000  0.250000 ;
      RECT  9.785000  0.800000  9.955000  0.970000 ;
      RECT  9.785000  1.160000  9.955000  1.330000 ;
      RECT  9.785000  1.520000  9.955000  1.690000 ;
      RECT  9.785000  1.880000  9.955000  2.050000 ;
      RECT  9.785000  2.240000  9.955000  2.410000 ;
      RECT  9.785000  2.600000  9.955000  2.770000 ;
      RECT  9.785000  2.960000  9.955000  3.130000 ;
      RECT  9.785000  3.320000  9.955000  3.490000 ;
      RECT  9.785000  3.680000  9.955000  3.850000 ;
      RECT  9.785000  4.040000  9.955000  4.210000 ;
      RECT  9.785000  4.400000  9.955000  4.570000 ;
      RECT  9.785000  4.760000  9.955000  4.930000 ;
      RECT  9.785000  5.120000  9.955000  5.290000 ;
      RECT  9.785000  5.840000  9.955000  6.010000 ;
      RECT  9.785000  6.560000  9.955000  6.730000 ;
      RECT  9.785000  6.920000  9.955000  7.090000 ;
      RECT  9.785000  7.280000  9.955000  7.450000 ;
      RECT  9.785000  7.640000  9.955000  7.810000 ;
      RECT  9.785000  8.000000  9.955000  8.170000 ;
      RECT  9.785000  8.360000  9.955000  8.530000 ;
      RECT  9.785000  8.720000  9.955000  8.890000 ;
      RECT  9.785000  9.080000  9.955000  9.250000 ;
      RECT  9.785000  9.440000  9.955000  9.610000 ;
      RECT  9.785000  9.800000  9.955000  9.970000 ;
      RECT  9.785000 10.160000  9.955000 10.330000 ;
      RECT  9.785000 10.520000  9.955000 10.690000 ;
      RECT  9.785000 10.880000  9.955000 11.050000 ;
      RECT  9.785000 11.600000  9.955000 11.770000 ;
      RECT 10.170000  0.080000 10.340000  0.250000 ;
      RECT 10.170000  5.840000 10.340000  6.010000 ;
      RECT 10.170000 11.600000 10.340000 11.770000 ;
      RECT 10.530000  0.080000 10.700000  0.250000 ;
      RECT 10.530000  5.840000 10.700000  6.010000 ;
      RECT 10.530000 11.600000 10.700000 11.770000 ;
      RECT 10.890000  0.080000 11.060000  0.250000 ;
      RECT 10.890000  5.840000 11.060000  6.010000 ;
      RECT 10.890000 11.600000 11.060000 11.770000 ;
      RECT 11.250000  0.080000 11.420000  0.250000 ;
      RECT 11.250000  5.840000 11.420000  6.010000 ;
      RECT 11.250000 11.600000 11.420000 11.770000 ;
      RECT 11.610000  0.080000 11.780000  0.250000 ;
      RECT 11.610000  5.840000 11.780000  6.010000 ;
      RECT 11.610000 11.600000 11.780000 11.770000 ;
      RECT 11.970000  0.080000 12.140000  0.250000 ;
      RECT 11.970000  5.840000 12.140000  6.010000 ;
      RECT 11.970000 11.600000 12.140000 11.770000 ;
      RECT 12.330000  0.080000 12.500000  0.250000 ;
      RECT 12.330000  5.840000 12.500000  6.010000 ;
      RECT 12.330000 11.600000 12.500000 11.770000 ;
      RECT 12.690000  0.080000 12.860000  0.250000 ;
      RECT 12.690000  5.840000 12.860000  6.010000 ;
      RECT 12.690000 11.600000 12.860000 11.770000 ;
      RECT 13.020000  0.440000 13.190000  0.610000 ;
      RECT 13.020000  0.800000 13.190000  0.970000 ;
      RECT 13.020000  1.160000 13.190000  1.330000 ;
      RECT 13.020000  1.520000 13.190000  1.690000 ;
      RECT 13.020000  1.880000 13.190000  2.050000 ;
      RECT 13.020000  2.240000 13.190000  2.410000 ;
      RECT 13.020000  2.600000 13.190000  2.770000 ;
      RECT 13.020000  2.960000 13.190000  3.130000 ;
      RECT 13.020000  3.320000 13.190000  3.490000 ;
      RECT 13.020000  3.680000 13.190000  3.850000 ;
      RECT 13.020000  4.040000 13.190000  4.210000 ;
      RECT 13.020000  4.400000 13.190000  4.570000 ;
      RECT 13.020000  4.760000 13.190000  4.930000 ;
      RECT 13.020000  5.120000 13.190000  5.290000 ;
      RECT 13.020000  5.480000 13.190000  5.650000 ;
      RECT 13.020000  6.200000 13.190000  6.370000 ;
      RECT 13.020000  6.560000 13.190000  6.730000 ;
      RECT 13.020000  6.920000 13.190000  7.090000 ;
      RECT 13.020000  7.280000 13.190000  7.450000 ;
      RECT 13.020000  7.640000 13.190000  7.810000 ;
      RECT 13.020000  8.000000 13.190000  8.170000 ;
      RECT 13.020000  8.360000 13.190000  8.530000 ;
      RECT 13.020000  8.720000 13.190000  8.890000 ;
      RECT 13.020000  9.080000 13.190000  9.250000 ;
      RECT 13.020000  9.440000 13.190000  9.610000 ;
      RECT 13.020000  9.800000 13.190000  9.970000 ;
      RECT 13.020000 10.160000 13.190000 10.330000 ;
      RECT 13.020000 10.520000 13.190000 10.690000 ;
      RECT 13.020000 10.880000 13.190000 11.050000 ;
      RECT 13.020000 11.240000 13.190000 11.410000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 13.270000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  5.760000 ;
      RECT  0.000000  5.760000 13.270000  6.090000 ;
      RECT  0.000000  6.090000  0.330000 11.520000 ;
      RECT  0.000000 11.520000 13.270000 11.850000 ;
      RECT  0.470000  0.470000  0.610000  2.885000 ;
      RECT  0.470000  2.885000  6.330000  3.205000 ;
      RECT  0.470000  3.205000  0.610000  5.620000 ;
      RECT  0.470000  6.230000  0.610000  8.645000 ;
      RECT  0.470000  8.645000  6.330000  8.965000 ;
      RECT  0.470000  8.965000  0.610000 11.380000 ;
      RECT  0.750000  0.330000  0.890000  2.745000 ;
      RECT  0.750000  3.345000  0.890000  5.760000 ;
      RECT  0.750000  6.090000  0.890000  8.505000 ;
      RECT  0.750000  9.105000  0.890000 11.520000 ;
      RECT  1.030000  0.470000  1.170000  2.885000 ;
      RECT  1.030000  3.205000  1.170000  5.620000 ;
      RECT  1.030000  6.230000  1.170000  8.645000 ;
      RECT  1.030000  8.965000  1.170000 11.380000 ;
      RECT  1.310000  0.330000  1.450000  2.745000 ;
      RECT  1.310000  3.345000  1.450000  5.760000 ;
      RECT  1.310000  6.090000  1.450000  8.505000 ;
      RECT  1.310000  9.105000  1.450000 11.520000 ;
      RECT  1.590000  0.470000  1.730000  2.885000 ;
      RECT  1.590000  3.205000  1.730000  5.620000 ;
      RECT  1.590000  6.230000  1.730000  8.645000 ;
      RECT  1.590000  8.965000  1.730000 11.380000 ;
      RECT  1.870000  0.330000  2.010000  2.745000 ;
      RECT  1.870000  3.345000  2.010000  5.760000 ;
      RECT  1.870000  6.090000  2.010000  8.505000 ;
      RECT  1.870000  9.105000  2.010000 11.520000 ;
      RECT  2.150000  0.470000  2.290000  2.885000 ;
      RECT  2.150000  3.205000  2.290000  5.620000 ;
      RECT  2.150000  6.230000  2.290000  8.645000 ;
      RECT  2.150000  8.965000  2.290000 11.380000 ;
      RECT  2.430000  0.330000  2.570000  2.745000 ;
      RECT  2.430000  3.345000  2.570000  5.760000 ;
      RECT  2.430000  6.090000  2.570000  8.505000 ;
      RECT  2.430000  9.105000  2.570000 11.520000 ;
      RECT  2.710000  0.470000  2.850000  2.885000 ;
      RECT  2.710000  3.205000  2.850000  5.620000 ;
      RECT  2.710000  6.230000  2.850000  8.645000 ;
      RECT  2.710000  8.965000  2.850000 11.380000 ;
      RECT  2.990000  0.330000  3.130000  2.745000 ;
      RECT  2.990000  3.345000  3.130000  5.760000 ;
      RECT  2.990000  6.090000  3.130000  8.505000 ;
      RECT  2.990000  9.105000  3.130000 11.520000 ;
      RECT  3.270000  0.470000  3.530000  2.885000 ;
      RECT  3.270000  3.205000  3.530000  5.620000 ;
      RECT  3.270000  6.230000  3.530000  8.645000 ;
      RECT  3.270000  8.965000  3.530000 11.380000 ;
      RECT  3.670000  0.330000  3.810000  2.745000 ;
      RECT  3.670000  3.345000  3.810000  5.760000 ;
      RECT  3.670000  6.090000  3.810000  8.505000 ;
      RECT  3.670000  9.105000  3.810000 11.520000 ;
      RECT  3.950000  0.470000  4.090000  2.885000 ;
      RECT  3.950000  3.205000  4.090000  5.620000 ;
      RECT  3.950000  6.230000  4.090000  8.645000 ;
      RECT  3.950000  8.965000  4.090000 11.380000 ;
      RECT  4.230000  0.330000  4.370000  2.745000 ;
      RECT  4.230000  3.345000  4.370000  5.760000 ;
      RECT  4.230000  6.090000  4.370000  8.505000 ;
      RECT  4.230000  9.105000  4.370000 11.520000 ;
      RECT  4.510000  0.470000  4.650000  2.885000 ;
      RECT  4.510000  3.205000  4.650000  5.620000 ;
      RECT  4.510000  6.230000  4.650000  8.645000 ;
      RECT  4.510000  8.965000  4.650000 11.380000 ;
      RECT  4.790000  0.330000  4.930000  2.745000 ;
      RECT  4.790000  3.345000  4.930000  5.760000 ;
      RECT  4.790000  6.090000  4.930000  8.505000 ;
      RECT  4.790000  9.105000  4.930000 11.520000 ;
      RECT  5.070000  0.470000  5.210000  2.885000 ;
      RECT  5.070000  3.205000  5.210000  5.620000 ;
      RECT  5.070000  6.230000  5.210000  8.645000 ;
      RECT  5.070000  8.965000  5.210000 11.380000 ;
      RECT  5.350000  0.330000  5.490000  2.745000 ;
      RECT  5.350000  3.345000  5.490000  5.760000 ;
      RECT  5.350000  6.090000  5.490000  8.505000 ;
      RECT  5.350000  9.105000  5.490000 11.520000 ;
      RECT  5.630000  0.470000  5.770000  2.885000 ;
      RECT  5.630000  3.205000  5.770000  5.620000 ;
      RECT  5.630000  6.230000  5.770000  8.645000 ;
      RECT  5.630000  8.965000  5.770000 11.380000 ;
      RECT  5.910000  0.330000  6.050000  2.745000 ;
      RECT  5.910000  3.345000  6.050000  5.760000 ;
      RECT  5.910000  6.090000  6.050000  8.505000 ;
      RECT  5.910000  9.105000  6.050000 11.520000 ;
      RECT  6.190000  0.470000  6.330000  2.885000 ;
      RECT  6.190000  3.205000  6.330000  5.620000 ;
      RECT  6.190000  6.230000  6.330000  8.645000 ;
      RECT  6.190000  8.965000  6.330000 11.380000 ;
      RECT  6.470000  0.330000  6.800000  5.760000 ;
      RECT  6.470000  6.090000  6.800000 11.520000 ;
      RECT  6.940000  0.470000  7.080000  2.885000 ;
      RECT  6.940000  2.885000 12.800000  3.205000 ;
      RECT  6.940000  3.205000  7.080000  5.620000 ;
      RECT  6.940000  6.230000  7.080000  8.645000 ;
      RECT  6.940000  8.645000 12.800000  8.965000 ;
      RECT  6.940000  8.965000  7.080000 11.380000 ;
      RECT  7.220000  0.330000  7.360000  2.745000 ;
      RECT  7.220000  3.345000  7.360000  5.760000 ;
      RECT  7.220000  6.090000  7.360000  8.505000 ;
      RECT  7.220000  9.105000  7.360000 11.520000 ;
      RECT  7.500000  0.470000  7.640000  2.885000 ;
      RECT  7.500000  3.205000  7.640000  5.620000 ;
      RECT  7.500000  6.230000  7.640000  8.645000 ;
      RECT  7.500000  8.965000  7.640000 11.380000 ;
      RECT  7.780000  0.330000  7.920000  2.745000 ;
      RECT  7.780000  3.345000  7.920000  5.760000 ;
      RECT  7.780000  6.090000  7.920000  8.505000 ;
      RECT  7.780000  9.105000  7.920000 11.520000 ;
      RECT  8.060000  0.470000  8.200000  2.885000 ;
      RECT  8.060000  3.205000  8.200000  5.620000 ;
      RECT  8.060000  6.230000  8.200000  8.645000 ;
      RECT  8.060000  8.965000  8.200000 11.380000 ;
      RECT  8.340000  0.330000  8.480000  2.745000 ;
      RECT  8.340000  3.345000  8.480000  5.760000 ;
      RECT  8.340000  6.090000  8.480000  8.505000 ;
      RECT  8.340000  9.105000  8.480000 11.520000 ;
      RECT  8.620000  0.470000  8.760000  2.885000 ;
      RECT  8.620000  3.205000  8.760000  5.620000 ;
      RECT  8.620000  6.230000  8.760000  8.645000 ;
      RECT  8.620000  8.965000  8.760000 11.380000 ;
      RECT  8.900000  0.330000  9.040000  2.745000 ;
      RECT  8.900000  3.345000  9.040000  5.760000 ;
      RECT  8.900000  6.090000  9.040000  8.505000 ;
      RECT  8.900000  9.105000  9.040000 11.520000 ;
      RECT  9.180000  0.470000  9.320000  2.885000 ;
      RECT  9.180000  3.205000  9.320000  5.620000 ;
      RECT  9.180000  6.230000  9.320000  8.645000 ;
      RECT  9.180000  8.965000  9.320000 11.380000 ;
      RECT  9.460000  0.330000  9.600000  2.745000 ;
      RECT  9.460000  3.345000  9.600000  5.760000 ;
      RECT  9.460000  6.090000  9.600000  8.505000 ;
      RECT  9.460000  9.105000  9.600000 11.520000 ;
      RECT  9.740000  0.470000 10.000000  2.885000 ;
      RECT  9.740000  3.205000 10.000000  5.620000 ;
      RECT  9.740000  6.230000 10.000000  8.645000 ;
      RECT  9.740000  8.965000 10.000000 11.380000 ;
      RECT 10.140000  0.330000 10.280000  2.745000 ;
      RECT 10.140000  3.345000 10.280000  5.760000 ;
      RECT 10.140000  6.090000 10.280000  8.505000 ;
      RECT 10.140000  9.105000 10.280000 11.520000 ;
      RECT 10.420000  0.470000 10.560000  2.885000 ;
      RECT 10.420000  3.205000 10.560000  5.620000 ;
      RECT 10.420000  6.230000 10.560000  8.645000 ;
      RECT 10.420000  8.965000 10.560000 11.380000 ;
      RECT 10.700000  0.330000 10.840000  2.745000 ;
      RECT 10.700000  3.345000 10.840000  5.760000 ;
      RECT 10.700000  6.090000 10.840000  8.505000 ;
      RECT 10.700000  9.105000 10.840000 11.520000 ;
      RECT 10.980000  0.470000 11.120000  2.885000 ;
      RECT 10.980000  3.205000 11.120000  5.620000 ;
      RECT 10.980000  6.230000 11.120000  8.645000 ;
      RECT 10.980000  8.965000 11.120000 11.380000 ;
      RECT 11.260000  0.330000 11.400000  2.745000 ;
      RECT 11.260000  3.345000 11.400000  5.760000 ;
      RECT 11.260000  6.090000 11.400000  8.505000 ;
      RECT 11.260000  9.105000 11.400000 11.520000 ;
      RECT 11.540000  0.470000 11.680000  2.885000 ;
      RECT 11.540000  3.205000 11.680000  5.620000 ;
      RECT 11.540000  6.230000 11.680000  8.645000 ;
      RECT 11.540000  8.965000 11.680000 11.380000 ;
      RECT 11.820000  0.330000 11.960000  2.745000 ;
      RECT 11.820000  3.345000 11.960000  5.760000 ;
      RECT 11.820000  6.090000 11.960000  8.505000 ;
      RECT 11.820000  9.105000 11.960000 11.520000 ;
      RECT 12.100000  0.470000 12.240000  2.885000 ;
      RECT 12.100000  3.205000 12.240000  5.620000 ;
      RECT 12.100000  6.230000 12.240000  8.645000 ;
      RECT 12.100000  8.965000 12.240000 11.380000 ;
      RECT 12.380000  0.330000 12.520000  2.745000 ;
      RECT 12.380000  3.345000 12.520000  5.760000 ;
      RECT 12.380000  6.090000 12.520000  8.505000 ;
      RECT 12.380000  9.105000 12.520000 11.520000 ;
      RECT 12.660000  0.470000 12.800000  2.885000 ;
      RECT 12.660000  3.205000 12.800000  5.620000 ;
      RECT 12.660000  6.230000 12.800000  8.645000 ;
      RECT 12.660000  8.965000 12.800000 11.380000 ;
      RECT 12.940000  0.330000 13.270000  5.760000 ;
      RECT 12.940000  6.090000 13.270000 11.520000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  3.095000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.750000 ;
      RECT  0.000000  0.750000  3.095000  0.890000 ;
      RECT  0.000000  0.890000  0.330000  1.310000 ;
      RECT  0.000000  1.310000  3.095000  1.450000 ;
      RECT  0.000000  1.450000  0.330000  1.870000 ;
      RECT  0.000000  1.870000  3.095000  2.010000 ;
      RECT  0.000000  2.010000  0.330000  2.430000 ;
      RECT  0.000000  2.430000  3.095000  2.765000 ;
      RECT  0.000000  2.905000 13.270000  3.185000 ;
      RECT  0.000000  3.325000  3.095000  3.660000 ;
      RECT  0.000000  3.660000  0.330000  4.080000 ;
      RECT  0.000000  4.080000  3.095000  4.220000 ;
      RECT  0.000000  4.220000  0.330000  4.640000 ;
      RECT  0.000000  4.640000  3.095000  4.780000 ;
      RECT  0.000000  4.780000  0.330000  5.200000 ;
      RECT  0.000000  5.200000  3.095000  5.340000 ;
      RECT  0.000000  5.340000  0.330000  5.760000 ;
      RECT  0.000000  5.760000  3.095000  6.090000 ;
      RECT  0.000000  6.090000  0.330000  6.510000 ;
      RECT  0.000000  6.510000  3.095000  6.650000 ;
      RECT  0.000000  6.650000  0.330000  7.070000 ;
      RECT  0.000000  7.070000  3.095000  7.210000 ;
      RECT  0.000000  7.210000  0.330000  7.630000 ;
      RECT  0.000000  7.630000  3.095000  7.770000 ;
      RECT  0.000000  7.770000  0.330000  8.190000 ;
      RECT  0.000000  8.190000  3.095000  8.525000 ;
      RECT  0.000000  8.665000 13.270000  8.945000 ;
      RECT  0.000000  9.085000  3.095000  9.420000 ;
      RECT  0.000000  9.420000  0.330000  9.840000 ;
      RECT  0.000000  9.840000  3.095000  9.980000 ;
      RECT  0.000000  9.980000  0.330000 10.400000 ;
      RECT  0.000000 10.400000  3.095000 10.540000 ;
      RECT  0.000000 10.540000  0.330000 10.960000 ;
      RECT  0.000000 10.960000  3.095000 11.100000 ;
      RECT  0.000000 11.100000  0.330000 11.520000 ;
      RECT  0.000000 11.520000  3.095000 11.850000 ;
      RECT  0.470000  0.470000  6.330000  0.610000 ;
      RECT  0.470000  1.030000  6.330000  1.170000 ;
      RECT  0.470000  1.590000  6.330000  1.730000 ;
      RECT  0.470000  2.150000  6.330000  2.290000 ;
      RECT  0.470000  3.800000  6.330000  3.940000 ;
      RECT  0.470000  4.360000  6.330000  4.500000 ;
      RECT  0.470000  4.920000  6.330000  5.060000 ;
      RECT  0.470000  5.480000  6.330000  5.620000 ;
      RECT  0.470000  6.230000  6.330000  6.370000 ;
      RECT  0.470000  6.790000  6.330000  6.930000 ;
      RECT  0.470000  7.350000  6.330000  7.490000 ;
      RECT  0.470000  7.910000  6.330000  8.050000 ;
      RECT  0.470000  9.560000  6.330000  9.700000 ;
      RECT  0.470000 10.120000  6.330000 10.260000 ;
      RECT  0.470000 10.680000  6.330000 10.820000 ;
      RECT  0.470000 11.240000  6.330000 11.380000 ;
      RECT  3.235000  0.000000  3.565000  0.470000 ;
      RECT  3.235000  0.610000  3.565000  1.030000 ;
      RECT  3.235000  1.170000  3.565000  1.590000 ;
      RECT  3.235000  1.730000  3.565000  2.150000 ;
      RECT  3.235000  2.290000  3.565000  2.905000 ;
      RECT  3.235000  3.185000  3.565000  3.800000 ;
      RECT  3.235000  3.940000  3.565000  4.360000 ;
      RECT  3.235000  4.500000  3.565000  4.920000 ;
      RECT  3.235000  5.060000  3.565000  5.480000 ;
      RECT  3.235000  5.620000  3.565000  6.230000 ;
      RECT  3.235000  6.370000  3.565000  6.790000 ;
      RECT  3.235000  6.930000  3.565000  7.350000 ;
      RECT  3.235000  7.490000  3.565000  7.910000 ;
      RECT  3.235000  8.050000  3.565000  8.665000 ;
      RECT  3.235000  8.945000  3.565000  9.560000 ;
      RECT  3.235000  9.700000  3.565000 10.120000 ;
      RECT  3.235000 10.260000  3.565000 10.680000 ;
      RECT  3.235000 10.820000  3.565000 11.240000 ;
      RECT  3.235000 11.380000  3.565000 11.850000 ;
      RECT  3.705000  0.000000  9.565000  0.330000 ;
      RECT  3.705000  0.750000  9.565000  0.890000 ;
      RECT  3.705000  1.310000  9.565000  1.450000 ;
      RECT  3.705000  1.870000  9.565000  2.010000 ;
      RECT  3.705000  2.430000  9.565000  2.765000 ;
      RECT  3.705000  3.325000  9.565000  3.660000 ;
      RECT  3.705000  4.080000  9.565000  4.220000 ;
      RECT  3.705000  4.640000  9.565000  4.780000 ;
      RECT  3.705000  5.200000  9.565000  5.340000 ;
      RECT  3.705000  5.760000  9.565000  6.090000 ;
      RECT  3.705000  6.510000  9.565000  6.650000 ;
      RECT  3.705000  7.070000  9.565000  7.210000 ;
      RECT  3.705000  7.630000  9.565000  7.770000 ;
      RECT  3.705000  8.190000  9.565000  8.525000 ;
      RECT  3.705000  9.085000  9.565000  9.420000 ;
      RECT  3.705000  9.840000  9.565000  9.980000 ;
      RECT  3.705000 10.400000  9.565000 10.540000 ;
      RECT  3.705000 10.960000  9.565000 11.100000 ;
      RECT  3.705000 11.520000  9.565000 11.850000 ;
      RECT  6.470000  0.330000  6.800000  0.750000 ;
      RECT  6.470000  0.890000  6.800000  1.310000 ;
      RECT  6.470000  1.450000  6.800000  1.870000 ;
      RECT  6.470000  2.010000  6.800000  2.430000 ;
      RECT  6.470000  3.660000  6.800000  4.080000 ;
      RECT  6.470000  4.220000  6.800000  4.640000 ;
      RECT  6.470000  4.780000  6.800000  5.200000 ;
      RECT  6.470000  5.340000  6.800000  5.760000 ;
      RECT  6.470000  6.090000  6.800000  6.510000 ;
      RECT  6.470000  6.650000  6.800000  7.070000 ;
      RECT  6.470000  7.210000  6.800000  7.630000 ;
      RECT  6.470000  7.770000  6.800000  8.190000 ;
      RECT  6.470000  9.420000  6.800000  9.840000 ;
      RECT  6.470000  9.980000  6.800000 10.400000 ;
      RECT  6.470000 10.540000  6.800000 10.960000 ;
      RECT  6.470000 11.100000  6.800000 11.520000 ;
      RECT  6.940000  0.470000 12.800000  0.610000 ;
      RECT  6.940000  1.030000 12.800000  1.170000 ;
      RECT  6.940000  1.590000 12.800000  1.730000 ;
      RECT  6.940000  2.150000 12.800000  2.290000 ;
      RECT  6.940000  3.800000 12.800000  3.940000 ;
      RECT  6.940000  4.360000 12.800000  4.500000 ;
      RECT  6.940000  4.920000 12.800000  5.060000 ;
      RECT  6.940000  5.480000 12.800000  5.620000 ;
      RECT  6.940000  6.230000 12.800000  6.370000 ;
      RECT  6.940000  6.790000 12.800000  6.930000 ;
      RECT  6.940000  7.350000 12.800000  7.490000 ;
      RECT  6.940000  7.910000 12.800000  8.050000 ;
      RECT  6.940000  9.560000 12.800000  9.700000 ;
      RECT  6.940000 10.120000 12.800000 10.260000 ;
      RECT  6.940000 10.680000 12.800000 10.820000 ;
      RECT  6.940000 11.240000 12.800000 11.380000 ;
      RECT  9.705000  0.000000 10.035000  0.470000 ;
      RECT  9.705000  0.610000 10.035000  1.030000 ;
      RECT  9.705000  1.170000 10.035000  1.590000 ;
      RECT  9.705000  1.730000 10.035000  2.150000 ;
      RECT  9.705000  2.290000 10.035000  2.905000 ;
      RECT  9.705000  3.185000 10.035000  3.800000 ;
      RECT  9.705000  3.940000 10.035000  4.360000 ;
      RECT  9.705000  4.500000 10.035000  4.920000 ;
      RECT  9.705000  5.060000 10.035000  5.480000 ;
      RECT  9.705000  5.620000 10.035000  6.230000 ;
      RECT  9.705000  6.370000 10.035000  6.790000 ;
      RECT  9.705000  6.930000 10.035000  7.350000 ;
      RECT  9.705000  7.490000 10.035000  7.910000 ;
      RECT  9.705000  8.050000 10.035000  8.665000 ;
      RECT  9.705000  8.945000 10.035000  9.560000 ;
      RECT  9.705000  9.700000 10.035000 10.120000 ;
      RECT  9.705000 10.260000 10.035000 10.680000 ;
      RECT  9.705000 10.820000 10.035000 11.240000 ;
      RECT  9.705000 11.380000 10.035000 11.850000 ;
      RECT 10.175000  0.000000 13.270000  0.330000 ;
      RECT 10.175000  0.750000 13.270000  0.890000 ;
      RECT 10.175000  1.310000 13.270000  1.450000 ;
      RECT 10.175000  1.870000 13.270000  2.010000 ;
      RECT 10.175000  2.430000 13.270000  2.765000 ;
      RECT 10.175000  3.325000 13.270000  3.660000 ;
      RECT 10.175000  4.080000 13.270000  4.220000 ;
      RECT 10.175000  4.640000 13.270000  4.780000 ;
      RECT 10.175000  5.200000 13.270000  5.340000 ;
      RECT 10.175000  5.760000 13.270000  6.090000 ;
      RECT 10.175000  6.510000 13.270000  6.650000 ;
      RECT 10.175000  7.070000 13.270000  7.210000 ;
      RECT 10.175000  7.630000 13.270000  7.770000 ;
      RECT 10.175000  8.190000 13.270000  8.525000 ;
      RECT 10.175000  9.085000 13.270000  9.420000 ;
      RECT 10.175000  9.840000 13.270000  9.980000 ;
      RECT 10.175000 10.400000 13.270000 10.540000 ;
      RECT 10.175000 10.960000 13.270000 11.100000 ;
      RECT 10.175000 11.520000 13.270000 11.850000 ;
      RECT 12.940000  0.330000 13.270000  0.750000 ;
      RECT 12.940000  0.890000 13.270000  1.310000 ;
      RECT 12.940000  1.450000 13.270000  1.870000 ;
      RECT 12.940000  2.010000 13.270000  2.430000 ;
      RECT 12.940000  3.660000 13.270000  4.080000 ;
      RECT 12.940000  4.220000 13.270000  4.640000 ;
      RECT 12.940000  4.780000 13.270000  5.200000 ;
      RECT 12.940000  5.340000 13.270000  5.760000 ;
      RECT 12.940000  6.090000 13.270000  6.510000 ;
      RECT 12.940000  6.650000 13.270000  7.070000 ;
      RECT 12.940000  7.210000 13.270000  7.630000 ;
      RECT 12.940000  7.770000 13.270000  8.190000 ;
      RECT 12.940000  9.420000 13.270000  9.840000 ;
      RECT 12.940000  9.980000 13.270000 10.400000 ;
      RECT 12.940000 10.540000 13.270000 10.960000 ;
      RECT 12.940000 11.100000 13.270000 11.520000 ;
    LAYER pwell ;
      RECT 2.735000  4.370000 2.840000  4.615000 ;
      RECT 2.735000 10.130000 2.840000 10.375000 ;
      RECT 9.205000  4.370000 9.310000  4.615000 ;
      RECT 9.205000 10.130000 9.310000 10.375000 ;
    LAYER via ;
      RECT  0.035000  0.355000  0.295000  0.615000 ;
      RECT  0.035000  0.675000  0.295000  0.935000 ;
      RECT  0.035000  0.995000  0.295000  1.255000 ;
      RECT  0.035000  1.315000  0.295000  1.575000 ;
      RECT  0.035000  1.635000  0.295000  1.895000 ;
      RECT  0.035000  1.955000  0.295000  2.215000 ;
      RECT  0.035000  2.275000  0.295000  2.535000 ;
      RECT  0.035000  3.555000  0.295000  3.815000 ;
      RECT  0.035000  3.875000  0.295000  4.135000 ;
      RECT  0.035000  4.195000  0.295000  4.455000 ;
      RECT  0.035000  4.515000  0.295000  4.775000 ;
      RECT  0.035000  4.835000  0.295000  5.095000 ;
      RECT  0.035000  5.155000  0.295000  5.415000 ;
      RECT  0.035000  5.475000  0.295000  5.735000 ;
      RECT  0.035000  6.115000  0.295000  6.375000 ;
      RECT  0.035000  6.435000  0.295000  6.695000 ;
      RECT  0.035000  6.755000  0.295000  7.015000 ;
      RECT  0.035000  7.075000  0.295000  7.335000 ;
      RECT  0.035000  7.395000  0.295000  7.655000 ;
      RECT  0.035000  7.715000  0.295000  7.975000 ;
      RECT  0.035000  8.035000  0.295000  8.295000 ;
      RECT  0.035000  9.315000  0.295000  9.575000 ;
      RECT  0.035000  9.635000  0.295000  9.895000 ;
      RECT  0.035000  9.955000  0.295000 10.215000 ;
      RECT  0.035000 10.275000  0.295000 10.535000 ;
      RECT  0.035000 10.595000  0.295000 10.855000 ;
      RECT  0.035000 10.915000  0.295000 11.175000 ;
      RECT  0.035000 11.235000  0.295000 11.495000 ;
      RECT  0.365000  0.035000  0.625000  0.295000 ;
      RECT  0.365000  5.795000  0.625000  6.055000 ;
      RECT  0.365000 11.555000  0.625000 11.815000 ;
      RECT  0.525000  2.915000  0.785000  3.175000 ;
      RECT  0.525000  8.675000  0.785000  8.935000 ;
      RECT  0.685000  0.035000  0.945000  0.295000 ;
      RECT  0.685000  5.795000  0.945000  6.055000 ;
      RECT  0.685000 11.555000  0.945000 11.815000 ;
      RECT  0.845000  2.915000  1.105000  3.175000 ;
      RECT  0.845000  8.675000  1.105000  8.935000 ;
      RECT  1.005000  0.035000  1.265000  0.295000 ;
      RECT  1.005000  5.795000  1.265000  6.055000 ;
      RECT  1.005000 11.555000  1.265000 11.815000 ;
      RECT  1.165000  2.915000  1.425000  3.175000 ;
      RECT  1.165000  8.675000  1.425000  8.935000 ;
      RECT  1.325000  0.035000  1.585000  0.295000 ;
      RECT  1.325000  5.795000  1.585000  6.055000 ;
      RECT  1.325000 11.555000  1.585000 11.815000 ;
      RECT  1.485000  2.915000  1.745000  3.175000 ;
      RECT  1.485000  8.675000  1.745000  8.935000 ;
      RECT  1.645000  0.035000  1.905000  0.295000 ;
      RECT  1.645000  5.795000  1.905000  6.055000 ;
      RECT  1.645000 11.555000  1.905000 11.815000 ;
      RECT  1.805000  2.915000  2.065000  3.175000 ;
      RECT  1.805000  8.675000  2.065000  8.935000 ;
      RECT  1.965000  0.035000  2.225000  0.295000 ;
      RECT  1.965000  5.795000  2.225000  6.055000 ;
      RECT  1.965000 11.555000  2.225000 11.815000 ;
      RECT  2.125000  2.915000  2.385000  3.175000 ;
      RECT  2.125000  8.675000  2.385000  8.935000 ;
      RECT  2.285000  0.035000  2.545000  0.295000 ;
      RECT  2.285000  5.795000  2.545000  6.055000 ;
      RECT  2.285000 11.555000  2.545000 11.815000 ;
      RECT  2.445000  2.915000  2.705000  3.175000 ;
      RECT  2.445000  8.675000  2.705000  8.935000 ;
      RECT  2.605000  0.035000  2.865000  0.295000 ;
      RECT  2.605000  5.795000  2.865000  6.055000 ;
      RECT  2.605000 11.555000  2.865000 11.815000 ;
      RECT  2.765000  2.915000  3.025000  3.175000 ;
      RECT  2.765000  8.675000  3.025000  8.935000 ;
      RECT  3.085000  2.915000  3.345000  3.175000 ;
      RECT  3.085000  8.675000  3.345000  8.935000 ;
      RECT  3.270000  0.515000  3.530000  0.775000 ;
      RECT  3.270000  0.835000  3.530000  1.095000 ;
      RECT  3.270000  1.155000  3.530000  1.415000 ;
      RECT  3.270000  1.475000  3.530000  1.735000 ;
      RECT  3.270000  1.795000  3.530000  2.055000 ;
      RECT  3.270000  2.115000  3.530000  2.375000 ;
      RECT  3.270000  2.435000  3.530000  2.695000 ;
      RECT  3.270000  3.395000  3.530000  3.655000 ;
      RECT  3.270000  3.715000  3.530000  3.975000 ;
      RECT  3.270000  4.035000  3.530000  4.295000 ;
      RECT  3.270000  4.355000  3.530000  4.615000 ;
      RECT  3.270000  4.675000  3.530000  4.935000 ;
      RECT  3.270000  4.995000  3.530000  5.255000 ;
      RECT  3.270000  5.315000  3.530000  5.575000 ;
      RECT  3.270000  6.275000  3.530000  6.535000 ;
      RECT  3.270000  6.595000  3.530000  6.855000 ;
      RECT  3.270000  6.915000  3.530000  7.175000 ;
      RECT  3.270000  7.235000  3.530000  7.495000 ;
      RECT  3.270000  7.555000  3.530000  7.815000 ;
      RECT  3.270000  7.875000  3.530000  8.135000 ;
      RECT  3.270000  8.195000  3.530000  8.455000 ;
      RECT  3.270000  9.155000  3.530000  9.415000 ;
      RECT  3.270000  9.475000  3.530000  9.735000 ;
      RECT  3.270000  9.795000  3.530000 10.055000 ;
      RECT  3.270000 10.115000  3.530000 10.375000 ;
      RECT  3.270000 10.435000  3.530000 10.695000 ;
      RECT  3.270000 10.755000  3.530000 11.015000 ;
      RECT  3.270000 11.075000  3.530000 11.335000 ;
      RECT  3.455000  2.915000  3.715000  3.175000 ;
      RECT  3.455000  8.675000  3.715000  8.935000 ;
      RECT  3.775000  2.915000  4.035000  3.175000 ;
      RECT  3.775000  8.675000  4.035000  8.935000 ;
      RECT  3.935000  0.035000  4.195000  0.295000 ;
      RECT  3.935000  5.795000  4.195000  6.055000 ;
      RECT  3.935000 11.555000  4.195000 11.815000 ;
      RECT  4.095000  2.915000  4.355000  3.175000 ;
      RECT  4.095000  8.675000  4.355000  8.935000 ;
      RECT  4.255000  0.035000  4.515000  0.295000 ;
      RECT  4.255000  5.795000  4.515000  6.055000 ;
      RECT  4.255000 11.555000  4.515000 11.815000 ;
      RECT  4.415000  2.915000  4.675000  3.175000 ;
      RECT  4.415000  8.675000  4.675000  8.935000 ;
      RECT  4.575000  0.035000  4.835000  0.295000 ;
      RECT  4.575000  5.795000  4.835000  6.055000 ;
      RECT  4.575000 11.555000  4.835000 11.815000 ;
      RECT  4.735000  2.915000  4.995000  3.175000 ;
      RECT  4.735000  8.675000  4.995000  8.935000 ;
      RECT  4.895000  0.035000  5.155000  0.295000 ;
      RECT  4.895000  5.795000  5.155000  6.055000 ;
      RECT  4.895000 11.555000  5.155000 11.815000 ;
      RECT  5.055000  2.915000  5.315000  3.175000 ;
      RECT  5.055000  8.675000  5.315000  8.935000 ;
      RECT  5.215000  0.035000  5.475000  0.295000 ;
      RECT  5.215000  5.795000  5.475000  6.055000 ;
      RECT  5.215000 11.555000  5.475000 11.815000 ;
      RECT  5.375000  2.915000  5.635000  3.175000 ;
      RECT  5.375000  8.675000  5.635000  8.935000 ;
      RECT  5.535000  0.035000  5.795000  0.295000 ;
      RECT  5.535000  5.795000  5.795000  6.055000 ;
      RECT  5.535000 11.555000  5.795000 11.815000 ;
      RECT  5.695000  2.915000  5.955000  3.175000 ;
      RECT  5.695000  8.675000  5.955000  8.935000 ;
      RECT  5.855000  0.035000  6.115000  0.295000 ;
      RECT  5.855000  5.795000  6.115000  6.055000 ;
      RECT  5.855000 11.555000  6.115000 11.815000 ;
      RECT  6.015000  2.915000  6.275000  3.175000 ;
      RECT  6.015000  8.675000  6.275000  8.935000 ;
      RECT  6.175000  0.035000  6.435000  0.295000 ;
      RECT  6.175000  5.795000  6.435000  6.055000 ;
      RECT  6.175000 11.555000  6.435000 11.815000 ;
      RECT  6.505000  0.355000  6.765000  0.615000 ;
      RECT  6.505000  0.675000  6.765000  0.935000 ;
      RECT  6.505000  0.995000  6.765000  1.255000 ;
      RECT  6.505000  1.315000  6.765000  1.575000 ;
      RECT  6.505000  1.635000  6.765000  1.895000 ;
      RECT  6.505000  1.955000  6.765000  2.215000 ;
      RECT  6.505000  2.275000  6.765000  2.535000 ;
      RECT  6.505000  3.555000  6.765000  3.815000 ;
      RECT  6.505000  3.875000  6.765000  4.135000 ;
      RECT  6.505000  4.195000  6.765000  4.455000 ;
      RECT  6.505000  4.515000  6.765000  4.775000 ;
      RECT  6.505000  4.835000  6.765000  5.095000 ;
      RECT  6.505000  5.155000  6.765000  5.415000 ;
      RECT  6.505000  5.475000  6.765000  5.735000 ;
      RECT  6.505000  6.115000  6.765000  6.375000 ;
      RECT  6.505000  6.435000  6.765000  6.695000 ;
      RECT  6.505000  6.755000  6.765000  7.015000 ;
      RECT  6.505000  7.075000  6.765000  7.335000 ;
      RECT  6.505000  7.395000  6.765000  7.655000 ;
      RECT  6.505000  7.715000  6.765000  7.975000 ;
      RECT  6.505000  8.035000  6.765000  8.295000 ;
      RECT  6.505000  9.315000  6.765000  9.575000 ;
      RECT  6.505000  9.635000  6.765000  9.895000 ;
      RECT  6.505000  9.955000  6.765000 10.215000 ;
      RECT  6.505000 10.275000  6.765000 10.535000 ;
      RECT  6.505000 10.595000  6.765000 10.855000 ;
      RECT  6.505000 10.915000  6.765000 11.175000 ;
      RECT  6.505000 11.235000  6.765000 11.495000 ;
      RECT  6.835000  0.035000  7.095000  0.295000 ;
      RECT  6.835000  5.795000  7.095000  6.055000 ;
      RECT  6.835000 11.555000  7.095000 11.815000 ;
      RECT  6.995000  2.915000  7.255000  3.175000 ;
      RECT  6.995000  8.675000  7.255000  8.935000 ;
      RECT  7.155000  0.035000  7.415000  0.295000 ;
      RECT  7.155000  5.795000  7.415000  6.055000 ;
      RECT  7.155000 11.555000  7.415000 11.815000 ;
      RECT  7.315000  2.915000  7.575000  3.175000 ;
      RECT  7.315000  8.675000  7.575000  8.935000 ;
      RECT  7.475000  0.035000  7.735000  0.295000 ;
      RECT  7.475000  5.795000  7.735000  6.055000 ;
      RECT  7.475000 11.555000  7.735000 11.815000 ;
      RECT  7.635000  2.915000  7.895000  3.175000 ;
      RECT  7.635000  8.675000  7.895000  8.935000 ;
      RECT  7.795000  0.035000  8.055000  0.295000 ;
      RECT  7.795000  5.795000  8.055000  6.055000 ;
      RECT  7.795000 11.555000  8.055000 11.815000 ;
      RECT  7.955000  2.915000  8.215000  3.175000 ;
      RECT  7.955000  8.675000  8.215000  8.935000 ;
      RECT  8.115000  0.035000  8.375000  0.295000 ;
      RECT  8.115000  5.795000  8.375000  6.055000 ;
      RECT  8.115000 11.555000  8.375000 11.815000 ;
      RECT  8.275000  2.915000  8.535000  3.175000 ;
      RECT  8.275000  8.675000  8.535000  8.935000 ;
      RECT  8.435000  0.035000  8.695000  0.295000 ;
      RECT  8.435000  5.795000  8.695000  6.055000 ;
      RECT  8.435000 11.555000  8.695000 11.815000 ;
      RECT  8.595000  2.915000  8.855000  3.175000 ;
      RECT  8.595000  8.675000  8.855000  8.935000 ;
      RECT  8.755000  0.035000  9.015000  0.295000 ;
      RECT  8.755000  5.795000  9.015000  6.055000 ;
      RECT  8.755000 11.555000  9.015000 11.815000 ;
      RECT  8.915000  2.915000  9.175000  3.175000 ;
      RECT  8.915000  8.675000  9.175000  8.935000 ;
      RECT  9.075000  0.035000  9.335000  0.295000 ;
      RECT  9.075000  5.795000  9.335000  6.055000 ;
      RECT  9.075000 11.555000  9.335000 11.815000 ;
      RECT  9.235000  2.915000  9.495000  3.175000 ;
      RECT  9.235000  8.675000  9.495000  8.935000 ;
      RECT  9.555000  2.915000  9.815000  3.175000 ;
      RECT  9.555000  8.675000  9.815000  8.935000 ;
      RECT  9.740000  0.515000 10.000000  0.775000 ;
      RECT  9.740000  0.835000 10.000000  1.095000 ;
      RECT  9.740000  1.155000 10.000000  1.415000 ;
      RECT  9.740000  1.475000 10.000000  1.735000 ;
      RECT  9.740000  1.795000 10.000000  2.055000 ;
      RECT  9.740000  2.115000 10.000000  2.375000 ;
      RECT  9.740000  2.435000 10.000000  2.695000 ;
      RECT  9.740000  3.395000 10.000000  3.655000 ;
      RECT  9.740000  3.715000 10.000000  3.975000 ;
      RECT  9.740000  4.035000 10.000000  4.295000 ;
      RECT  9.740000  4.355000 10.000000  4.615000 ;
      RECT  9.740000  4.675000 10.000000  4.935000 ;
      RECT  9.740000  4.995000 10.000000  5.255000 ;
      RECT  9.740000  5.315000 10.000000  5.575000 ;
      RECT  9.740000  6.275000 10.000000  6.535000 ;
      RECT  9.740000  6.595000 10.000000  6.855000 ;
      RECT  9.740000  6.915000 10.000000  7.175000 ;
      RECT  9.740000  7.235000 10.000000  7.495000 ;
      RECT  9.740000  7.555000 10.000000  7.815000 ;
      RECT  9.740000  7.875000 10.000000  8.135000 ;
      RECT  9.740000  8.195000 10.000000  8.455000 ;
      RECT  9.740000  9.155000 10.000000  9.415000 ;
      RECT  9.740000  9.475000 10.000000  9.735000 ;
      RECT  9.740000  9.795000 10.000000 10.055000 ;
      RECT  9.740000 10.115000 10.000000 10.375000 ;
      RECT  9.740000 10.435000 10.000000 10.695000 ;
      RECT  9.740000 10.755000 10.000000 11.015000 ;
      RECT  9.740000 11.075000 10.000000 11.335000 ;
      RECT  9.925000  2.915000 10.185000  3.175000 ;
      RECT  9.925000  8.675000 10.185000  8.935000 ;
      RECT 10.245000  2.915000 10.505000  3.175000 ;
      RECT 10.245000  8.675000 10.505000  8.935000 ;
      RECT 10.405000  0.035000 10.665000  0.295000 ;
      RECT 10.405000  5.795000 10.665000  6.055000 ;
      RECT 10.405000 11.555000 10.665000 11.815000 ;
      RECT 10.565000  2.915000 10.825000  3.175000 ;
      RECT 10.565000  8.675000 10.825000  8.935000 ;
      RECT 10.725000  0.035000 10.985000  0.295000 ;
      RECT 10.725000  5.795000 10.985000  6.055000 ;
      RECT 10.725000 11.555000 10.985000 11.815000 ;
      RECT 10.885000  2.915000 11.145000  3.175000 ;
      RECT 10.885000  8.675000 11.145000  8.935000 ;
      RECT 11.045000  0.035000 11.305000  0.295000 ;
      RECT 11.045000  5.795000 11.305000  6.055000 ;
      RECT 11.045000 11.555000 11.305000 11.815000 ;
      RECT 11.205000  2.915000 11.465000  3.175000 ;
      RECT 11.205000  8.675000 11.465000  8.935000 ;
      RECT 11.365000  0.035000 11.625000  0.295000 ;
      RECT 11.365000  5.795000 11.625000  6.055000 ;
      RECT 11.365000 11.555000 11.625000 11.815000 ;
      RECT 11.525000  2.915000 11.785000  3.175000 ;
      RECT 11.525000  8.675000 11.785000  8.935000 ;
      RECT 11.685000  0.035000 11.945000  0.295000 ;
      RECT 11.685000  5.795000 11.945000  6.055000 ;
      RECT 11.685000 11.555000 11.945000 11.815000 ;
      RECT 11.845000  2.915000 12.105000  3.175000 ;
      RECT 11.845000  8.675000 12.105000  8.935000 ;
      RECT 12.005000  0.035000 12.265000  0.295000 ;
      RECT 12.005000  5.795000 12.265000  6.055000 ;
      RECT 12.005000 11.555000 12.265000 11.815000 ;
      RECT 12.165000  2.915000 12.425000  3.175000 ;
      RECT 12.165000  8.675000 12.425000  8.935000 ;
      RECT 12.325000  0.035000 12.585000  0.295000 ;
      RECT 12.325000  5.795000 12.585000  6.055000 ;
      RECT 12.325000 11.555000 12.585000 11.815000 ;
      RECT 12.485000  2.915000 12.745000  3.175000 ;
      RECT 12.485000  8.675000 12.745000  8.935000 ;
      RECT 12.645000  0.035000 12.905000  0.295000 ;
      RECT 12.645000  5.795000 12.905000  6.055000 ;
      RECT 12.645000 11.555000 12.905000 11.815000 ;
      RECT 12.975000  0.355000 13.235000  0.615000 ;
      RECT 12.975000  0.675000 13.235000  0.935000 ;
      RECT 12.975000  0.995000 13.235000  1.255000 ;
      RECT 12.975000  1.315000 13.235000  1.575000 ;
      RECT 12.975000  1.635000 13.235000  1.895000 ;
      RECT 12.975000  1.955000 13.235000  2.215000 ;
      RECT 12.975000  2.275000 13.235000  2.535000 ;
      RECT 12.975000  3.555000 13.235000  3.815000 ;
      RECT 12.975000  3.875000 13.235000  4.135000 ;
      RECT 12.975000  4.195000 13.235000  4.455000 ;
      RECT 12.975000  4.515000 13.235000  4.775000 ;
      RECT 12.975000  4.835000 13.235000  5.095000 ;
      RECT 12.975000  5.155000 13.235000  5.415000 ;
      RECT 12.975000  5.475000 13.235000  5.735000 ;
      RECT 12.975000  6.115000 13.235000  6.375000 ;
      RECT 12.975000  6.435000 13.235000  6.695000 ;
      RECT 12.975000  6.755000 13.235000  7.015000 ;
      RECT 12.975000  7.075000 13.235000  7.335000 ;
      RECT 12.975000  7.395000 13.235000  7.655000 ;
      RECT 12.975000  7.715000 13.235000  7.975000 ;
      RECT 12.975000  8.035000 13.235000  8.295000 ;
      RECT 12.975000  9.315000 13.235000  9.575000 ;
      RECT 12.975000  9.635000 13.235000  9.895000 ;
      RECT 12.975000  9.955000 13.235000 10.215000 ;
      RECT 12.975000 10.275000 13.235000 10.535000 ;
      RECT 12.975000 10.595000 13.235000 10.855000 ;
      RECT 12.975000 10.915000 13.235000 11.175000 ;
      RECT 12.975000 11.235000 13.235000 11.495000 ;
    LAYER via2 ;
      RECT  0.025000  0.400000  0.305000  0.680000 ;
      RECT  0.025000  0.800000  0.305000  1.080000 ;
      RECT  0.025000  1.200000  0.305000  1.480000 ;
      RECT  0.025000  1.600000  0.305000  1.880000 ;
      RECT  0.025000  2.000000  0.305000  2.280000 ;
      RECT  0.025000  2.400000  0.305000  2.680000 ;
      RECT  0.025000  3.410000  0.305000  3.690000 ;
      RECT  0.025000  3.810000  0.305000  4.090000 ;
      RECT  0.025000  4.210000  0.305000  4.490000 ;
      RECT  0.025000  4.610000  0.305000  4.890000 ;
      RECT  0.025000  5.010000  0.305000  5.290000 ;
      RECT  0.025000  5.410000  0.305000  5.690000 ;
      RECT  0.025000  6.160000  0.305000  6.440000 ;
      RECT  0.025000  6.560000  0.305000  6.840000 ;
      RECT  0.025000  6.960000  0.305000  7.240000 ;
      RECT  0.025000  7.360000  0.305000  7.640000 ;
      RECT  0.025000  7.760000  0.305000  8.040000 ;
      RECT  0.025000  8.160000  0.305000  8.440000 ;
      RECT  0.025000  9.170000  0.305000  9.450000 ;
      RECT  0.025000  9.570000  0.305000  9.850000 ;
      RECT  0.025000  9.970000  0.305000 10.250000 ;
      RECT  0.025000 10.370000  0.305000 10.650000 ;
      RECT  0.025000 10.770000  0.305000 11.050000 ;
      RECT  0.025000 11.170000  0.305000 11.450000 ;
      RECT  0.440000  0.025000  0.720000  0.305000 ;
      RECT  0.440000  5.785000  0.720000  6.065000 ;
      RECT  0.440000 11.545000  0.720000 11.825000 ;
      RECT  0.835000  2.905000  1.115000  3.185000 ;
      RECT  0.835000  8.665000  1.115000  8.945000 ;
      RECT  0.840000  0.025000  1.120000  0.305000 ;
      RECT  0.840000  5.785000  1.120000  6.065000 ;
      RECT  0.840000 11.545000  1.120000 11.825000 ;
      RECT  1.235000  2.905000  1.515000  3.185000 ;
      RECT  1.235000  8.665000  1.515000  8.945000 ;
      RECT  1.240000  0.025000  1.520000  0.305000 ;
      RECT  1.240000  5.785000  1.520000  6.065000 ;
      RECT  1.240000 11.545000  1.520000 11.825000 ;
      RECT  1.635000  2.905000  1.915000  3.185000 ;
      RECT  1.635000  8.665000  1.915000  8.945000 ;
      RECT  1.640000  0.025000  1.920000  0.305000 ;
      RECT  1.640000  5.785000  1.920000  6.065000 ;
      RECT  1.640000 11.545000  1.920000 11.825000 ;
      RECT  2.035000  2.905000  2.315000  3.185000 ;
      RECT  2.035000  8.665000  2.315000  8.945000 ;
      RECT  2.040000  0.025000  2.320000  0.305000 ;
      RECT  2.040000  5.785000  2.320000  6.065000 ;
      RECT  2.040000 11.545000  2.320000 11.825000 ;
      RECT  2.435000  2.905000  2.715000  3.185000 ;
      RECT  2.435000  8.665000  2.715000  8.945000 ;
      RECT  2.440000  0.025000  2.720000  0.305000 ;
      RECT  2.440000  5.785000  2.720000  6.065000 ;
      RECT  2.440000 11.545000  2.720000 11.825000 ;
      RECT  2.835000  2.905000  3.115000  3.185000 ;
      RECT  2.835000  8.665000  3.115000  8.945000 ;
      RECT  3.255000  0.705000  3.535000  0.985000 ;
      RECT  3.255000  1.105000  3.535000  1.385000 ;
      RECT  3.255000  1.505000  3.535000  1.785000 ;
      RECT  3.255000  1.905000  3.535000  2.185000 ;
      RECT  3.255000  2.305000  3.535000  2.585000 ;
      RECT  3.255000  3.505000  3.535000  3.785000 ;
      RECT  3.255000  3.905000  3.535000  4.185000 ;
      RECT  3.255000  4.305000  3.535000  4.585000 ;
      RECT  3.255000  4.705000  3.535000  4.985000 ;
      RECT  3.255000  5.105000  3.535000  5.385000 ;
      RECT  3.255000  6.465000  3.535000  6.745000 ;
      RECT  3.255000  6.865000  3.535000  7.145000 ;
      RECT  3.255000  7.265000  3.535000  7.545000 ;
      RECT  3.255000  7.665000  3.535000  7.945000 ;
      RECT  3.255000  8.065000  3.535000  8.345000 ;
      RECT  3.255000  9.265000  3.535000  9.545000 ;
      RECT  3.255000  9.665000  3.535000  9.945000 ;
      RECT  3.255000 10.065000  3.535000 10.345000 ;
      RECT  3.255000 10.465000  3.535000 10.745000 ;
      RECT  3.255000 10.865000  3.535000 11.145000 ;
      RECT  3.260000  2.905000  3.540000  3.185000 ;
      RECT  3.260000  8.665000  3.540000  8.945000 ;
      RECT  3.685000  2.905000  3.965000  3.185000 ;
      RECT  3.685000  8.665000  3.965000  8.945000 ;
      RECT  4.085000  2.905000  4.365000  3.185000 ;
      RECT  4.085000  8.665000  4.365000  8.945000 ;
      RECT  4.090000  0.025000  4.370000  0.305000 ;
      RECT  4.090000  5.785000  4.370000  6.065000 ;
      RECT  4.090000 11.545000  4.370000 11.825000 ;
      RECT  4.485000  2.905000  4.765000  3.185000 ;
      RECT  4.485000  8.665000  4.765000  8.945000 ;
      RECT  4.490000  0.025000  4.770000  0.305000 ;
      RECT  4.490000  5.785000  4.770000  6.065000 ;
      RECT  4.490000 11.545000  4.770000 11.825000 ;
      RECT  4.885000  2.905000  5.165000  3.185000 ;
      RECT  4.885000  8.665000  5.165000  8.945000 ;
      RECT  4.890000  0.025000  5.170000  0.305000 ;
      RECT  4.890000  5.785000  5.170000  6.065000 ;
      RECT  4.890000 11.545000  5.170000 11.825000 ;
      RECT  5.285000  2.905000  5.565000  3.185000 ;
      RECT  5.285000  8.665000  5.565000  8.945000 ;
      RECT  5.290000  0.025000  5.570000  0.305000 ;
      RECT  5.290000  5.785000  5.570000  6.065000 ;
      RECT  5.290000 11.545000  5.570000 11.825000 ;
      RECT  5.685000  2.905000  5.965000  3.185000 ;
      RECT  5.685000  8.665000  5.965000  8.945000 ;
      RECT  5.690000  0.025000  5.970000  0.305000 ;
      RECT  5.690000  5.785000  5.970000  6.065000 ;
      RECT  5.690000 11.545000  5.970000 11.825000 ;
      RECT  6.090000  0.025000  6.370000  0.305000 ;
      RECT  6.090000  5.785000  6.370000  6.065000 ;
      RECT  6.090000 11.545000  6.370000 11.825000 ;
      RECT  6.495000  0.400000  6.775000  0.680000 ;
      RECT  6.495000  0.800000  6.775000  1.080000 ;
      RECT  6.495000  1.200000  6.775000  1.480000 ;
      RECT  6.495000  1.600000  6.775000  1.880000 ;
      RECT  6.495000  2.000000  6.775000  2.280000 ;
      RECT  6.495000  2.400000  6.775000  2.680000 ;
      RECT  6.495000  3.410000  6.775000  3.690000 ;
      RECT  6.495000  3.810000  6.775000  4.090000 ;
      RECT  6.495000  4.210000  6.775000  4.490000 ;
      RECT  6.495000  4.610000  6.775000  4.890000 ;
      RECT  6.495000  5.010000  6.775000  5.290000 ;
      RECT  6.495000  5.410000  6.775000  5.690000 ;
      RECT  6.495000  6.160000  6.775000  6.440000 ;
      RECT  6.495000  6.560000  6.775000  6.840000 ;
      RECT  6.495000  6.960000  6.775000  7.240000 ;
      RECT  6.495000  7.360000  6.775000  7.640000 ;
      RECT  6.495000  7.760000  6.775000  8.040000 ;
      RECT  6.495000  8.160000  6.775000  8.440000 ;
      RECT  6.495000  9.170000  6.775000  9.450000 ;
      RECT  6.495000  9.570000  6.775000  9.850000 ;
      RECT  6.495000  9.970000  6.775000 10.250000 ;
      RECT  6.495000 10.370000  6.775000 10.650000 ;
      RECT  6.495000 10.770000  6.775000 11.050000 ;
      RECT  6.495000 11.170000  6.775000 11.450000 ;
      RECT  6.910000  0.025000  7.190000  0.305000 ;
      RECT  6.910000  5.785000  7.190000  6.065000 ;
      RECT  6.910000 11.545000  7.190000 11.825000 ;
      RECT  7.305000  2.905000  7.585000  3.185000 ;
      RECT  7.305000  8.665000  7.585000  8.945000 ;
      RECT  7.310000  0.025000  7.590000  0.305000 ;
      RECT  7.310000  5.785000  7.590000  6.065000 ;
      RECT  7.310000 11.545000  7.590000 11.825000 ;
      RECT  7.705000  2.905000  7.985000  3.185000 ;
      RECT  7.705000  8.665000  7.985000  8.945000 ;
      RECT  7.710000  0.025000  7.990000  0.305000 ;
      RECT  7.710000  5.785000  7.990000  6.065000 ;
      RECT  7.710000 11.545000  7.990000 11.825000 ;
      RECT  8.105000  2.905000  8.385000  3.185000 ;
      RECT  8.105000  8.665000  8.385000  8.945000 ;
      RECT  8.110000  0.025000  8.390000  0.305000 ;
      RECT  8.110000  5.785000  8.390000  6.065000 ;
      RECT  8.110000 11.545000  8.390000 11.825000 ;
      RECT  8.505000  2.905000  8.785000  3.185000 ;
      RECT  8.505000  8.665000  8.785000  8.945000 ;
      RECT  8.510000  0.025000  8.790000  0.305000 ;
      RECT  8.510000  5.785000  8.790000  6.065000 ;
      RECT  8.510000 11.545000  8.790000 11.825000 ;
      RECT  8.905000  2.905000  9.185000  3.185000 ;
      RECT  8.905000  8.665000  9.185000  8.945000 ;
      RECT  8.910000  0.025000  9.190000  0.305000 ;
      RECT  8.910000  5.785000  9.190000  6.065000 ;
      RECT  8.910000 11.545000  9.190000 11.825000 ;
      RECT  9.305000  2.905000  9.585000  3.185000 ;
      RECT  9.305000  8.665000  9.585000  8.945000 ;
      RECT  9.725000  0.705000 10.005000  0.985000 ;
      RECT  9.725000  1.105000 10.005000  1.385000 ;
      RECT  9.725000  1.505000 10.005000  1.785000 ;
      RECT  9.725000  1.905000 10.005000  2.185000 ;
      RECT  9.725000  2.305000 10.005000  2.585000 ;
      RECT  9.725000  3.505000 10.005000  3.785000 ;
      RECT  9.725000  3.905000 10.005000  4.185000 ;
      RECT  9.725000  4.305000 10.005000  4.585000 ;
      RECT  9.725000  4.705000 10.005000  4.985000 ;
      RECT  9.725000  5.105000 10.005000  5.385000 ;
      RECT  9.725000  6.465000 10.005000  6.745000 ;
      RECT  9.725000  6.865000 10.005000  7.145000 ;
      RECT  9.725000  7.265000 10.005000  7.545000 ;
      RECT  9.725000  7.665000 10.005000  7.945000 ;
      RECT  9.725000  8.065000 10.005000  8.345000 ;
      RECT  9.725000  9.265000 10.005000  9.545000 ;
      RECT  9.725000  9.665000 10.005000  9.945000 ;
      RECT  9.725000 10.065000 10.005000 10.345000 ;
      RECT  9.725000 10.465000 10.005000 10.745000 ;
      RECT  9.725000 10.865000 10.005000 11.145000 ;
      RECT  9.730000  2.905000 10.010000  3.185000 ;
      RECT  9.730000  8.665000 10.010000  8.945000 ;
      RECT 10.155000  2.905000 10.435000  3.185000 ;
      RECT 10.155000  8.665000 10.435000  8.945000 ;
      RECT 10.555000  2.905000 10.835000  3.185000 ;
      RECT 10.555000  8.665000 10.835000  8.945000 ;
      RECT 10.560000  0.025000 10.840000  0.305000 ;
      RECT 10.560000  5.785000 10.840000  6.065000 ;
      RECT 10.560000 11.545000 10.840000 11.825000 ;
      RECT 10.955000  2.905000 11.235000  3.185000 ;
      RECT 10.955000  8.665000 11.235000  8.945000 ;
      RECT 10.960000  0.025000 11.240000  0.305000 ;
      RECT 10.960000  5.785000 11.240000  6.065000 ;
      RECT 10.960000 11.545000 11.240000 11.825000 ;
      RECT 11.355000  2.905000 11.635000  3.185000 ;
      RECT 11.355000  8.665000 11.635000  8.945000 ;
      RECT 11.360000  0.025000 11.640000  0.305000 ;
      RECT 11.360000  5.785000 11.640000  6.065000 ;
      RECT 11.360000 11.545000 11.640000 11.825000 ;
      RECT 11.755000  2.905000 12.035000  3.185000 ;
      RECT 11.755000  8.665000 12.035000  8.945000 ;
      RECT 11.760000  0.025000 12.040000  0.305000 ;
      RECT 11.760000  5.785000 12.040000  6.065000 ;
      RECT 11.760000 11.545000 12.040000 11.825000 ;
      RECT 12.155000  2.905000 12.435000  3.185000 ;
      RECT 12.155000  8.665000 12.435000  8.945000 ;
      RECT 12.160000  0.025000 12.440000  0.305000 ;
      RECT 12.160000  5.785000 12.440000  6.065000 ;
      RECT 12.160000 11.545000 12.440000 11.825000 ;
      RECT 12.560000  0.025000 12.840000  0.305000 ;
      RECT 12.560000  5.785000 12.840000  6.065000 ;
      RECT 12.560000 11.545000 12.840000 11.825000 ;
      RECT 12.965000  0.400000 13.245000  0.680000 ;
      RECT 12.965000  0.800000 13.245000  1.080000 ;
      RECT 12.965000  1.200000 13.245000  1.480000 ;
      RECT 12.965000  1.600000 13.245000  1.880000 ;
      RECT 12.965000  2.000000 13.245000  2.280000 ;
      RECT 12.965000  2.400000 13.245000  2.680000 ;
      RECT 12.965000  3.410000 13.245000  3.690000 ;
      RECT 12.965000  3.810000 13.245000  4.090000 ;
      RECT 12.965000  4.210000 13.245000  4.490000 ;
      RECT 12.965000  4.610000 13.245000  4.890000 ;
      RECT 12.965000  5.010000 13.245000  5.290000 ;
      RECT 12.965000  5.410000 13.245000  5.690000 ;
      RECT 12.965000  6.160000 13.245000  6.440000 ;
      RECT 12.965000  6.560000 13.245000  6.840000 ;
      RECT 12.965000  6.960000 13.245000  7.240000 ;
      RECT 12.965000  7.360000 13.245000  7.640000 ;
      RECT 12.965000  7.760000 13.245000  8.040000 ;
      RECT 12.965000  8.160000 13.245000  8.440000 ;
      RECT 12.965000  9.170000 13.245000  9.450000 ;
      RECT 12.965000  9.570000 13.245000  9.850000 ;
      RECT 12.965000  9.970000 13.245000 10.250000 ;
      RECT 12.965000 10.370000 13.245000 10.650000 ;
      RECT 12.965000 10.770000 13.245000 11.050000 ;
      RECT 12.965000 11.170000 13.245000 11.450000 ;
  END
END sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4_top
END LIBRARY
