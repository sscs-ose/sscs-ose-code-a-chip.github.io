MACRO NMOS_S_12565100_X2_Y74
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_12565100_X2_Y74 0 0 ;
  SIZE 3440 BY 436800 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 429820 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 4460 1860 434020 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 680 2290 436120 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 144985 ;
    LAYER M1 ;
      RECT 1165 145235 1415 146245 ;
    LAYER M1 ;
      RECT 1165 147335 1415 150865 ;
    LAYER M1 ;
      RECT 1165 151115 1415 152125 ;
    LAYER M1 ;
      RECT 1165 153215 1415 156745 ;
    LAYER M1 ;
      RECT 1165 156995 1415 158005 ;
    LAYER M1 ;
      RECT 1165 159095 1415 162625 ;
    LAYER M1 ;
      RECT 1165 162875 1415 163885 ;
    LAYER M1 ;
      RECT 1165 164975 1415 168505 ;
    LAYER M1 ;
      RECT 1165 168755 1415 169765 ;
    LAYER M1 ;
      RECT 1165 170855 1415 174385 ;
    LAYER M1 ;
      RECT 1165 174635 1415 175645 ;
    LAYER M1 ;
      RECT 1165 176735 1415 180265 ;
    LAYER M1 ;
      RECT 1165 180515 1415 181525 ;
    LAYER M1 ;
      RECT 1165 182615 1415 186145 ;
    LAYER M1 ;
      RECT 1165 186395 1415 187405 ;
    LAYER M1 ;
      RECT 1165 188495 1415 192025 ;
    LAYER M1 ;
      RECT 1165 192275 1415 193285 ;
    LAYER M1 ;
      RECT 1165 194375 1415 197905 ;
    LAYER M1 ;
      RECT 1165 198155 1415 199165 ;
    LAYER M1 ;
      RECT 1165 200255 1415 203785 ;
    LAYER M1 ;
      RECT 1165 204035 1415 205045 ;
    LAYER M1 ;
      RECT 1165 206135 1415 209665 ;
    LAYER M1 ;
      RECT 1165 209915 1415 210925 ;
    LAYER M1 ;
      RECT 1165 212015 1415 215545 ;
    LAYER M1 ;
      RECT 1165 215795 1415 216805 ;
    LAYER M1 ;
      RECT 1165 217895 1415 221425 ;
    LAYER M1 ;
      RECT 1165 221675 1415 222685 ;
    LAYER M1 ;
      RECT 1165 223775 1415 227305 ;
    LAYER M1 ;
      RECT 1165 227555 1415 228565 ;
    LAYER M1 ;
      RECT 1165 229655 1415 233185 ;
    LAYER M1 ;
      RECT 1165 233435 1415 234445 ;
    LAYER M1 ;
      RECT 1165 235535 1415 239065 ;
    LAYER M1 ;
      RECT 1165 239315 1415 240325 ;
    LAYER M1 ;
      RECT 1165 241415 1415 244945 ;
    LAYER M1 ;
      RECT 1165 245195 1415 246205 ;
    LAYER M1 ;
      RECT 1165 247295 1415 250825 ;
    LAYER M1 ;
      RECT 1165 251075 1415 252085 ;
    LAYER M1 ;
      RECT 1165 253175 1415 256705 ;
    LAYER M1 ;
      RECT 1165 256955 1415 257965 ;
    LAYER M1 ;
      RECT 1165 259055 1415 262585 ;
    LAYER M1 ;
      RECT 1165 262835 1415 263845 ;
    LAYER M1 ;
      RECT 1165 264935 1415 268465 ;
    LAYER M1 ;
      RECT 1165 268715 1415 269725 ;
    LAYER M1 ;
      RECT 1165 270815 1415 274345 ;
    LAYER M1 ;
      RECT 1165 274595 1415 275605 ;
    LAYER M1 ;
      RECT 1165 276695 1415 280225 ;
    LAYER M1 ;
      RECT 1165 280475 1415 281485 ;
    LAYER M1 ;
      RECT 1165 282575 1415 286105 ;
    LAYER M1 ;
      RECT 1165 286355 1415 287365 ;
    LAYER M1 ;
      RECT 1165 288455 1415 291985 ;
    LAYER M1 ;
      RECT 1165 292235 1415 293245 ;
    LAYER M1 ;
      RECT 1165 294335 1415 297865 ;
    LAYER M1 ;
      RECT 1165 298115 1415 299125 ;
    LAYER M1 ;
      RECT 1165 300215 1415 303745 ;
    LAYER M1 ;
      RECT 1165 303995 1415 305005 ;
    LAYER M1 ;
      RECT 1165 306095 1415 309625 ;
    LAYER M1 ;
      RECT 1165 309875 1415 310885 ;
    LAYER M1 ;
      RECT 1165 311975 1415 315505 ;
    LAYER M1 ;
      RECT 1165 315755 1415 316765 ;
    LAYER M1 ;
      RECT 1165 317855 1415 321385 ;
    LAYER M1 ;
      RECT 1165 321635 1415 322645 ;
    LAYER M1 ;
      RECT 1165 323735 1415 327265 ;
    LAYER M1 ;
      RECT 1165 327515 1415 328525 ;
    LAYER M1 ;
      RECT 1165 329615 1415 333145 ;
    LAYER M1 ;
      RECT 1165 333395 1415 334405 ;
    LAYER M1 ;
      RECT 1165 335495 1415 339025 ;
    LAYER M1 ;
      RECT 1165 339275 1415 340285 ;
    LAYER M1 ;
      RECT 1165 341375 1415 344905 ;
    LAYER M1 ;
      RECT 1165 345155 1415 346165 ;
    LAYER M1 ;
      RECT 1165 347255 1415 350785 ;
    LAYER M1 ;
      RECT 1165 351035 1415 352045 ;
    LAYER M1 ;
      RECT 1165 353135 1415 356665 ;
    LAYER M1 ;
      RECT 1165 356915 1415 357925 ;
    LAYER M1 ;
      RECT 1165 359015 1415 362545 ;
    LAYER M1 ;
      RECT 1165 362795 1415 363805 ;
    LAYER M1 ;
      RECT 1165 364895 1415 368425 ;
    LAYER M1 ;
      RECT 1165 368675 1415 369685 ;
    LAYER M1 ;
      RECT 1165 370775 1415 374305 ;
    LAYER M1 ;
      RECT 1165 374555 1415 375565 ;
    LAYER M1 ;
      RECT 1165 376655 1415 380185 ;
    LAYER M1 ;
      RECT 1165 380435 1415 381445 ;
    LAYER M1 ;
      RECT 1165 382535 1415 386065 ;
    LAYER M1 ;
      RECT 1165 386315 1415 387325 ;
    LAYER M1 ;
      RECT 1165 388415 1415 391945 ;
    LAYER M1 ;
      RECT 1165 392195 1415 393205 ;
    LAYER M1 ;
      RECT 1165 394295 1415 397825 ;
    LAYER M1 ;
      RECT 1165 398075 1415 399085 ;
    LAYER M1 ;
      RECT 1165 400175 1415 403705 ;
    LAYER M1 ;
      RECT 1165 403955 1415 404965 ;
    LAYER M1 ;
      RECT 1165 406055 1415 409585 ;
    LAYER M1 ;
      RECT 1165 409835 1415 410845 ;
    LAYER M1 ;
      RECT 1165 411935 1415 415465 ;
    LAYER M1 ;
      RECT 1165 415715 1415 416725 ;
    LAYER M1 ;
      RECT 1165 417815 1415 421345 ;
    LAYER M1 ;
      RECT 1165 421595 1415 422605 ;
    LAYER M1 ;
      RECT 1165 423695 1415 427225 ;
    LAYER M1 ;
      RECT 1165 427475 1415 428485 ;
    LAYER M1 ;
      RECT 1165 429575 1415 433105 ;
    LAYER M1 ;
      RECT 1165 433355 1415 434365 ;
    LAYER M1 ;
      RECT 1165 435455 1415 436465 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 735 141455 985 144985 ;
    LAYER M1 ;
      RECT 735 147335 985 150865 ;
    LAYER M1 ;
      RECT 735 153215 985 156745 ;
    LAYER M1 ;
      RECT 735 159095 985 162625 ;
    LAYER M1 ;
      RECT 735 164975 985 168505 ;
    LAYER M1 ;
      RECT 735 170855 985 174385 ;
    LAYER M1 ;
      RECT 735 176735 985 180265 ;
    LAYER M1 ;
      RECT 735 182615 985 186145 ;
    LAYER M1 ;
      RECT 735 188495 985 192025 ;
    LAYER M1 ;
      RECT 735 194375 985 197905 ;
    LAYER M1 ;
      RECT 735 200255 985 203785 ;
    LAYER M1 ;
      RECT 735 206135 985 209665 ;
    LAYER M1 ;
      RECT 735 212015 985 215545 ;
    LAYER M1 ;
      RECT 735 217895 985 221425 ;
    LAYER M1 ;
      RECT 735 223775 985 227305 ;
    LAYER M1 ;
      RECT 735 229655 985 233185 ;
    LAYER M1 ;
      RECT 735 235535 985 239065 ;
    LAYER M1 ;
      RECT 735 241415 985 244945 ;
    LAYER M1 ;
      RECT 735 247295 985 250825 ;
    LAYER M1 ;
      RECT 735 253175 985 256705 ;
    LAYER M1 ;
      RECT 735 259055 985 262585 ;
    LAYER M1 ;
      RECT 735 264935 985 268465 ;
    LAYER M1 ;
      RECT 735 270815 985 274345 ;
    LAYER M1 ;
      RECT 735 276695 985 280225 ;
    LAYER M1 ;
      RECT 735 282575 985 286105 ;
    LAYER M1 ;
      RECT 735 288455 985 291985 ;
    LAYER M1 ;
      RECT 735 294335 985 297865 ;
    LAYER M1 ;
      RECT 735 300215 985 303745 ;
    LAYER M1 ;
      RECT 735 306095 985 309625 ;
    LAYER M1 ;
      RECT 735 311975 985 315505 ;
    LAYER M1 ;
      RECT 735 317855 985 321385 ;
    LAYER M1 ;
      RECT 735 323735 985 327265 ;
    LAYER M1 ;
      RECT 735 329615 985 333145 ;
    LAYER M1 ;
      RECT 735 335495 985 339025 ;
    LAYER M1 ;
      RECT 735 341375 985 344905 ;
    LAYER M1 ;
      RECT 735 347255 985 350785 ;
    LAYER M1 ;
      RECT 735 353135 985 356665 ;
    LAYER M1 ;
      RECT 735 359015 985 362545 ;
    LAYER M1 ;
      RECT 735 364895 985 368425 ;
    LAYER M1 ;
      RECT 735 370775 985 374305 ;
    LAYER M1 ;
      RECT 735 376655 985 380185 ;
    LAYER M1 ;
      RECT 735 382535 985 386065 ;
    LAYER M1 ;
      RECT 735 388415 985 391945 ;
    LAYER M1 ;
      RECT 735 394295 985 397825 ;
    LAYER M1 ;
      RECT 735 400175 985 403705 ;
    LAYER M1 ;
      RECT 735 406055 985 409585 ;
    LAYER M1 ;
      RECT 735 411935 985 415465 ;
    LAYER M1 ;
      RECT 735 417815 985 421345 ;
    LAYER M1 ;
      RECT 735 423695 985 427225 ;
    LAYER M1 ;
      RECT 735 429575 985 433105 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 1595 141455 1845 144985 ;
    LAYER M1 ;
      RECT 1595 147335 1845 150865 ;
    LAYER M1 ;
      RECT 1595 153215 1845 156745 ;
    LAYER M1 ;
      RECT 1595 159095 1845 162625 ;
    LAYER M1 ;
      RECT 1595 164975 1845 168505 ;
    LAYER M1 ;
      RECT 1595 170855 1845 174385 ;
    LAYER M1 ;
      RECT 1595 176735 1845 180265 ;
    LAYER M1 ;
      RECT 1595 182615 1845 186145 ;
    LAYER M1 ;
      RECT 1595 188495 1845 192025 ;
    LAYER M1 ;
      RECT 1595 194375 1845 197905 ;
    LAYER M1 ;
      RECT 1595 200255 1845 203785 ;
    LAYER M1 ;
      RECT 1595 206135 1845 209665 ;
    LAYER M1 ;
      RECT 1595 212015 1845 215545 ;
    LAYER M1 ;
      RECT 1595 217895 1845 221425 ;
    LAYER M1 ;
      RECT 1595 223775 1845 227305 ;
    LAYER M1 ;
      RECT 1595 229655 1845 233185 ;
    LAYER M1 ;
      RECT 1595 235535 1845 239065 ;
    LAYER M1 ;
      RECT 1595 241415 1845 244945 ;
    LAYER M1 ;
      RECT 1595 247295 1845 250825 ;
    LAYER M1 ;
      RECT 1595 253175 1845 256705 ;
    LAYER M1 ;
      RECT 1595 259055 1845 262585 ;
    LAYER M1 ;
      RECT 1595 264935 1845 268465 ;
    LAYER M1 ;
      RECT 1595 270815 1845 274345 ;
    LAYER M1 ;
      RECT 1595 276695 1845 280225 ;
    LAYER M1 ;
      RECT 1595 282575 1845 286105 ;
    LAYER M1 ;
      RECT 1595 288455 1845 291985 ;
    LAYER M1 ;
      RECT 1595 294335 1845 297865 ;
    LAYER M1 ;
      RECT 1595 300215 1845 303745 ;
    LAYER M1 ;
      RECT 1595 306095 1845 309625 ;
    LAYER M1 ;
      RECT 1595 311975 1845 315505 ;
    LAYER M1 ;
      RECT 1595 317855 1845 321385 ;
    LAYER M1 ;
      RECT 1595 323735 1845 327265 ;
    LAYER M1 ;
      RECT 1595 329615 1845 333145 ;
    LAYER M1 ;
      RECT 1595 335495 1845 339025 ;
    LAYER M1 ;
      RECT 1595 341375 1845 344905 ;
    LAYER M1 ;
      RECT 1595 347255 1845 350785 ;
    LAYER M1 ;
      RECT 1595 353135 1845 356665 ;
    LAYER M1 ;
      RECT 1595 359015 1845 362545 ;
    LAYER M1 ;
      RECT 1595 364895 1845 368425 ;
    LAYER M1 ;
      RECT 1595 370775 1845 374305 ;
    LAYER M1 ;
      RECT 1595 376655 1845 380185 ;
    LAYER M1 ;
      RECT 1595 382535 1845 386065 ;
    LAYER M1 ;
      RECT 1595 388415 1845 391945 ;
    LAYER M1 ;
      RECT 1595 394295 1845 397825 ;
    LAYER M1 ;
      RECT 1595 400175 1845 403705 ;
    LAYER M1 ;
      RECT 1595 406055 1845 409585 ;
    LAYER M1 ;
      RECT 1595 411935 1845 415465 ;
    LAYER M1 ;
      RECT 1595 417815 1845 421345 ;
    LAYER M1 ;
      RECT 1595 423695 1845 427225 ;
    LAYER M1 ;
      RECT 1595 429575 1845 433105 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 68545 ;
    LAYER M1 ;
      RECT 2025 68795 2275 69805 ;
    LAYER M1 ;
      RECT 2025 70895 2275 74425 ;
    LAYER M1 ;
      RECT 2025 74675 2275 75685 ;
    LAYER M1 ;
      RECT 2025 76775 2275 80305 ;
    LAYER M1 ;
      RECT 2025 80555 2275 81565 ;
    LAYER M1 ;
      RECT 2025 82655 2275 86185 ;
    LAYER M1 ;
      RECT 2025 86435 2275 87445 ;
    LAYER M1 ;
      RECT 2025 88535 2275 92065 ;
    LAYER M1 ;
      RECT 2025 92315 2275 93325 ;
    LAYER M1 ;
      RECT 2025 94415 2275 97945 ;
    LAYER M1 ;
      RECT 2025 98195 2275 99205 ;
    LAYER M1 ;
      RECT 2025 100295 2275 103825 ;
    LAYER M1 ;
      RECT 2025 104075 2275 105085 ;
    LAYER M1 ;
      RECT 2025 106175 2275 109705 ;
    LAYER M1 ;
      RECT 2025 109955 2275 110965 ;
    LAYER M1 ;
      RECT 2025 112055 2275 115585 ;
    LAYER M1 ;
      RECT 2025 115835 2275 116845 ;
    LAYER M1 ;
      RECT 2025 117935 2275 121465 ;
    LAYER M1 ;
      RECT 2025 121715 2275 122725 ;
    LAYER M1 ;
      RECT 2025 123815 2275 127345 ;
    LAYER M1 ;
      RECT 2025 127595 2275 128605 ;
    LAYER M1 ;
      RECT 2025 129695 2275 133225 ;
    LAYER M1 ;
      RECT 2025 133475 2275 134485 ;
    LAYER M1 ;
      RECT 2025 135575 2275 139105 ;
    LAYER M1 ;
      RECT 2025 139355 2275 140365 ;
    LAYER M1 ;
      RECT 2025 141455 2275 144985 ;
    LAYER M1 ;
      RECT 2025 145235 2275 146245 ;
    LAYER M1 ;
      RECT 2025 147335 2275 150865 ;
    LAYER M1 ;
      RECT 2025 151115 2275 152125 ;
    LAYER M1 ;
      RECT 2025 153215 2275 156745 ;
    LAYER M1 ;
      RECT 2025 156995 2275 158005 ;
    LAYER M1 ;
      RECT 2025 159095 2275 162625 ;
    LAYER M1 ;
      RECT 2025 162875 2275 163885 ;
    LAYER M1 ;
      RECT 2025 164975 2275 168505 ;
    LAYER M1 ;
      RECT 2025 168755 2275 169765 ;
    LAYER M1 ;
      RECT 2025 170855 2275 174385 ;
    LAYER M1 ;
      RECT 2025 174635 2275 175645 ;
    LAYER M1 ;
      RECT 2025 176735 2275 180265 ;
    LAYER M1 ;
      RECT 2025 180515 2275 181525 ;
    LAYER M1 ;
      RECT 2025 182615 2275 186145 ;
    LAYER M1 ;
      RECT 2025 186395 2275 187405 ;
    LAYER M1 ;
      RECT 2025 188495 2275 192025 ;
    LAYER M1 ;
      RECT 2025 192275 2275 193285 ;
    LAYER M1 ;
      RECT 2025 194375 2275 197905 ;
    LAYER M1 ;
      RECT 2025 198155 2275 199165 ;
    LAYER M1 ;
      RECT 2025 200255 2275 203785 ;
    LAYER M1 ;
      RECT 2025 204035 2275 205045 ;
    LAYER M1 ;
      RECT 2025 206135 2275 209665 ;
    LAYER M1 ;
      RECT 2025 209915 2275 210925 ;
    LAYER M1 ;
      RECT 2025 212015 2275 215545 ;
    LAYER M1 ;
      RECT 2025 215795 2275 216805 ;
    LAYER M1 ;
      RECT 2025 217895 2275 221425 ;
    LAYER M1 ;
      RECT 2025 221675 2275 222685 ;
    LAYER M1 ;
      RECT 2025 223775 2275 227305 ;
    LAYER M1 ;
      RECT 2025 227555 2275 228565 ;
    LAYER M1 ;
      RECT 2025 229655 2275 233185 ;
    LAYER M1 ;
      RECT 2025 233435 2275 234445 ;
    LAYER M1 ;
      RECT 2025 235535 2275 239065 ;
    LAYER M1 ;
      RECT 2025 239315 2275 240325 ;
    LAYER M1 ;
      RECT 2025 241415 2275 244945 ;
    LAYER M1 ;
      RECT 2025 245195 2275 246205 ;
    LAYER M1 ;
      RECT 2025 247295 2275 250825 ;
    LAYER M1 ;
      RECT 2025 251075 2275 252085 ;
    LAYER M1 ;
      RECT 2025 253175 2275 256705 ;
    LAYER M1 ;
      RECT 2025 256955 2275 257965 ;
    LAYER M1 ;
      RECT 2025 259055 2275 262585 ;
    LAYER M1 ;
      RECT 2025 262835 2275 263845 ;
    LAYER M1 ;
      RECT 2025 264935 2275 268465 ;
    LAYER M1 ;
      RECT 2025 268715 2275 269725 ;
    LAYER M1 ;
      RECT 2025 270815 2275 274345 ;
    LAYER M1 ;
      RECT 2025 274595 2275 275605 ;
    LAYER M1 ;
      RECT 2025 276695 2275 280225 ;
    LAYER M1 ;
      RECT 2025 280475 2275 281485 ;
    LAYER M1 ;
      RECT 2025 282575 2275 286105 ;
    LAYER M1 ;
      RECT 2025 286355 2275 287365 ;
    LAYER M1 ;
      RECT 2025 288455 2275 291985 ;
    LAYER M1 ;
      RECT 2025 292235 2275 293245 ;
    LAYER M1 ;
      RECT 2025 294335 2275 297865 ;
    LAYER M1 ;
      RECT 2025 298115 2275 299125 ;
    LAYER M1 ;
      RECT 2025 300215 2275 303745 ;
    LAYER M1 ;
      RECT 2025 303995 2275 305005 ;
    LAYER M1 ;
      RECT 2025 306095 2275 309625 ;
    LAYER M1 ;
      RECT 2025 309875 2275 310885 ;
    LAYER M1 ;
      RECT 2025 311975 2275 315505 ;
    LAYER M1 ;
      RECT 2025 315755 2275 316765 ;
    LAYER M1 ;
      RECT 2025 317855 2275 321385 ;
    LAYER M1 ;
      RECT 2025 321635 2275 322645 ;
    LAYER M1 ;
      RECT 2025 323735 2275 327265 ;
    LAYER M1 ;
      RECT 2025 327515 2275 328525 ;
    LAYER M1 ;
      RECT 2025 329615 2275 333145 ;
    LAYER M1 ;
      RECT 2025 333395 2275 334405 ;
    LAYER M1 ;
      RECT 2025 335495 2275 339025 ;
    LAYER M1 ;
      RECT 2025 339275 2275 340285 ;
    LAYER M1 ;
      RECT 2025 341375 2275 344905 ;
    LAYER M1 ;
      RECT 2025 345155 2275 346165 ;
    LAYER M1 ;
      RECT 2025 347255 2275 350785 ;
    LAYER M1 ;
      RECT 2025 351035 2275 352045 ;
    LAYER M1 ;
      RECT 2025 353135 2275 356665 ;
    LAYER M1 ;
      RECT 2025 356915 2275 357925 ;
    LAYER M1 ;
      RECT 2025 359015 2275 362545 ;
    LAYER M1 ;
      RECT 2025 362795 2275 363805 ;
    LAYER M1 ;
      RECT 2025 364895 2275 368425 ;
    LAYER M1 ;
      RECT 2025 368675 2275 369685 ;
    LAYER M1 ;
      RECT 2025 370775 2275 374305 ;
    LAYER M1 ;
      RECT 2025 374555 2275 375565 ;
    LAYER M1 ;
      RECT 2025 376655 2275 380185 ;
    LAYER M1 ;
      RECT 2025 380435 2275 381445 ;
    LAYER M1 ;
      RECT 2025 382535 2275 386065 ;
    LAYER M1 ;
      RECT 2025 386315 2275 387325 ;
    LAYER M1 ;
      RECT 2025 388415 2275 391945 ;
    LAYER M1 ;
      RECT 2025 392195 2275 393205 ;
    LAYER M1 ;
      RECT 2025 394295 2275 397825 ;
    LAYER M1 ;
      RECT 2025 398075 2275 399085 ;
    LAYER M1 ;
      RECT 2025 400175 2275 403705 ;
    LAYER M1 ;
      RECT 2025 403955 2275 404965 ;
    LAYER M1 ;
      RECT 2025 406055 2275 409585 ;
    LAYER M1 ;
      RECT 2025 409835 2275 410845 ;
    LAYER M1 ;
      RECT 2025 411935 2275 415465 ;
    LAYER M1 ;
      RECT 2025 415715 2275 416725 ;
    LAYER M1 ;
      RECT 2025 417815 2275 421345 ;
    LAYER M1 ;
      RECT 2025 421595 2275 422605 ;
    LAYER M1 ;
      RECT 2025 423695 2275 427225 ;
    LAYER M1 ;
      RECT 2025 427475 2275 428485 ;
    LAYER M1 ;
      RECT 2025 429575 2275 433105 ;
    LAYER M1 ;
      RECT 2025 433355 2275 434365 ;
    LAYER M1 ;
      RECT 2025 435455 2275 436465 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M1 ;
      RECT 2455 65015 2705 68545 ;
    LAYER M1 ;
      RECT 2455 70895 2705 74425 ;
    LAYER M1 ;
      RECT 2455 76775 2705 80305 ;
    LAYER M1 ;
      RECT 2455 82655 2705 86185 ;
    LAYER M1 ;
      RECT 2455 88535 2705 92065 ;
    LAYER M1 ;
      RECT 2455 94415 2705 97945 ;
    LAYER M1 ;
      RECT 2455 100295 2705 103825 ;
    LAYER M1 ;
      RECT 2455 106175 2705 109705 ;
    LAYER M1 ;
      RECT 2455 112055 2705 115585 ;
    LAYER M1 ;
      RECT 2455 117935 2705 121465 ;
    LAYER M1 ;
      RECT 2455 123815 2705 127345 ;
    LAYER M1 ;
      RECT 2455 129695 2705 133225 ;
    LAYER M1 ;
      RECT 2455 135575 2705 139105 ;
    LAYER M1 ;
      RECT 2455 141455 2705 144985 ;
    LAYER M1 ;
      RECT 2455 147335 2705 150865 ;
    LAYER M1 ;
      RECT 2455 153215 2705 156745 ;
    LAYER M1 ;
      RECT 2455 159095 2705 162625 ;
    LAYER M1 ;
      RECT 2455 164975 2705 168505 ;
    LAYER M1 ;
      RECT 2455 170855 2705 174385 ;
    LAYER M1 ;
      RECT 2455 176735 2705 180265 ;
    LAYER M1 ;
      RECT 2455 182615 2705 186145 ;
    LAYER M1 ;
      RECT 2455 188495 2705 192025 ;
    LAYER M1 ;
      RECT 2455 194375 2705 197905 ;
    LAYER M1 ;
      RECT 2455 200255 2705 203785 ;
    LAYER M1 ;
      RECT 2455 206135 2705 209665 ;
    LAYER M1 ;
      RECT 2455 212015 2705 215545 ;
    LAYER M1 ;
      RECT 2455 217895 2705 221425 ;
    LAYER M1 ;
      RECT 2455 223775 2705 227305 ;
    LAYER M1 ;
      RECT 2455 229655 2705 233185 ;
    LAYER M1 ;
      RECT 2455 235535 2705 239065 ;
    LAYER M1 ;
      RECT 2455 241415 2705 244945 ;
    LAYER M1 ;
      RECT 2455 247295 2705 250825 ;
    LAYER M1 ;
      RECT 2455 253175 2705 256705 ;
    LAYER M1 ;
      RECT 2455 259055 2705 262585 ;
    LAYER M1 ;
      RECT 2455 264935 2705 268465 ;
    LAYER M1 ;
      RECT 2455 270815 2705 274345 ;
    LAYER M1 ;
      RECT 2455 276695 2705 280225 ;
    LAYER M1 ;
      RECT 2455 282575 2705 286105 ;
    LAYER M1 ;
      RECT 2455 288455 2705 291985 ;
    LAYER M1 ;
      RECT 2455 294335 2705 297865 ;
    LAYER M1 ;
      RECT 2455 300215 2705 303745 ;
    LAYER M1 ;
      RECT 2455 306095 2705 309625 ;
    LAYER M1 ;
      RECT 2455 311975 2705 315505 ;
    LAYER M1 ;
      RECT 2455 317855 2705 321385 ;
    LAYER M1 ;
      RECT 2455 323735 2705 327265 ;
    LAYER M1 ;
      RECT 2455 329615 2705 333145 ;
    LAYER M1 ;
      RECT 2455 335495 2705 339025 ;
    LAYER M1 ;
      RECT 2455 341375 2705 344905 ;
    LAYER M1 ;
      RECT 2455 347255 2705 350785 ;
    LAYER M1 ;
      RECT 2455 353135 2705 356665 ;
    LAYER M1 ;
      RECT 2455 359015 2705 362545 ;
    LAYER M1 ;
      RECT 2455 364895 2705 368425 ;
    LAYER M1 ;
      RECT 2455 370775 2705 374305 ;
    LAYER M1 ;
      RECT 2455 376655 2705 380185 ;
    LAYER M1 ;
      RECT 2455 382535 2705 386065 ;
    LAYER M1 ;
      RECT 2455 388415 2705 391945 ;
    LAYER M1 ;
      RECT 2455 394295 2705 397825 ;
    LAYER M1 ;
      RECT 2455 400175 2705 403705 ;
    LAYER M1 ;
      RECT 2455 406055 2705 409585 ;
    LAYER M1 ;
      RECT 2455 411935 2705 415465 ;
    LAYER M1 ;
      RECT 2455 417815 2705 421345 ;
    LAYER M1 ;
      RECT 2455 423695 2705 427225 ;
    LAYER M1 ;
      RECT 2455 429575 2705 433105 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 690 700 2750 980 ;
    LAYER M2 ;
      RECT 1120 6160 2320 6440 ;
    LAYER M2 ;
      RECT 1120 10360 2320 10640 ;
    LAYER M2 ;
      RECT 690 6580 2750 6860 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 1120 16240 2320 16520 ;
    LAYER M2 ;
      RECT 690 12460 2750 12740 ;
    LAYER M2 ;
      RECT 1120 17920 2320 18200 ;
    LAYER M2 ;
      RECT 1120 22120 2320 22400 ;
    LAYER M2 ;
      RECT 690 18340 2750 18620 ;
    LAYER M2 ;
      RECT 1120 23800 2320 24080 ;
    LAYER M2 ;
      RECT 1120 28000 2320 28280 ;
    LAYER M2 ;
      RECT 690 24220 2750 24500 ;
    LAYER M2 ;
      RECT 1120 29680 2320 29960 ;
    LAYER M2 ;
      RECT 1120 33880 2320 34160 ;
    LAYER M2 ;
      RECT 690 30100 2750 30380 ;
    LAYER M2 ;
      RECT 1120 35560 2320 35840 ;
    LAYER M2 ;
      RECT 1120 39760 2320 40040 ;
    LAYER M2 ;
      RECT 690 35980 2750 36260 ;
    LAYER M2 ;
      RECT 1120 41440 2320 41720 ;
    LAYER M2 ;
      RECT 1120 45640 2320 45920 ;
    LAYER M2 ;
      RECT 690 41860 2750 42140 ;
    LAYER M2 ;
      RECT 1120 47320 2320 47600 ;
    LAYER M2 ;
      RECT 1120 51520 2320 51800 ;
    LAYER M2 ;
      RECT 690 47740 2750 48020 ;
    LAYER M2 ;
      RECT 1120 53200 2320 53480 ;
    LAYER M2 ;
      RECT 1120 57400 2320 57680 ;
    LAYER M2 ;
      RECT 690 53620 2750 53900 ;
    LAYER M2 ;
      RECT 1120 59080 2320 59360 ;
    LAYER M2 ;
      RECT 1120 63280 2320 63560 ;
    LAYER M2 ;
      RECT 690 59500 2750 59780 ;
    LAYER M2 ;
      RECT 1120 64960 2320 65240 ;
    LAYER M2 ;
      RECT 1120 69160 2320 69440 ;
    LAYER M2 ;
      RECT 690 65380 2750 65660 ;
    LAYER M2 ;
      RECT 1120 70840 2320 71120 ;
    LAYER M2 ;
      RECT 1120 75040 2320 75320 ;
    LAYER M2 ;
      RECT 690 71260 2750 71540 ;
    LAYER M2 ;
      RECT 1120 76720 2320 77000 ;
    LAYER M2 ;
      RECT 1120 80920 2320 81200 ;
    LAYER M2 ;
      RECT 690 77140 2750 77420 ;
    LAYER M2 ;
      RECT 1120 82600 2320 82880 ;
    LAYER M2 ;
      RECT 1120 86800 2320 87080 ;
    LAYER M2 ;
      RECT 690 83020 2750 83300 ;
    LAYER M2 ;
      RECT 1120 88480 2320 88760 ;
    LAYER M2 ;
      RECT 1120 92680 2320 92960 ;
    LAYER M2 ;
      RECT 690 88900 2750 89180 ;
    LAYER M2 ;
      RECT 1120 94360 2320 94640 ;
    LAYER M2 ;
      RECT 1120 98560 2320 98840 ;
    LAYER M2 ;
      RECT 690 94780 2750 95060 ;
    LAYER M2 ;
      RECT 1120 100240 2320 100520 ;
    LAYER M2 ;
      RECT 1120 104440 2320 104720 ;
    LAYER M2 ;
      RECT 690 100660 2750 100940 ;
    LAYER M2 ;
      RECT 1120 106120 2320 106400 ;
    LAYER M2 ;
      RECT 1120 110320 2320 110600 ;
    LAYER M2 ;
      RECT 690 106540 2750 106820 ;
    LAYER M2 ;
      RECT 1120 112000 2320 112280 ;
    LAYER M2 ;
      RECT 1120 116200 2320 116480 ;
    LAYER M2 ;
      RECT 690 112420 2750 112700 ;
    LAYER M2 ;
      RECT 1120 117880 2320 118160 ;
    LAYER M2 ;
      RECT 1120 122080 2320 122360 ;
    LAYER M2 ;
      RECT 690 118300 2750 118580 ;
    LAYER M2 ;
      RECT 1120 123760 2320 124040 ;
    LAYER M2 ;
      RECT 1120 127960 2320 128240 ;
    LAYER M2 ;
      RECT 690 124180 2750 124460 ;
    LAYER M2 ;
      RECT 1120 129640 2320 129920 ;
    LAYER M2 ;
      RECT 1120 133840 2320 134120 ;
    LAYER M2 ;
      RECT 690 130060 2750 130340 ;
    LAYER M2 ;
      RECT 1120 135520 2320 135800 ;
    LAYER M2 ;
      RECT 1120 139720 2320 140000 ;
    LAYER M2 ;
      RECT 690 135940 2750 136220 ;
    LAYER M2 ;
      RECT 1120 141400 2320 141680 ;
    LAYER M2 ;
      RECT 1120 145600 2320 145880 ;
    LAYER M2 ;
      RECT 690 141820 2750 142100 ;
    LAYER M2 ;
      RECT 1120 147280 2320 147560 ;
    LAYER M2 ;
      RECT 1120 151480 2320 151760 ;
    LAYER M2 ;
      RECT 690 147700 2750 147980 ;
    LAYER M2 ;
      RECT 1120 153160 2320 153440 ;
    LAYER M2 ;
      RECT 1120 157360 2320 157640 ;
    LAYER M2 ;
      RECT 690 153580 2750 153860 ;
    LAYER M2 ;
      RECT 1120 159040 2320 159320 ;
    LAYER M2 ;
      RECT 1120 163240 2320 163520 ;
    LAYER M2 ;
      RECT 690 159460 2750 159740 ;
    LAYER M2 ;
      RECT 1120 164920 2320 165200 ;
    LAYER M2 ;
      RECT 1120 169120 2320 169400 ;
    LAYER M2 ;
      RECT 690 165340 2750 165620 ;
    LAYER M2 ;
      RECT 1120 170800 2320 171080 ;
    LAYER M2 ;
      RECT 1120 175000 2320 175280 ;
    LAYER M2 ;
      RECT 690 171220 2750 171500 ;
    LAYER M2 ;
      RECT 1120 176680 2320 176960 ;
    LAYER M2 ;
      RECT 1120 180880 2320 181160 ;
    LAYER M2 ;
      RECT 690 177100 2750 177380 ;
    LAYER M2 ;
      RECT 1120 182560 2320 182840 ;
    LAYER M2 ;
      RECT 1120 186760 2320 187040 ;
    LAYER M2 ;
      RECT 690 182980 2750 183260 ;
    LAYER M2 ;
      RECT 1120 188440 2320 188720 ;
    LAYER M2 ;
      RECT 1120 192640 2320 192920 ;
    LAYER M2 ;
      RECT 690 188860 2750 189140 ;
    LAYER M2 ;
      RECT 1120 194320 2320 194600 ;
    LAYER M2 ;
      RECT 1120 198520 2320 198800 ;
    LAYER M2 ;
      RECT 690 194740 2750 195020 ;
    LAYER M2 ;
      RECT 1120 200200 2320 200480 ;
    LAYER M2 ;
      RECT 1120 204400 2320 204680 ;
    LAYER M2 ;
      RECT 690 200620 2750 200900 ;
    LAYER M2 ;
      RECT 1120 206080 2320 206360 ;
    LAYER M2 ;
      RECT 1120 210280 2320 210560 ;
    LAYER M2 ;
      RECT 690 206500 2750 206780 ;
    LAYER M2 ;
      RECT 1120 211960 2320 212240 ;
    LAYER M2 ;
      RECT 1120 216160 2320 216440 ;
    LAYER M2 ;
      RECT 690 212380 2750 212660 ;
    LAYER M2 ;
      RECT 1120 217840 2320 218120 ;
    LAYER M2 ;
      RECT 1120 222040 2320 222320 ;
    LAYER M2 ;
      RECT 690 218260 2750 218540 ;
    LAYER M2 ;
      RECT 1120 223720 2320 224000 ;
    LAYER M2 ;
      RECT 1120 227920 2320 228200 ;
    LAYER M2 ;
      RECT 690 224140 2750 224420 ;
    LAYER M2 ;
      RECT 1120 229600 2320 229880 ;
    LAYER M2 ;
      RECT 1120 233800 2320 234080 ;
    LAYER M2 ;
      RECT 690 230020 2750 230300 ;
    LAYER M2 ;
      RECT 1120 235480 2320 235760 ;
    LAYER M2 ;
      RECT 1120 239680 2320 239960 ;
    LAYER M2 ;
      RECT 690 235900 2750 236180 ;
    LAYER M2 ;
      RECT 1120 241360 2320 241640 ;
    LAYER M2 ;
      RECT 1120 245560 2320 245840 ;
    LAYER M2 ;
      RECT 690 241780 2750 242060 ;
    LAYER M2 ;
      RECT 1120 247240 2320 247520 ;
    LAYER M2 ;
      RECT 1120 251440 2320 251720 ;
    LAYER M2 ;
      RECT 690 247660 2750 247940 ;
    LAYER M2 ;
      RECT 1120 253120 2320 253400 ;
    LAYER M2 ;
      RECT 1120 257320 2320 257600 ;
    LAYER M2 ;
      RECT 690 253540 2750 253820 ;
    LAYER M2 ;
      RECT 1120 259000 2320 259280 ;
    LAYER M2 ;
      RECT 1120 263200 2320 263480 ;
    LAYER M2 ;
      RECT 690 259420 2750 259700 ;
    LAYER M2 ;
      RECT 1120 264880 2320 265160 ;
    LAYER M2 ;
      RECT 1120 269080 2320 269360 ;
    LAYER M2 ;
      RECT 690 265300 2750 265580 ;
    LAYER M2 ;
      RECT 1120 270760 2320 271040 ;
    LAYER M2 ;
      RECT 1120 274960 2320 275240 ;
    LAYER M2 ;
      RECT 690 271180 2750 271460 ;
    LAYER M2 ;
      RECT 1120 276640 2320 276920 ;
    LAYER M2 ;
      RECT 1120 280840 2320 281120 ;
    LAYER M2 ;
      RECT 690 277060 2750 277340 ;
    LAYER M2 ;
      RECT 1120 282520 2320 282800 ;
    LAYER M2 ;
      RECT 1120 286720 2320 287000 ;
    LAYER M2 ;
      RECT 690 282940 2750 283220 ;
    LAYER M2 ;
      RECT 1120 288400 2320 288680 ;
    LAYER M2 ;
      RECT 1120 292600 2320 292880 ;
    LAYER M2 ;
      RECT 690 288820 2750 289100 ;
    LAYER M2 ;
      RECT 1120 294280 2320 294560 ;
    LAYER M2 ;
      RECT 1120 298480 2320 298760 ;
    LAYER M2 ;
      RECT 690 294700 2750 294980 ;
    LAYER M2 ;
      RECT 1120 300160 2320 300440 ;
    LAYER M2 ;
      RECT 1120 304360 2320 304640 ;
    LAYER M2 ;
      RECT 690 300580 2750 300860 ;
    LAYER M2 ;
      RECT 1120 306040 2320 306320 ;
    LAYER M2 ;
      RECT 1120 310240 2320 310520 ;
    LAYER M2 ;
      RECT 690 306460 2750 306740 ;
    LAYER M2 ;
      RECT 1120 311920 2320 312200 ;
    LAYER M2 ;
      RECT 1120 316120 2320 316400 ;
    LAYER M2 ;
      RECT 690 312340 2750 312620 ;
    LAYER M2 ;
      RECT 1120 317800 2320 318080 ;
    LAYER M2 ;
      RECT 1120 322000 2320 322280 ;
    LAYER M2 ;
      RECT 690 318220 2750 318500 ;
    LAYER M2 ;
      RECT 1120 323680 2320 323960 ;
    LAYER M2 ;
      RECT 1120 327880 2320 328160 ;
    LAYER M2 ;
      RECT 690 324100 2750 324380 ;
    LAYER M2 ;
      RECT 1120 329560 2320 329840 ;
    LAYER M2 ;
      RECT 1120 333760 2320 334040 ;
    LAYER M2 ;
      RECT 690 329980 2750 330260 ;
    LAYER M2 ;
      RECT 1120 335440 2320 335720 ;
    LAYER M2 ;
      RECT 1120 339640 2320 339920 ;
    LAYER M2 ;
      RECT 690 335860 2750 336140 ;
    LAYER M2 ;
      RECT 1120 341320 2320 341600 ;
    LAYER M2 ;
      RECT 1120 345520 2320 345800 ;
    LAYER M2 ;
      RECT 690 341740 2750 342020 ;
    LAYER M2 ;
      RECT 1120 347200 2320 347480 ;
    LAYER M2 ;
      RECT 1120 351400 2320 351680 ;
    LAYER M2 ;
      RECT 690 347620 2750 347900 ;
    LAYER M2 ;
      RECT 1120 353080 2320 353360 ;
    LAYER M2 ;
      RECT 1120 357280 2320 357560 ;
    LAYER M2 ;
      RECT 690 353500 2750 353780 ;
    LAYER M2 ;
      RECT 1120 358960 2320 359240 ;
    LAYER M2 ;
      RECT 1120 363160 2320 363440 ;
    LAYER M2 ;
      RECT 690 359380 2750 359660 ;
    LAYER M2 ;
      RECT 1120 364840 2320 365120 ;
    LAYER M2 ;
      RECT 1120 369040 2320 369320 ;
    LAYER M2 ;
      RECT 690 365260 2750 365540 ;
    LAYER M2 ;
      RECT 1120 370720 2320 371000 ;
    LAYER M2 ;
      RECT 1120 374920 2320 375200 ;
    LAYER M2 ;
      RECT 690 371140 2750 371420 ;
    LAYER M2 ;
      RECT 1120 376600 2320 376880 ;
    LAYER M2 ;
      RECT 1120 380800 2320 381080 ;
    LAYER M2 ;
      RECT 690 377020 2750 377300 ;
    LAYER M2 ;
      RECT 1120 382480 2320 382760 ;
    LAYER M2 ;
      RECT 1120 386680 2320 386960 ;
    LAYER M2 ;
      RECT 690 382900 2750 383180 ;
    LAYER M2 ;
      RECT 1120 388360 2320 388640 ;
    LAYER M2 ;
      RECT 1120 392560 2320 392840 ;
    LAYER M2 ;
      RECT 690 388780 2750 389060 ;
    LAYER M2 ;
      RECT 1120 394240 2320 394520 ;
    LAYER M2 ;
      RECT 1120 398440 2320 398720 ;
    LAYER M2 ;
      RECT 690 394660 2750 394940 ;
    LAYER M2 ;
      RECT 1120 400120 2320 400400 ;
    LAYER M2 ;
      RECT 1120 404320 2320 404600 ;
    LAYER M2 ;
      RECT 690 400540 2750 400820 ;
    LAYER M2 ;
      RECT 1120 406000 2320 406280 ;
    LAYER M2 ;
      RECT 1120 410200 2320 410480 ;
    LAYER M2 ;
      RECT 690 406420 2750 406700 ;
    LAYER M2 ;
      RECT 1120 411880 2320 412160 ;
    LAYER M2 ;
      RECT 1120 416080 2320 416360 ;
    LAYER M2 ;
      RECT 690 412300 2750 412580 ;
    LAYER M2 ;
      RECT 1120 417760 2320 418040 ;
    LAYER M2 ;
      RECT 1120 421960 2320 422240 ;
    LAYER M2 ;
      RECT 690 418180 2750 418460 ;
    LAYER M2 ;
      RECT 1120 423640 2320 423920 ;
    LAYER M2 ;
      RECT 1120 427840 2320 428120 ;
    LAYER M2 ;
      RECT 690 424060 2750 424340 ;
    LAYER M2 ;
      RECT 1120 429520 2320 429800 ;
    LAYER M2 ;
      RECT 1120 433720 2320 434000 ;
    LAYER M2 ;
      RECT 1120 435820 2320 436100 ;
    LAYER M2 ;
      RECT 690 429940 2750 430220 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141455 1375 141625 ;
    LAYER V1 ;
      RECT 1205 145655 1375 145825 ;
    LAYER V1 ;
      RECT 1205 147335 1375 147505 ;
    LAYER V1 ;
      RECT 1205 151535 1375 151705 ;
    LAYER V1 ;
      RECT 1205 153215 1375 153385 ;
    LAYER V1 ;
      RECT 1205 157415 1375 157585 ;
    LAYER V1 ;
      RECT 1205 159095 1375 159265 ;
    LAYER V1 ;
      RECT 1205 163295 1375 163465 ;
    LAYER V1 ;
      RECT 1205 164975 1375 165145 ;
    LAYER V1 ;
      RECT 1205 169175 1375 169345 ;
    LAYER V1 ;
      RECT 1205 170855 1375 171025 ;
    LAYER V1 ;
      RECT 1205 175055 1375 175225 ;
    LAYER V1 ;
      RECT 1205 176735 1375 176905 ;
    LAYER V1 ;
      RECT 1205 180935 1375 181105 ;
    LAYER V1 ;
      RECT 1205 182615 1375 182785 ;
    LAYER V1 ;
      RECT 1205 186815 1375 186985 ;
    LAYER V1 ;
      RECT 1205 188495 1375 188665 ;
    LAYER V1 ;
      RECT 1205 192695 1375 192865 ;
    LAYER V1 ;
      RECT 1205 194375 1375 194545 ;
    LAYER V1 ;
      RECT 1205 198575 1375 198745 ;
    LAYER V1 ;
      RECT 1205 200255 1375 200425 ;
    LAYER V1 ;
      RECT 1205 204455 1375 204625 ;
    LAYER V1 ;
      RECT 1205 206135 1375 206305 ;
    LAYER V1 ;
      RECT 1205 210335 1375 210505 ;
    LAYER V1 ;
      RECT 1205 212015 1375 212185 ;
    LAYER V1 ;
      RECT 1205 216215 1375 216385 ;
    LAYER V1 ;
      RECT 1205 217895 1375 218065 ;
    LAYER V1 ;
      RECT 1205 222095 1375 222265 ;
    LAYER V1 ;
      RECT 1205 223775 1375 223945 ;
    LAYER V1 ;
      RECT 1205 227975 1375 228145 ;
    LAYER V1 ;
      RECT 1205 229655 1375 229825 ;
    LAYER V1 ;
      RECT 1205 233855 1375 234025 ;
    LAYER V1 ;
      RECT 1205 235535 1375 235705 ;
    LAYER V1 ;
      RECT 1205 239735 1375 239905 ;
    LAYER V1 ;
      RECT 1205 241415 1375 241585 ;
    LAYER V1 ;
      RECT 1205 245615 1375 245785 ;
    LAYER V1 ;
      RECT 1205 247295 1375 247465 ;
    LAYER V1 ;
      RECT 1205 251495 1375 251665 ;
    LAYER V1 ;
      RECT 1205 253175 1375 253345 ;
    LAYER V1 ;
      RECT 1205 257375 1375 257545 ;
    LAYER V1 ;
      RECT 1205 259055 1375 259225 ;
    LAYER V1 ;
      RECT 1205 263255 1375 263425 ;
    LAYER V1 ;
      RECT 1205 264935 1375 265105 ;
    LAYER V1 ;
      RECT 1205 269135 1375 269305 ;
    LAYER V1 ;
      RECT 1205 270815 1375 270985 ;
    LAYER V1 ;
      RECT 1205 275015 1375 275185 ;
    LAYER V1 ;
      RECT 1205 276695 1375 276865 ;
    LAYER V1 ;
      RECT 1205 280895 1375 281065 ;
    LAYER V1 ;
      RECT 1205 282575 1375 282745 ;
    LAYER V1 ;
      RECT 1205 286775 1375 286945 ;
    LAYER V1 ;
      RECT 1205 288455 1375 288625 ;
    LAYER V1 ;
      RECT 1205 292655 1375 292825 ;
    LAYER V1 ;
      RECT 1205 294335 1375 294505 ;
    LAYER V1 ;
      RECT 1205 298535 1375 298705 ;
    LAYER V1 ;
      RECT 1205 300215 1375 300385 ;
    LAYER V1 ;
      RECT 1205 304415 1375 304585 ;
    LAYER V1 ;
      RECT 1205 306095 1375 306265 ;
    LAYER V1 ;
      RECT 1205 310295 1375 310465 ;
    LAYER V1 ;
      RECT 1205 311975 1375 312145 ;
    LAYER V1 ;
      RECT 1205 316175 1375 316345 ;
    LAYER V1 ;
      RECT 1205 317855 1375 318025 ;
    LAYER V1 ;
      RECT 1205 322055 1375 322225 ;
    LAYER V1 ;
      RECT 1205 323735 1375 323905 ;
    LAYER V1 ;
      RECT 1205 327935 1375 328105 ;
    LAYER V1 ;
      RECT 1205 329615 1375 329785 ;
    LAYER V1 ;
      RECT 1205 333815 1375 333985 ;
    LAYER V1 ;
      RECT 1205 335495 1375 335665 ;
    LAYER V1 ;
      RECT 1205 339695 1375 339865 ;
    LAYER V1 ;
      RECT 1205 341375 1375 341545 ;
    LAYER V1 ;
      RECT 1205 345575 1375 345745 ;
    LAYER V1 ;
      RECT 1205 347255 1375 347425 ;
    LAYER V1 ;
      RECT 1205 351455 1375 351625 ;
    LAYER V1 ;
      RECT 1205 353135 1375 353305 ;
    LAYER V1 ;
      RECT 1205 357335 1375 357505 ;
    LAYER V1 ;
      RECT 1205 359015 1375 359185 ;
    LAYER V1 ;
      RECT 1205 363215 1375 363385 ;
    LAYER V1 ;
      RECT 1205 364895 1375 365065 ;
    LAYER V1 ;
      RECT 1205 369095 1375 369265 ;
    LAYER V1 ;
      RECT 1205 370775 1375 370945 ;
    LAYER V1 ;
      RECT 1205 374975 1375 375145 ;
    LAYER V1 ;
      RECT 1205 376655 1375 376825 ;
    LAYER V1 ;
      RECT 1205 380855 1375 381025 ;
    LAYER V1 ;
      RECT 1205 382535 1375 382705 ;
    LAYER V1 ;
      RECT 1205 386735 1375 386905 ;
    LAYER V1 ;
      RECT 1205 388415 1375 388585 ;
    LAYER V1 ;
      RECT 1205 392615 1375 392785 ;
    LAYER V1 ;
      RECT 1205 394295 1375 394465 ;
    LAYER V1 ;
      RECT 1205 398495 1375 398665 ;
    LAYER V1 ;
      RECT 1205 400175 1375 400345 ;
    LAYER V1 ;
      RECT 1205 404375 1375 404545 ;
    LAYER V1 ;
      RECT 1205 406055 1375 406225 ;
    LAYER V1 ;
      RECT 1205 410255 1375 410425 ;
    LAYER V1 ;
      RECT 1205 411935 1375 412105 ;
    LAYER V1 ;
      RECT 1205 416135 1375 416305 ;
    LAYER V1 ;
      RECT 1205 417815 1375 417985 ;
    LAYER V1 ;
      RECT 1205 422015 1375 422185 ;
    LAYER V1 ;
      RECT 1205 423695 1375 423865 ;
    LAYER V1 ;
      RECT 1205 427895 1375 428065 ;
    LAYER V1 ;
      RECT 1205 429575 1375 429745 ;
    LAYER V1 ;
      RECT 1205 433775 1375 433945 ;
    LAYER V1 ;
      RECT 1205 435875 1375 436045 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59135 2235 59305 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65015 2235 65185 ;
    LAYER V1 ;
      RECT 2065 69215 2235 69385 ;
    LAYER V1 ;
      RECT 2065 70895 2235 71065 ;
    LAYER V1 ;
      RECT 2065 75095 2235 75265 ;
    LAYER V1 ;
      RECT 2065 76775 2235 76945 ;
    LAYER V1 ;
      RECT 2065 80975 2235 81145 ;
    LAYER V1 ;
      RECT 2065 82655 2235 82825 ;
    LAYER V1 ;
      RECT 2065 86855 2235 87025 ;
    LAYER V1 ;
      RECT 2065 88535 2235 88705 ;
    LAYER V1 ;
      RECT 2065 92735 2235 92905 ;
    LAYER V1 ;
      RECT 2065 94415 2235 94585 ;
    LAYER V1 ;
      RECT 2065 98615 2235 98785 ;
    LAYER V1 ;
      RECT 2065 100295 2235 100465 ;
    LAYER V1 ;
      RECT 2065 104495 2235 104665 ;
    LAYER V1 ;
      RECT 2065 106175 2235 106345 ;
    LAYER V1 ;
      RECT 2065 110375 2235 110545 ;
    LAYER V1 ;
      RECT 2065 112055 2235 112225 ;
    LAYER V1 ;
      RECT 2065 116255 2235 116425 ;
    LAYER V1 ;
      RECT 2065 117935 2235 118105 ;
    LAYER V1 ;
      RECT 2065 122135 2235 122305 ;
    LAYER V1 ;
      RECT 2065 123815 2235 123985 ;
    LAYER V1 ;
      RECT 2065 128015 2235 128185 ;
    LAYER V1 ;
      RECT 2065 129695 2235 129865 ;
    LAYER V1 ;
      RECT 2065 133895 2235 134065 ;
    LAYER V1 ;
      RECT 2065 135575 2235 135745 ;
    LAYER V1 ;
      RECT 2065 139775 2235 139945 ;
    LAYER V1 ;
      RECT 2065 141455 2235 141625 ;
    LAYER V1 ;
      RECT 2065 145655 2235 145825 ;
    LAYER V1 ;
      RECT 2065 147335 2235 147505 ;
    LAYER V1 ;
      RECT 2065 151535 2235 151705 ;
    LAYER V1 ;
      RECT 2065 153215 2235 153385 ;
    LAYER V1 ;
      RECT 2065 157415 2235 157585 ;
    LAYER V1 ;
      RECT 2065 159095 2235 159265 ;
    LAYER V1 ;
      RECT 2065 163295 2235 163465 ;
    LAYER V1 ;
      RECT 2065 164975 2235 165145 ;
    LAYER V1 ;
      RECT 2065 169175 2235 169345 ;
    LAYER V1 ;
      RECT 2065 170855 2235 171025 ;
    LAYER V1 ;
      RECT 2065 175055 2235 175225 ;
    LAYER V1 ;
      RECT 2065 176735 2235 176905 ;
    LAYER V1 ;
      RECT 2065 180935 2235 181105 ;
    LAYER V1 ;
      RECT 2065 182615 2235 182785 ;
    LAYER V1 ;
      RECT 2065 186815 2235 186985 ;
    LAYER V1 ;
      RECT 2065 188495 2235 188665 ;
    LAYER V1 ;
      RECT 2065 192695 2235 192865 ;
    LAYER V1 ;
      RECT 2065 194375 2235 194545 ;
    LAYER V1 ;
      RECT 2065 198575 2235 198745 ;
    LAYER V1 ;
      RECT 2065 200255 2235 200425 ;
    LAYER V1 ;
      RECT 2065 204455 2235 204625 ;
    LAYER V1 ;
      RECT 2065 206135 2235 206305 ;
    LAYER V1 ;
      RECT 2065 210335 2235 210505 ;
    LAYER V1 ;
      RECT 2065 212015 2235 212185 ;
    LAYER V1 ;
      RECT 2065 216215 2235 216385 ;
    LAYER V1 ;
      RECT 2065 217895 2235 218065 ;
    LAYER V1 ;
      RECT 2065 222095 2235 222265 ;
    LAYER V1 ;
      RECT 2065 223775 2235 223945 ;
    LAYER V1 ;
      RECT 2065 227975 2235 228145 ;
    LAYER V1 ;
      RECT 2065 229655 2235 229825 ;
    LAYER V1 ;
      RECT 2065 233855 2235 234025 ;
    LAYER V1 ;
      RECT 2065 235535 2235 235705 ;
    LAYER V1 ;
      RECT 2065 239735 2235 239905 ;
    LAYER V1 ;
      RECT 2065 241415 2235 241585 ;
    LAYER V1 ;
      RECT 2065 245615 2235 245785 ;
    LAYER V1 ;
      RECT 2065 247295 2235 247465 ;
    LAYER V1 ;
      RECT 2065 251495 2235 251665 ;
    LAYER V1 ;
      RECT 2065 253175 2235 253345 ;
    LAYER V1 ;
      RECT 2065 257375 2235 257545 ;
    LAYER V1 ;
      RECT 2065 259055 2235 259225 ;
    LAYER V1 ;
      RECT 2065 263255 2235 263425 ;
    LAYER V1 ;
      RECT 2065 264935 2235 265105 ;
    LAYER V1 ;
      RECT 2065 269135 2235 269305 ;
    LAYER V1 ;
      RECT 2065 270815 2235 270985 ;
    LAYER V1 ;
      RECT 2065 275015 2235 275185 ;
    LAYER V1 ;
      RECT 2065 276695 2235 276865 ;
    LAYER V1 ;
      RECT 2065 280895 2235 281065 ;
    LAYER V1 ;
      RECT 2065 282575 2235 282745 ;
    LAYER V1 ;
      RECT 2065 286775 2235 286945 ;
    LAYER V1 ;
      RECT 2065 288455 2235 288625 ;
    LAYER V1 ;
      RECT 2065 292655 2235 292825 ;
    LAYER V1 ;
      RECT 2065 294335 2235 294505 ;
    LAYER V1 ;
      RECT 2065 298535 2235 298705 ;
    LAYER V1 ;
      RECT 2065 300215 2235 300385 ;
    LAYER V1 ;
      RECT 2065 304415 2235 304585 ;
    LAYER V1 ;
      RECT 2065 306095 2235 306265 ;
    LAYER V1 ;
      RECT 2065 310295 2235 310465 ;
    LAYER V1 ;
      RECT 2065 311975 2235 312145 ;
    LAYER V1 ;
      RECT 2065 316175 2235 316345 ;
    LAYER V1 ;
      RECT 2065 317855 2235 318025 ;
    LAYER V1 ;
      RECT 2065 322055 2235 322225 ;
    LAYER V1 ;
      RECT 2065 323735 2235 323905 ;
    LAYER V1 ;
      RECT 2065 327935 2235 328105 ;
    LAYER V1 ;
      RECT 2065 329615 2235 329785 ;
    LAYER V1 ;
      RECT 2065 333815 2235 333985 ;
    LAYER V1 ;
      RECT 2065 335495 2235 335665 ;
    LAYER V1 ;
      RECT 2065 339695 2235 339865 ;
    LAYER V1 ;
      RECT 2065 341375 2235 341545 ;
    LAYER V1 ;
      RECT 2065 345575 2235 345745 ;
    LAYER V1 ;
      RECT 2065 347255 2235 347425 ;
    LAYER V1 ;
      RECT 2065 351455 2235 351625 ;
    LAYER V1 ;
      RECT 2065 353135 2235 353305 ;
    LAYER V1 ;
      RECT 2065 357335 2235 357505 ;
    LAYER V1 ;
      RECT 2065 359015 2235 359185 ;
    LAYER V1 ;
      RECT 2065 363215 2235 363385 ;
    LAYER V1 ;
      RECT 2065 364895 2235 365065 ;
    LAYER V1 ;
      RECT 2065 369095 2235 369265 ;
    LAYER V1 ;
      RECT 2065 370775 2235 370945 ;
    LAYER V1 ;
      RECT 2065 374975 2235 375145 ;
    LAYER V1 ;
      RECT 2065 376655 2235 376825 ;
    LAYER V1 ;
      RECT 2065 380855 2235 381025 ;
    LAYER V1 ;
      RECT 2065 382535 2235 382705 ;
    LAYER V1 ;
      RECT 2065 386735 2235 386905 ;
    LAYER V1 ;
      RECT 2065 388415 2235 388585 ;
    LAYER V1 ;
      RECT 2065 392615 2235 392785 ;
    LAYER V1 ;
      RECT 2065 394295 2235 394465 ;
    LAYER V1 ;
      RECT 2065 398495 2235 398665 ;
    LAYER V1 ;
      RECT 2065 400175 2235 400345 ;
    LAYER V1 ;
      RECT 2065 404375 2235 404545 ;
    LAYER V1 ;
      RECT 2065 406055 2235 406225 ;
    LAYER V1 ;
      RECT 2065 410255 2235 410425 ;
    LAYER V1 ;
      RECT 2065 411935 2235 412105 ;
    LAYER V1 ;
      RECT 2065 416135 2235 416305 ;
    LAYER V1 ;
      RECT 2065 417815 2235 417985 ;
    LAYER V1 ;
      RECT 2065 422015 2235 422185 ;
    LAYER V1 ;
      RECT 2065 423695 2235 423865 ;
    LAYER V1 ;
      RECT 2065 427895 2235 428065 ;
    LAYER V1 ;
      RECT 2065 429575 2235 429745 ;
    LAYER V1 ;
      RECT 2065 433775 2235 433945 ;
    LAYER V1 ;
      RECT 2065 435875 2235 436045 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 775 141875 945 142045 ;
    LAYER V1 ;
      RECT 775 147755 945 147925 ;
    LAYER V1 ;
      RECT 775 153635 945 153805 ;
    LAYER V1 ;
      RECT 775 159515 945 159685 ;
    LAYER V1 ;
      RECT 775 165395 945 165565 ;
    LAYER V1 ;
      RECT 775 171275 945 171445 ;
    LAYER V1 ;
      RECT 775 177155 945 177325 ;
    LAYER V1 ;
      RECT 775 183035 945 183205 ;
    LAYER V1 ;
      RECT 775 188915 945 189085 ;
    LAYER V1 ;
      RECT 775 194795 945 194965 ;
    LAYER V1 ;
      RECT 775 200675 945 200845 ;
    LAYER V1 ;
      RECT 775 206555 945 206725 ;
    LAYER V1 ;
      RECT 775 212435 945 212605 ;
    LAYER V1 ;
      RECT 775 218315 945 218485 ;
    LAYER V1 ;
      RECT 775 224195 945 224365 ;
    LAYER V1 ;
      RECT 775 230075 945 230245 ;
    LAYER V1 ;
      RECT 775 235955 945 236125 ;
    LAYER V1 ;
      RECT 775 241835 945 242005 ;
    LAYER V1 ;
      RECT 775 247715 945 247885 ;
    LAYER V1 ;
      RECT 775 253595 945 253765 ;
    LAYER V1 ;
      RECT 775 259475 945 259645 ;
    LAYER V1 ;
      RECT 775 265355 945 265525 ;
    LAYER V1 ;
      RECT 775 271235 945 271405 ;
    LAYER V1 ;
      RECT 775 277115 945 277285 ;
    LAYER V1 ;
      RECT 775 282995 945 283165 ;
    LAYER V1 ;
      RECT 775 288875 945 289045 ;
    LAYER V1 ;
      RECT 775 294755 945 294925 ;
    LAYER V1 ;
      RECT 775 300635 945 300805 ;
    LAYER V1 ;
      RECT 775 306515 945 306685 ;
    LAYER V1 ;
      RECT 775 312395 945 312565 ;
    LAYER V1 ;
      RECT 775 318275 945 318445 ;
    LAYER V1 ;
      RECT 775 324155 945 324325 ;
    LAYER V1 ;
      RECT 775 330035 945 330205 ;
    LAYER V1 ;
      RECT 775 335915 945 336085 ;
    LAYER V1 ;
      RECT 775 341795 945 341965 ;
    LAYER V1 ;
      RECT 775 347675 945 347845 ;
    LAYER V1 ;
      RECT 775 353555 945 353725 ;
    LAYER V1 ;
      RECT 775 359435 945 359605 ;
    LAYER V1 ;
      RECT 775 365315 945 365485 ;
    LAYER V1 ;
      RECT 775 371195 945 371365 ;
    LAYER V1 ;
      RECT 775 377075 945 377245 ;
    LAYER V1 ;
      RECT 775 382955 945 383125 ;
    LAYER V1 ;
      RECT 775 388835 945 389005 ;
    LAYER V1 ;
      RECT 775 394715 945 394885 ;
    LAYER V1 ;
      RECT 775 400595 945 400765 ;
    LAYER V1 ;
      RECT 775 406475 945 406645 ;
    LAYER V1 ;
      RECT 775 412355 945 412525 ;
    LAYER V1 ;
      RECT 775 418235 945 418405 ;
    LAYER V1 ;
      RECT 775 424115 945 424285 ;
    LAYER V1 ;
      RECT 775 429995 945 430165 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 1635 141875 1805 142045 ;
    LAYER V1 ;
      RECT 1635 147755 1805 147925 ;
    LAYER V1 ;
      RECT 1635 153635 1805 153805 ;
    LAYER V1 ;
      RECT 1635 159515 1805 159685 ;
    LAYER V1 ;
      RECT 1635 165395 1805 165565 ;
    LAYER V1 ;
      RECT 1635 171275 1805 171445 ;
    LAYER V1 ;
      RECT 1635 177155 1805 177325 ;
    LAYER V1 ;
      RECT 1635 183035 1805 183205 ;
    LAYER V1 ;
      RECT 1635 188915 1805 189085 ;
    LAYER V1 ;
      RECT 1635 194795 1805 194965 ;
    LAYER V1 ;
      RECT 1635 200675 1805 200845 ;
    LAYER V1 ;
      RECT 1635 206555 1805 206725 ;
    LAYER V1 ;
      RECT 1635 212435 1805 212605 ;
    LAYER V1 ;
      RECT 1635 218315 1805 218485 ;
    LAYER V1 ;
      RECT 1635 224195 1805 224365 ;
    LAYER V1 ;
      RECT 1635 230075 1805 230245 ;
    LAYER V1 ;
      RECT 1635 235955 1805 236125 ;
    LAYER V1 ;
      RECT 1635 241835 1805 242005 ;
    LAYER V1 ;
      RECT 1635 247715 1805 247885 ;
    LAYER V1 ;
      RECT 1635 253595 1805 253765 ;
    LAYER V1 ;
      RECT 1635 259475 1805 259645 ;
    LAYER V1 ;
      RECT 1635 265355 1805 265525 ;
    LAYER V1 ;
      RECT 1635 271235 1805 271405 ;
    LAYER V1 ;
      RECT 1635 277115 1805 277285 ;
    LAYER V1 ;
      RECT 1635 282995 1805 283165 ;
    LAYER V1 ;
      RECT 1635 288875 1805 289045 ;
    LAYER V1 ;
      RECT 1635 294755 1805 294925 ;
    LAYER V1 ;
      RECT 1635 300635 1805 300805 ;
    LAYER V1 ;
      RECT 1635 306515 1805 306685 ;
    LAYER V1 ;
      RECT 1635 312395 1805 312565 ;
    LAYER V1 ;
      RECT 1635 318275 1805 318445 ;
    LAYER V1 ;
      RECT 1635 324155 1805 324325 ;
    LAYER V1 ;
      RECT 1635 330035 1805 330205 ;
    LAYER V1 ;
      RECT 1635 335915 1805 336085 ;
    LAYER V1 ;
      RECT 1635 341795 1805 341965 ;
    LAYER V1 ;
      RECT 1635 347675 1805 347845 ;
    LAYER V1 ;
      RECT 1635 353555 1805 353725 ;
    LAYER V1 ;
      RECT 1635 359435 1805 359605 ;
    LAYER V1 ;
      RECT 1635 365315 1805 365485 ;
    LAYER V1 ;
      RECT 1635 371195 1805 371365 ;
    LAYER V1 ;
      RECT 1635 377075 1805 377245 ;
    LAYER V1 ;
      RECT 1635 382955 1805 383125 ;
    LAYER V1 ;
      RECT 1635 388835 1805 389005 ;
    LAYER V1 ;
      RECT 1635 394715 1805 394885 ;
    LAYER V1 ;
      RECT 1635 400595 1805 400765 ;
    LAYER V1 ;
      RECT 1635 406475 1805 406645 ;
    LAYER V1 ;
      RECT 1635 412355 1805 412525 ;
    LAYER V1 ;
      RECT 1635 418235 1805 418405 ;
    LAYER V1 ;
      RECT 1635 424115 1805 424285 ;
    LAYER V1 ;
      RECT 1635 429995 1805 430165 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V1 ;
      RECT 2495 53675 2665 53845 ;
    LAYER V1 ;
      RECT 2495 59555 2665 59725 ;
    LAYER V1 ;
      RECT 2495 65435 2665 65605 ;
    LAYER V1 ;
      RECT 2495 71315 2665 71485 ;
    LAYER V1 ;
      RECT 2495 77195 2665 77365 ;
    LAYER V1 ;
      RECT 2495 83075 2665 83245 ;
    LAYER V1 ;
      RECT 2495 88955 2665 89125 ;
    LAYER V1 ;
      RECT 2495 94835 2665 95005 ;
    LAYER V1 ;
      RECT 2495 100715 2665 100885 ;
    LAYER V1 ;
      RECT 2495 106595 2665 106765 ;
    LAYER V1 ;
      RECT 2495 112475 2665 112645 ;
    LAYER V1 ;
      RECT 2495 118355 2665 118525 ;
    LAYER V1 ;
      RECT 2495 124235 2665 124405 ;
    LAYER V1 ;
      RECT 2495 130115 2665 130285 ;
    LAYER V1 ;
      RECT 2495 135995 2665 136165 ;
    LAYER V1 ;
      RECT 2495 141875 2665 142045 ;
    LAYER V1 ;
      RECT 2495 147755 2665 147925 ;
    LAYER V1 ;
      RECT 2495 153635 2665 153805 ;
    LAYER V1 ;
      RECT 2495 159515 2665 159685 ;
    LAYER V1 ;
      RECT 2495 165395 2665 165565 ;
    LAYER V1 ;
      RECT 2495 171275 2665 171445 ;
    LAYER V1 ;
      RECT 2495 177155 2665 177325 ;
    LAYER V1 ;
      RECT 2495 183035 2665 183205 ;
    LAYER V1 ;
      RECT 2495 188915 2665 189085 ;
    LAYER V1 ;
      RECT 2495 194795 2665 194965 ;
    LAYER V1 ;
      RECT 2495 200675 2665 200845 ;
    LAYER V1 ;
      RECT 2495 206555 2665 206725 ;
    LAYER V1 ;
      RECT 2495 212435 2665 212605 ;
    LAYER V1 ;
      RECT 2495 218315 2665 218485 ;
    LAYER V1 ;
      RECT 2495 224195 2665 224365 ;
    LAYER V1 ;
      RECT 2495 230075 2665 230245 ;
    LAYER V1 ;
      RECT 2495 235955 2665 236125 ;
    LAYER V1 ;
      RECT 2495 241835 2665 242005 ;
    LAYER V1 ;
      RECT 2495 247715 2665 247885 ;
    LAYER V1 ;
      RECT 2495 253595 2665 253765 ;
    LAYER V1 ;
      RECT 2495 259475 2665 259645 ;
    LAYER V1 ;
      RECT 2495 265355 2665 265525 ;
    LAYER V1 ;
      RECT 2495 271235 2665 271405 ;
    LAYER V1 ;
      RECT 2495 277115 2665 277285 ;
    LAYER V1 ;
      RECT 2495 282995 2665 283165 ;
    LAYER V1 ;
      RECT 2495 288875 2665 289045 ;
    LAYER V1 ;
      RECT 2495 294755 2665 294925 ;
    LAYER V1 ;
      RECT 2495 300635 2665 300805 ;
    LAYER V1 ;
      RECT 2495 306515 2665 306685 ;
    LAYER V1 ;
      RECT 2495 312395 2665 312565 ;
    LAYER V1 ;
      RECT 2495 318275 2665 318445 ;
    LAYER V1 ;
      RECT 2495 324155 2665 324325 ;
    LAYER V1 ;
      RECT 2495 330035 2665 330205 ;
    LAYER V1 ;
      RECT 2495 335915 2665 336085 ;
    LAYER V1 ;
      RECT 2495 341795 2665 341965 ;
    LAYER V1 ;
      RECT 2495 347675 2665 347845 ;
    LAYER V1 ;
      RECT 2495 353555 2665 353725 ;
    LAYER V1 ;
      RECT 2495 359435 2665 359605 ;
    LAYER V1 ;
      RECT 2495 365315 2665 365485 ;
    LAYER V1 ;
      RECT 2495 371195 2665 371365 ;
    LAYER V1 ;
      RECT 2495 377075 2665 377245 ;
    LAYER V1 ;
      RECT 2495 382955 2665 383125 ;
    LAYER V1 ;
      RECT 2495 388835 2665 389005 ;
    LAYER V1 ;
      RECT 2495 394715 2665 394885 ;
    LAYER V1 ;
      RECT 2495 400595 2665 400765 ;
    LAYER V1 ;
      RECT 2495 406475 2665 406645 ;
    LAYER V1 ;
      RECT 2495 412355 2665 412525 ;
    LAYER V1 ;
      RECT 2495 418235 2665 418405 ;
    LAYER V1 ;
      RECT 2495 424115 2665 424285 ;
    LAYER V1 ;
      RECT 2495 429995 2665 430165 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 6225 1365 6375 ;
    LAYER V2 ;
      RECT 1215 12105 1365 12255 ;
    LAYER V2 ;
      RECT 1215 17985 1365 18135 ;
    LAYER V2 ;
      RECT 1215 23865 1365 24015 ;
    LAYER V2 ;
      RECT 1215 29745 1365 29895 ;
    LAYER V2 ;
      RECT 1215 35625 1365 35775 ;
    LAYER V2 ;
      RECT 1215 41505 1365 41655 ;
    LAYER V2 ;
      RECT 1215 47385 1365 47535 ;
    LAYER V2 ;
      RECT 1215 53265 1365 53415 ;
    LAYER V2 ;
      RECT 1215 59145 1365 59295 ;
    LAYER V2 ;
      RECT 1215 65025 1365 65175 ;
    LAYER V2 ;
      RECT 1215 70905 1365 71055 ;
    LAYER V2 ;
      RECT 1215 76785 1365 76935 ;
    LAYER V2 ;
      RECT 1215 82665 1365 82815 ;
    LAYER V2 ;
      RECT 1215 88545 1365 88695 ;
    LAYER V2 ;
      RECT 1215 94425 1365 94575 ;
    LAYER V2 ;
      RECT 1215 100305 1365 100455 ;
    LAYER V2 ;
      RECT 1215 106185 1365 106335 ;
    LAYER V2 ;
      RECT 1215 112065 1365 112215 ;
    LAYER V2 ;
      RECT 1215 117945 1365 118095 ;
    LAYER V2 ;
      RECT 1215 123825 1365 123975 ;
    LAYER V2 ;
      RECT 1215 129705 1365 129855 ;
    LAYER V2 ;
      RECT 1215 135585 1365 135735 ;
    LAYER V2 ;
      RECT 1215 141465 1365 141615 ;
    LAYER V2 ;
      RECT 1215 147345 1365 147495 ;
    LAYER V2 ;
      RECT 1215 153225 1365 153375 ;
    LAYER V2 ;
      RECT 1215 159105 1365 159255 ;
    LAYER V2 ;
      RECT 1215 164985 1365 165135 ;
    LAYER V2 ;
      RECT 1215 170865 1365 171015 ;
    LAYER V2 ;
      RECT 1215 176745 1365 176895 ;
    LAYER V2 ;
      RECT 1215 182625 1365 182775 ;
    LAYER V2 ;
      RECT 1215 188505 1365 188655 ;
    LAYER V2 ;
      RECT 1215 194385 1365 194535 ;
    LAYER V2 ;
      RECT 1215 200265 1365 200415 ;
    LAYER V2 ;
      RECT 1215 206145 1365 206295 ;
    LAYER V2 ;
      RECT 1215 212025 1365 212175 ;
    LAYER V2 ;
      RECT 1215 217905 1365 218055 ;
    LAYER V2 ;
      RECT 1215 223785 1365 223935 ;
    LAYER V2 ;
      RECT 1215 229665 1365 229815 ;
    LAYER V2 ;
      RECT 1215 235545 1365 235695 ;
    LAYER V2 ;
      RECT 1215 241425 1365 241575 ;
    LAYER V2 ;
      RECT 1215 247305 1365 247455 ;
    LAYER V2 ;
      RECT 1215 253185 1365 253335 ;
    LAYER V2 ;
      RECT 1215 259065 1365 259215 ;
    LAYER V2 ;
      RECT 1215 264945 1365 265095 ;
    LAYER V2 ;
      RECT 1215 270825 1365 270975 ;
    LAYER V2 ;
      RECT 1215 276705 1365 276855 ;
    LAYER V2 ;
      RECT 1215 282585 1365 282735 ;
    LAYER V2 ;
      RECT 1215 288465 1365 288615 ;
    LAYER V2 ;
      RECT 1215 294345 1365 294495 ;
    LAYER V2 ;
      RECT 1215 300225 1365 300375 ;
    LAYER V2 ;
      RECT 1215 306105 1365 306255 ;
    LAYER V2 ;
      RECT 1215 311985 1365 312135 ;
    LAYER V2 ;
      RECT 1215 317865 1365 318015 ;
    LAYER V2 ;
      RECT 1215 323745 1365 323895 ;
    LAYER V2 ;
      RECT 1215 329625 1365 329775 ;
    LAYER V2 ;
      RECT 1215 335505 1365 335655 ;
    LAYER V2 ;
      RECT 1215 341385 1365 341535 ;
    LAYER V2 ;
      RECT 1215 347265 1365 347415 ;
    LAYER V2 ;
      RECT 1215 353145 1365 353295 ;
    LAYER V2 ;
      RECT 1215 359025 1365 359175 ;
    LAYER V2 ;
      RECT 1215 364905 1365 365055 ;
    LAYER V2 ;
      RECT 1215 370785 1365 370935 ;
    LAYER V2 ;
      RECT 1215 376665 1365 376815 ;
    LAYER V2 ;
      RECT 1215 382545 1365 382695 ;
    LAYER V2 ;
      RECT 1215 388425 1365 388575 ;
    LAYER V2 ;
      RECT 1215 394305 1365 394455 ;
    LAYER V2 ;
      RECT 1215 400185 1365 400335 ;
    LAYER V2 ;
      RECT 1215 406065 1365 406215 ;
    LAYER V2 ;
      RECT 1215 411945 1365 412095 ;
    LAYER V2 ;
      RECT 1215 417825 1365 417975 ;
    LAYER V2 ;
      RECT 1215 423705 1365 423855 ;
    LAYER V2 ;
      RECT 1215 429585 1365 429735 ;
    LAYER V2 ;
      RECT 1645 4545 1795 4695 ;
    LAYER V2 ;
      RECT 1645 10425 1795 10575 ;
    LAYER V2 ;
      RECT 1645 16305 1795 16455 ;
    LAYER V2 ;
      RECT 1645 22185 1795 22335 ;
    LAYER V2 ;
      RECT 1645 28065 1795 28215 ;
    LAYER V2 ;
      RECT 1645 33945 1795 34095 ;
    LAYER V2 ;
      RECT 1645 39825 1795 39975 ;
    LAYER V2 ;
      RECT 1645 45705 1795 45855 ;
    LAYER V2 ;
      RECT 1645 51585 1795 51735 ;
    LAYER V2 ;
      RECT 1645 57465 1795 57615 ;
    LAYER V2 ;
      RECT 1645 63345 1795 63495 ;
    LAYER V2 ;
      RECT 1645 69225 1795 69375 ;
    LAYER V2 ;
      RECT 1645 75105 1795 75255 ;
    LAYER V2 ;
      RECT 1645 80985 1795 81135 ;
    LAYER V2 ;
      RECT 1645 86865 1795 87015 ;
    LAYER V2 ;
      RECT 1645 92745 1795 92895 ;
    LAYER V2 ;
      RECT 1645 98625 1795 98775 ;
    LAYER V2 ;
      RECT 1645 104505 1795 104655 ;
    LAYER V2 ;
      RECT 1645 110385 1795 110535 ;
    LAYER V2 ;
      RECT 1645 116265 1795 116415 ;
    LAYER V2 ;
      RECT 1645 122145 1795 122295 ;
    LAYER V2 ;
      RECT 1645 128025 1795 128175 ;
    LAYER V2 ;
      RECT 1645 133905 1795 134055 ;
    LAYER V2 ;
      RECT 1645 139785 1795 139935 ;
    LAYER V2 ;
      RECT 1645 145665 1795 145815 ;
    LAYER V2 ;
      RECT 1645 151545 1795 151695 ;
    LAYER V2 ;
      RECT 1645 157425 1795 157575 ;
    LAYER V2 ;
      RECT 1645 163305 1795 163455 ;
    LAYER V2 ;
      RECT 1645 169185 1795 169335 ;
    LAYER V2 ;
      RECT 1645 175065 1795 175215 ;
    LAYER V2 ;
      RECT 1645 180945 1795 181095 ;
    LAYER V2 ;
      RECT 1645 186825 1795 186975 ;
    LAYER V2 ;
      RECT 1645 192705 1795 192855 ;
    LAYER V2 ;
      RECT 1645 198585 1795 198735 ;
    LAYER V2 ;
      RECT 1645 204465 1795 204615 ;
    LAYER V2 ;
      RECT 1645 210345 1795 210495 ;
    LAYER V2 ;
      RECT 1645 216225 1795 216375 ;
    LAYER V2 ;
      RECT 1645 222105 1795 222255 ;
    LAYER V2 ;
      RECT 1645 227985 1795 228135 ;
    LAYER V2 ;
      RECT 1645 233865 1795 234015 ;
    LAYER V2 ;
      RECT 1645 239745 1795 239895 ;
    LAYER V2 ;
      RECT 1645 245625 1795 245775 ;
    LAYER V2 ;
      RECT 1645 251505 1795 251655 ;
    LAYER V2 ;
      RECT 1645 257385 1795 257535 ;
    LAYER V2 ;
      RECT 1645 263265 1795 263415 ;
    LAYER V2 ;
      RECT 1645 269145 1795 269295 ;
    LAYER V2 ;
      RECT 1645 275025 1795 275175 ;
    LAYER V2 ;
      RECT 1645 280905 1795 281055 ;
    LAYER V2 ;
      RECT 1645 286785 1795 286935 ;
    LAYER V2 ;
      RECT 1645 292665 1795 292815 ;
    LAYER V2 ;
      RECT 1645 298545 1795 298695 ;
    LAYER V2 ;
      RECT 1645 304425 1795 304575 ;
    LAYER V2 ;
      RECT 1645 310305 1795 310455 ;
    LAYER V2 ;
      RECT 1645 316185 1795 316335 ;
    LAYER V2 ;
      RECT 1645 322065 1795 322215 ;
    LAYER V2 ;
      RECT 1645 327945 1795 328095 ;
    LAYER V2 ;
      RECT 1645 333825 1795 333975 ;
    LAYER V2 ;
      RECT 1645 339705 1795 339855 ;
    LAYER V2 ;
      RECT 1645 345585 1795 345735 ;
    LAYER V2 ;
      RECT 1645 351465 1795 351615 ;
    LAYER V2 ;
      RECT 1645 357345 1795 357495 ;
    LAYER V2 ;
      RECT 1645 363225 1795 363375 ;
    LAYER V2 ;
      RECT 1645 369105 1795 369255 ;
    LAYER V2 ;
      RECT 1645 374985 1795 375135 ;
    LAYER V2 ;
      RECT 1645 380865 1795 381015 ;
    LAYER V2 ;
      RECT 1645 386745 1795 386895 ;
    LAYER V2 ;
      RECT 1645 392625 1795 392775 ;
    LAYER V2 ;
      RECT 1645 398505 1795 398655 ;
    LAYER V2 ;
      RECT 1645 404385 1795 404535 ;
    LAYER V2 ;
      RECT 1645 410265 1795 410415 ;
    LAYER V2 ;
      RECT 1645 416145 1795 416295 ;
    LAYER V2 ;
      RECT 1645 422025 1795 422175 ;
    LAYER V2 ;
      RECT 1645 427905 1795 428055 ;
    LAYER V2 ;
      RECT 1645 433785 1795 433935 ;
    LAYER V2 ;
      RECT 2075 765 2225 915 ;
    LAYER V2 ;
      RECT 2075 6645 2225 6795 ;
    LAYER V2 ;
      RECT 2075 12525 2225 12675 ;
    LAYER V2 ;
      RECT 2075 18405 2225 18555 ;
    LAYER V2 ;
      RECT 2075 24285 2225 24435 ;
    LAYER V2 ;
      RECT 2075 30165 2225 30315 ;
    LAYER V2 ;
      RECT 2075 36045 2225 36195 ;
    LAYER V2 ;
      RECT 2075 41925 2225 42075 ;
    LAYER V2 ;
      RECT 2075 47805 2225 47955 ;
    LAYER V2 ;
      RECT 2075 53685 2225 53835 ;
    LAYER V2 ;
      RECT 2075 59565 2225 59715 ;
    LAYER V2 ;
      RECT 2075 65445 2225 65595 ;
    LAYER V2 ;
      RECT 2075 71325 2225 71475 ;
    LAYER V2 ;
      RECT 2075 77205 2225 77355 ;
    LAYER V2 ;
      RECT 2075 83085 2225 83235 ;
    LAYER V2 ;
      RECT 2075 88965 2225 89115 ;
    LAYER V2 ;
      RECT 2075 94845 2225 94995 ;
    LAYER V2 ;
      RECT 2075 100725 2225 100875 ;
    LAYER V2 ;
      RECT 2075 106605 2225 106755 ;
    LAYER V2 ;
      RECT 2075 112485 2225 112635 ;
    LAYER V2 ;
      RECT 2075 118365 2225 118515 ;
    LAYER V2 ;
      RECT 2075 124245 2225 124395 ;
    LAYER V2 ;
      RECT 2075 130125 2225 130275 ;
    LAYER V2 ;
      RECT 2075 136005 2225 136155 ;
    LAYER V2 ;
      RECT 2075 141885 2225 142035 ;
    LAYER V2 ;
      RECT 2075 147765 2225 147915 ;
    LAYER V2 ;
      RECT 2075 153645 2225 153795 ;
    LAYER V2 ;
      RECT 2075 159525 2225 159675 ;
    LAYER V2 ;
      RECT 2075 165405 2225 165555 ;
    LAYER V2 ;
      RECT 2075 171285 2225 171435 ;
    LAYER V2 ;
      RECT 2075 177165 2225 177315 ;
    LAYER V2 ;
      RECT 2075 183045 2225 183195 ;
    LAYER V2 ;
      RECT 2075 188925 2225 189075 ;
    LAYER V2 ;
      RECT 2075 194805 2225 194955 ;
    LAYER V2 ;
      RECT 2075 200685 2225 200835 ;
    LAYER V2 ;
      RECT 2075 206565 2225 206715 ;
    LAYER V2 ;
      RECT 2075 212445 2225 212595 ;
    LAYER V2 ;
      RECT 2075 218325 2225 218475 ;
    LAYER V2 ;
      RECT 2075 224205 2225 224355 ;
    LAYER V2 ;
      RECT 2075 230085 2225 230235 ;
    LAYER V2 ;
      RECT 2075 235965 2225 236115 ;
    LAYER V2 ;
      RECT 2075 241845 2225 241995 ;
    LAYER V2 ;
      RECT 2075 247725 2225 247875 ;
    LAYER V2 ;
      RECT 2075 253605 2225 253755 ;
    LAYER V2 ;
      RECT 2075 259485 2225 259635 ;
    LAYER V2 ;
      RECT 2075 265365 2225 265515 ;
    LAYER V2 ;
      RECT 2075 271245 2225 271395 ;
    LAYER V2 ;
      RECT 2075 277125 2225 277275 ;
    LAYER V2 ;
      RECT 2075 283005 2225 283155 ;
    LAYER V2 ;
      RECT 2075 288885 2225 289035 ;
    LAYER V2 ;
      RECT 2075 294765 2225 294915 ;
    LAYER V2 ;
      RECT 2075 300645 2225 300795 ;
    LAYER V2 ;
      RECT 2075 306525 2225 306675 ;
    LAYER V2 ;
      RECT 2075 312405 2225 312555 ;
    LAYER V2 ;
      RECT 2075 318285 2225 318435 ;
    LAYER V2 ;
      RECT 2075 324165 2225 324315 ;
    LAYER V2 ;
      RECT 2075 330045 2225 330195 ;
    LAYER V2 ;
      RECT 2075 335925 2225 336075 ;
    LAYER V2 ;
      RECT 2075 341805 2225 341955 ;
    LAYER V2 ;
      RECT 2075 347685 2225 347835 ;
    LAYER V2 ;
      RECT 2075 353565 2225 353715 ;
    LAYER V2 ;
      RECT 2075 359445 2225 359595 ;
    LAYER V2 ;
      RECT 2075 365325 2225 365475 ;
    LAYER V2 ;
      RECT 2075 371205 2225 371355 ;
    LAYER V2 ;
      RECT 2075 377085 2225 377235 ;
    LAYER V2 ;
      RECT 2075 382965 2225 383115 ;
    LAYER V2 ;
      RECT 2075 388845 2225 388995 ;
    LAYER V2 ;
      RECT 2075 394725 2225 394875 ;
    LAYER V2 ;
      RECT 2075 400605 2225 400755 ;
    LAYER V2 ;
      RECT 2075 406485 2225 406635 ;
    LAYER V2 ;
      RECT 2075 412365 2225 412515 ;
    LAYER V2 ;
      RECT 2075 418245 2225 418395 ;
    LAYER V2 ;
      RECT 2075 424125 2225 424275 ;
    LAYER V2 ;
      RECT 2075 430005 2225 430155 ;
    LAYER V2 ;
      RECT 2075 435885 2225 436035 ;
  END
END NMOS_S_12565100_X2_Y74
