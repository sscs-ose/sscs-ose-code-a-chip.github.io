# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  3.720000 BY  4.110000 ;
  PIN DRAIN
    ANTENNADIFFAREA  3.360000 ;
    PORT
      LAYER met3 ;
        RECT 0.585000 2.365000 0.915000 2.805000 ;
        RECT 0.585000 2.805000 3.495000 3.135000 ;
        RECT 1.445000 2.365000 1.775000 2.805000 ;
        RECT 2.305000 2.365000 2.635000 2.805000 ;
        RECT 3.165000 2.365000 3.495000 2.805000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.600000 ;
    PORT
      LAYER met1 ;
        RECT 0.635000 3.355000 3.445000 3.645000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.200000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 3.875000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  3.105000 ;
        RECT 1.065000 -0.145000 1.295000  3.105000 ;
        RECT 1.925000 -0.145000 2.155000  3.105000 ;
        RECT 2.785000 -0.145000 3.015000  3.105000 ;
        RECT 3.645000 -0.145000 3.875000  3.105000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.395000 3.195000 0.445000 3.290000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.255000 0.405000 3.105000 ;
      RECT 0.665000 0.255000 0.835000 3.105000 ;
      RECT 0.685000 3.335000 3.395000 3.665000 ;
      RECT 1.095000 0.255000 1.265000 3.105000 ;
      RECT 1.525000 0.255000 1.695000 3.105000 ;
      RECT 1.955000 0.255000 2.125000 3.105000 ;
      RECT 2.385000 0.255000 2.555000 3.105000 ;
      RECT 2.815000 0.255000 2.985000 3.105000 ;
      RECT 3.245000 0.255000 3.415000 3.105000 ;
      RECT 3.675000 0.255000 3.845000 3.105000 ;
    LAYER mcon ;
      RECT 0.235000 0.335000 0.405000 0.505000 ;
      RECT 0.235000 0.695000 0.405000 0.865000 ;
      RECT 0.235000 1.055000 0.405000 1.225000 ;
      RECT 0.235000 1.415000 0.405000 1.585000 ;
      RECT 0.235000 1.775000 0.405000 1.945000 ;
      RECT 0.235000 2.135000 0.405000 2.305000 ;
      RECT 0.235000 2.495000 0.405000 2.665000 ;
      RECT 0.235000 2.855000 0.405000 3.025000 ;
      RECT 0.665000 0.335000 0.835000 0.505000 ;
      RECT 0.665000 0.695000 0.835000 0.865000 ;
      RECT 0.665000 1.055000 0.835000 1.225000 ;
      RECT 0.665000 1.415000 0.835000 1.585000 ;
      RECT 0.665000 1.775000 0.835000 1.945000 ;
      RECT 0.665000 2.135000 0.835000 2.305000 ;
      RECT 0.665000 2.495000 0.835000 2.665000 ;
      RECT 0.665000 2.855000 0.835000 3.025000 ;
      RECT 0.695000 3.415000 0.865000 3.585000 ;
      RECT 1.055000 3.415000 1.225000 3.585000 ;
      RECT 1.095000 0.335000 1.265000 0.505000 ;
      RECT 1.095000 0.695000 1.265000 0.865000 ;
      RECT 1.095000 1.055000 1.265000 1.225000 ;
      RECT 1.095000 1.415000 1.265000 1.585000 ;
      RECT 1.095000 1.775000 1.265000 1.945000 ;
      RECT 1.095000 2.135000 1.265000 2.305000 ;
      RECT 1.095000 2.495000 1.265000 2.665000 ;
      RECT 1.095000 2.855000 1.265000 3.025000 ;
      RECT 1.415000 3.415000 1.585000 3.585000 ;
      RECT 1.525000 0.335000 1.695000 0.505000 ;
      RECT 1.525000 0.695000 1.695000 0.865000 ;
      RECT 1.525000 1.055000 1.695000 1.225000 ;
      RECT 1.525000 1.415000 1.695000 1.585000 ;
      RECT 1.525000 1.775000 1.695000 1.945000 ;
      RECT 1.525000 2.135000 1.695000 2.305000 ;
      RECT 1.525000 2.495000 1.695000 2.665000 ;
      RECT 1.525000 2.855000 1.695000 3.025000 ;
      RECT 1.775000 3.415000 1.945000 3.585000 ;
      RECT 1.955000 0.335000 2.125000 0.505000 ;
      RECT 1.955000 0.695000 2.125000 0.865000 ;
      RECT 1.955000 1.055000 2.125000 1.225000 ;
      RECT 1.955000 1.415000 2.125000 1.585000 ;
      RECT 1.955000 1.775000 2.125000 1.945000 ;
      RECT 1.955000 2.135000 2.125000 2.305000 ;
      RECT 1.955000 2.495000 2.125000 2.665000 ;
      RECT 1.955000 2.855000 2.125000 3.025000 ;
      RECT 2.135000 3.415000 2.305000 3.585000 ;
      RECT 2.385000 0.335000 2.555000 0.505000 ;
      RECT 2.385000 0.695000 2.555000 0.865000 ;
      RECT 2.385000 1.055000 2.555000 1.225000 ;
      RECT 2.385000 1.415000 2.555000 1.585000 ;
      RECT 2.385000 1.775000 2.555000 1.945000 ;
      RECT 2.385000 2.135000 2.555000 2.305000 ;
      RECT 2.385000 2.495000 2.555000 2.665000 ;
      RECT 2.385000 2.855000 2.555000 3.025000 ;
      RECT 2.495000 3.415000 2.665000 3.585000 ;
      RECT 2.815000 0.335000 2.985000 0.505000 ;
      RECT 2.815000 0.695000 2.985000 0.865000 ;
      RECT 2.815000 1.055000 2.985000 1.225000 ;
      RECT 2.815000 1.415000 2.985000 1.585000 ;
      RECT 2.815000 1.775000 2.985000 1.945000 ;
      RECT 2.815000 2.135000 2.985000 2.305000 ;
      RECT 2.815000 2.495000 2.985000 2.665000 ;
      RECT 2.815000 2.855000 2.985000 3.025000 ;
      RECT 2.855000 3.415000 3.025000 3.585000 ;
      RECT 3.215000 3.415000 3.385000 3.585000 ;
      RECT 3.245000 0.335000 3.415000 0.505000 ;
      RECT 3.245000 0.695000 3.415000 0.865000 ;
      RECT 3.245000 1.055000 3.415000 1.225000 ;
      RECT 3.245000 1.415000 3.415000 1.585000 ;
      RECT 3.245000 1.775000 3.415000 1.945000 ;
      RECT 3.245000 2.135000 3.415000 2.305000 ;
      RECT 3.245000 2.495000 3.415000 2.665000 ;
      RECT 3.245000 2.855000 3.415000 3.025000 ;
      RECT 3.675000 0.335000 3.845000 0.505000 ;
      RECT 3.675000 0.695000 3.845000 0.865000 ;
      RECT 3.675000 1.055000 3.845000 1.225000 ;
      RECT 3.675000 1.415000 3.845000 1.585000 ;
      RECT 3.675000 1.775000 3.845000 1.945000 ;
      RECT 3.675000 2.135000 3.845000 2.305000 ;
      RECT 3.675000 2.495000 3.845000 2.665000 ;
      RECT 3.675000 2.855000 3.845000 3.025000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 3.105000 ;
      RECT 1.480000 0.255000 1.740000 3.105000 ;
      RECT 2.340000 0.255000 2.600000 3.105000 ;
      RECT 3.200000 0.255000 3.460000 3.105000 ;
    LAYER met2 ;
      RECT 0.585000 2.365000 0.915000 3.135000 ;
      RECT 1.445000 2.365000 1.775000 3.135000 ;
      RECT 2.305000 2.365000 2.635000 3.135000 ;
      RECT 3.165000 2.365000 3.495000 3.135000 ;
    LAYER via ;
      RECT 0.620000 2.460000 0.880000 2.720000 ;
      RECT 0.620000 2.780000 0.880000 3.040000 ;
      RECT 1.480000 2.460000 1.740000 2.720000 ;
      RECT 1.480000 2.780000 1.740000 3.040000 ;
      RECT 2.340000 2.460000 2.600000 2.720000 ;
      RECT 2.340000 2.780000 2.600000 3.040000 ;
      RECT 3.200000 2.460000 3.460000 2.720000 ;
      RECT 3.200000 2.780000 3.460000 3.040000 ;
    LAYER via2 ;
      RECT 0.610000 2.410000 0.890000 2.690000 ;
      RECT 0.610000 2.810000 0.890000 3.090000 ;
      RECT 1.470000 2.410000 1.750000 2.690000 ;
      RECT 1.470000 2.810000 1.750000 3.090000 ;
      RECT 2.330000 2.410000 2.610000 2.690000 ;
      RECT 2.330000 2.810000 2.610000 3.090000 ;
      RECT 3.190000 2.410000 3.470000 2.690000 ;
      RECT 3.190000 2.810000 3.470000 3.090000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15
END LIBRARY
