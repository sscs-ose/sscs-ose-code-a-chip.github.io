* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+ sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult = 1.042
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult = 1.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult = 0.99758
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult = 1.1193e+0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult = 1.1801e+0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff = -1.21275e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff = 2.252e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff = -1.21275e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff = 2.252e-8
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0 = 0.30329
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0 = 0.01726
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0 = 0.00068868
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0 = 0.024431
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0 = 1583.3
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0 = 1.32e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0 = 1.6741e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1 = 0.28901
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1 = 0.01659
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1 = 0.0023767
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1 = 0.025579
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1 = 1895.9
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1 = 1.438e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1 = 2.8248e-12
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2 = 0.28823
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2 = 0.016801
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2 = 0.00060123
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2 = 0.024939
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2 = 3195.6
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2 = 1.4202e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2 = 1.0136e-11
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3 = 1.3648e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3 = 0.29555
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3 = 0.016145
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3 = 0.00028215
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3 = 0.023983
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3 = 3192.2
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3 = 1.3881e-18
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4 = 1.3703e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4 = 1.7829e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4 = 0.2895
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4 = 0.017958
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4 = 0.00077795
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4 = 0.022447
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4 = 2279.7
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5 = -2.1985e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5 = 6.9289e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5 = 0.33754
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5 = 0.049359
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5 = 0.071277
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5 = 0.043943
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5 = -0.0080434
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5 = 0.013646
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6 = 1.7407e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6 = 1.9509e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6 = 0.29323
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6 = 0.017035
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6 = 0.0011167
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6 = 0.021986
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6 = 4980.3
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7 = 6726.2
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7 = 2.17e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7 = 1.9011e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7 = 0.25951
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7 = 0.017543
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7 = 0.00080633
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7 = 0.021766
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8 = -0.010132
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8 = -0.0032051
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8 = -2.1641e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8 = 6.8574e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8 = 0.31944
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8 = 0.10492
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8 = 0.15983
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8 = 0.00845
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9 = 0.0060854
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9 = 0.0032612
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9 = 0.012301
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9 = 3335.1
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9 = 2.5113e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9 = 1.4426e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9 = 0.27036
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10 = 1.0694e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10 = -198.96
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10 = 7.208e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10 = 0.0071747
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10 = 0.31463
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10 = -0.00052628
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10 = 0.024124
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10 = 0.0
.include "sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"
