magic
tech sky130A
magscale 1 2
timestamp 1666543010
<< nwell >>
rect 2246 8934 2546 8936
rect 2246 8930 6050 8934
rect 522 6680 6050 8930
rect 2472 4686 6050 6680
rect 515 3092 1125 3634
rect 1536 2200 2174 2872
<< nmos >>
rect 613 3785 643 3985
rect 709 3785 739 3985
rect 805 3785 835 3985
rect 901 3785 931 3985
rect 997 3785 1027 3985
<< pmos >>
rect 613 3334 643 3534
rect 709 3334 739 3534
rect 805 3334 835 3534
rect 901 3334 931 3534
rect 997 3334 1027 3534
<< mvnmos >>
rect 646 4320 746 6320
rect 804 4320 904 6320
rect 962 4320 1062 6320
rect 1120 4320 1220 6320
rect 1278 4320 1378 6320
rect 1436 4320 1536 6320
rect 1594 4320 1694 6320
rect 1752 4320 1852 6320
rect 1910 4320 2010 6320
rect 2068 4320 2168 6320
rect 1348 3132 1448 3932
rect 1506 3132 1606 3932
rect 1664 3132 1764 3932
rect 1962 3132 2062 3932
rect 2120 3132 2220 3932
rect 2278 3132 2378 3932
rect 2714 206 2814 4206
rect 2872 206 2972 4206
rect 3030 206 3130 4206
rect 3188 206 3288 4206
rect 3346 206 3446 4206
rect 3504 206 3604 4206
rect 3662 206 3762 4206
rect 3820 206 3920 4206
rect 3978 206 4078 4206
rect 4136 206 4236 4206
rect 4294 206 4394 4206
rect 4452 206 4552 4206
rect 4610 206 4710 4206
rect 4768 206 4868 4206
rect 4926 206 5026 4206
rect 5084 206 5184 4206
rect 5242 206 5342 4206
rect 5400 206 5500 4206
rect 5558 206 5658 4206
rect 5716 206 5816 4206
<< mvpmos >>
rect 646 6746 746 8746
rect 804 6746 904 8746
rect 962 6746 1062 8746
rect 1120 6746 1220 8746
rect 1278 6746 1378 8746
rect 1436 6746 1536 8746
rect 1594 6746 1694 8746
rect 1752 6746 1852 8746
rect 1910 6746 2010 8746
rect 2068 6746 2168 8746
rect 2714 4754 2814 8754
rect 2872 4754 2972 8754
rect 3030 4754 3130 8754
rect 3188 4754 3288 8754
rect 3346 4754 3446 8754
rect 3504 4754 3604 8754
rect 3662 4754 3762 8754
rect 3820 4754 3920 8754
rect 3978 4754 4078 8754
rect 4136 4754 4236 8754
rect 4294 4754 4394 8754
rect 4452 4754 4552 8754
rect 4610 4754 4710 8754
rect 4768 4754 4868 8754
rect 4926 4754 5026 8754
rect 5084 4754 5184 8754
rect 5242 4754 5342 8754
rect 5400 4754 5500 8754
rect 5558 4754 5658 8754
rect 5716 4754 5816 8754
rect 1660 2372 1760 2772
rect 1950 2372 2050 2772
<< ndiff >>
rect 551 3973 613 3985
rect 551 3797 563 3973
rect 597 3797 613 3973
rect 551 3785 613 3797
rect 643 3973 709 3985
rect 643 3797 659 3973
rect 693 3797 709 3973
rect 643 3785 709 3797
rect 739 3973 805 3985
rect 739 3797 755 3973
rect 789 3797 805 3973
rect 739 3785 805 3797
rect 835 3973 901 3985
rect 835 3797 851 3973
rect 885 3797 901 3973
rect 835 3785 901 3797
rect 931 3973 997 3985
rect 931 3797 947 3973
rect 981 3797 997 3973
rect 931 3785 997 3797
rect 1027 3973 1089 3985
rect 1027 3797 1043 3973
rect 1077 3797 1089 3973
rect 1027 3785 1089 3797
<< pdiff >>
rect 551 3522 613 3534
rect 551 3346 563 3522
rect 597 3346 613 3522
rect 551 3334 613 3346
rect 643 3522 709 3534
rect 643 3346 659 3522
rect 693 3346 709 3522
rect 643 3334 709 3346
rect 739 3522 805 3534
rect 739 3346 755 3522
rect 789 3346 805 3522
rect 739 3334 805 3346
rect 835 3522 901 3534
rect 835 3346 851 3522
rect 885 3346 901 3522
rect 835 3334 901 3346
rect 931 3522 997 3534
rect 931 3346 947 3522
rect 981 3346 997 3522
rect 931 3334 997 3346
rect 1027 3522 1089 3534
rect 1027 3346 1043 3522
rect 1077 3346 1089 3522
rect 1027 3334 1089 3346
<< mvndiff >>
rect 588 6308 646 6320
rect 588 4332 600 6308
rect 634 4332 646 6308
rect 588 4320 646 4332
rect 746 6308 804 6320
rect 746 4332 758 6308
rect 792 4332 804 6308
rect 746 4320 804 4332
rect 904 6308 962 6320
rect 904 4332 916 6308
rect 950 4332 962 6308
rect 904 4320 962 4332
rect 1062 6308 1120 6320
rect 1062 4332 1074 6308
rect 1108 4332 1120 6308
rect 1062 4320 1120 4332
rect 1220 6308 1278 6320
rect 1220 4332 1232 6308
rect 1266 4332 1278 6308
rect 1220 4320 1278 4332
rect 1378 6308 1436 6320
rect 1378 4332 1390 6308
rect 1424 4332 1436 6308
rect 1378 4320 1436 4332
rect 1536 6308 1594 6320
rect 1536 4332 1548 6308
rect 1582 4332 1594 6308
rect 1536 4320 1594 4332
rect 1694 6308 1752 6320
rect 1694 4332 1706 6308
rect 1740 4332 1752 6308
rect 1694 4320 1752 4332
rect 1852 6308 1910 6320
rect 1852 4332 1864 6308
rect 1898 4332 1910 6308
rect 1852 4320 1910 4332
rect 2010 6308 2068 6320
rect 2010 4332 2022 6308
rect 2056 4332 2068 6308
rect 2010 4320 2068 4332
rect 2168 6308 2226 6320
rect 2168 4332 2180 6308
rect 2214 4332 2226 6308
rect 2168 4320 2226 4332
rect 2656 4194 2714 4206
rect 1290 3920 1348 3932
rect 1290 3144 1302 3920
rect 1336 3144 1348 3920
rect 1290 3132 1348 3144
rect 1448 3920 1506 3932
rect 1448 3144 1460 3920
rect 1494 3144 1506 3920
rect 1448 3132 1506 3144
rect 1606 3920 1664 3932
rect 1606 3144 1618 3920
rect 1652 3144 1664 3920
rect 1606 3132 1664 3144
rect 1764 3920 1822 3932
rect 1764 3144 1776 3920
rect 1810 3144 1822 3920
rect 1764 3132 1822 3144
rect 1904 3920 1962 3932
rect 1904 3144 1916 3920
rect 1950 3144 1962 3920
rect 1904 3132 1962 3144
rect 2062 3920 2120 3932
rect 2062 3144 2074 3920
rect 2108 3144 2120 3920
rect 2062 3132 2120 3144
rect 2220 3920 2278 3932
rect 2220 3144 2232 3920
rect 2266 3144 2278 3920
rect 2220 3132 2278 3144
rect 2378 3920 2436 3932
rect 2378 3144 2390 3920
rect 2424 3144 2436 3920
rect 2378 3132 2436 3144
rect 2656 218 2668 4194
rect 2702 218 2714 4194
rect 2656 206 2714 218
rect 2814 4194 2872 4206
rect 2814 218 2826 4194
rect 2860 218 2872 4194
rect 2814 206 2872 218
rect 2972 4194 3030 4206
rect 2972 218 2984 4194
rect 3018 218 3030 4194
rect 2972 206 3030 218
rect 3130 4194 3188 4206
rect 3130 218 3142 4194
rect 3176 218 3188 4194
rect 3130 206 3188 218
rect 3288 4194 3346 4206
rect 3288 218 3300 4194
rect 3334 218 3346 4194
rect 3288 206 3346 218
rect 3446 4194 3504 4206
rect 3446 218 3458 4194
rect 3492 218 3504 4194
rect 3446 206 3504 218
rect 3604 4194 3662 4206
rect 3604 218 3616 4194
rect 3650 218 3662 4194
rect 3604 206 3662 218
rect 3762 4194 3820 4206
rect 3762 218 3774 4194
rect 3808 218 3820 4194
rect 3762 206 3820 218
rect 3920 4194 3978 4206
rect 3920 218 3932 4194
rect 3966 218 3978 4194
rect 3920 206 3978 218
rect 4078 4194 4136 4206
rect 4078 218 4090 4194
rect 4124 218 4136 4194
rect 4078 206 4136 218
rect 4236 4194 4294 4206
rect 4236 218 4248 4194
rect 4282 218 4294 4194
rect 4236 206 4294 218
rect 4394 4194 4452 4206
rect 4394 218 4406 4194
rect 4440 218 4452 4194
rect 4394 206 4452 218
rect 4552 4194 4610 4206
rect 4552 218 4564 4194
rect 4598 218 4610 4194
rect 4552 206 4610 218
rect 4710 4194 4768 4206
rect 4710 218 4722 4194
rect 4756 218 4768 4194
rect 4710 206 4768 218
rect 4868 4194 4926 4206
rect 4868 218 4880 4194
rect 4914 218 4926 4194
rect 4868 206 4926 218
rect 5026 4194 5084 4206
rect 5026 218 5038 4194
rect 5072 218 5084 4194
rect 5026 206 5084 218
rect 5184 4194 5242 4206
rect 5184 218 5196 4194
rect 5230 218 5242 4194
rect 5184 206 5242 218
rect 5342 4194 5400 4206
rect 5342 218 5354 4194
rect 5388 218 5400 4194
rect 5342 206 5400 218
rect 5500 4194 5558 4206
rect 5500 218 5512 4194
rect 5546 218 5558 4194
rect 5500 206 5558 218
rect 5658 4194 5716 4206
rect 5658 218 5670 4194
rect 5704 218 5716 4194
rect 5658 206 5716 218
rect 5816 4194 5874 4206
rect 5816 218 5828 4194
rect 5862 218 5874 4194
rect 5816 206 5874 218
<< mvpdiff >>
rect 588 8734 646 8746
rect 588 6758 600 8734
rect 634 6758 646 8734
rect 588 6746 646 6758
rect 746 8734 804 8746
rect 746 6758 758 8734
rect 792 6758 804 8734
rect 746 6746 804 6758
rect 904 8734 962 8746
rect 904 6758 916 8734
rect 950 6758 962 8734
rect 904 6746 962 6758
rect 1062 8734 1120 8746
rect 1062 6758 1074 8734
rect 1108 6758 1120 8734
rect 1062 6746 1120 6758
rect 1220 8734 1278 8746
rect 1220 6758 1232 8734
rect 1266 6758 1278 8734
rect 1220 6746 1278 6758
rect 1378 8734 1436 8746
rect 1378 6758 1390 8734
rect 1424 6758 1436 8734
rect 1378 6746 1436 6758
rect 1536 8734 1594 8746
rect 1536 6758 1548 8734
rect 1582 6758 1594 8734
rect 1536 6746 1594 6758
rect 1694 8734 1752 8746
rect 1694 6758 1706 8734
rect 1740 6758 1752 8734
rect 1694 6746 1752 6758
rect 1852 8734 1910 8746
rect 1852 6758 1864 8734
rect 1898 6758 1910 8734
rect 1852 6746 1910 6758
rect 2010 8734 2068 8746
rect 2010 6758 2022 8734
rect 2056 6758 2068 8734
rect 2010 6746 2068 6758
rect 2168 8734 2226 8746
rect 2168 6758 2180 8734
rect 2214 6758 2226 8734
rect 2656 8742 2714 8754
rect 2168 6746 2226 6758
rect 2656 4766 2668 8742
rect 2702 4766 2714 8742
rect 2656 4754 2714 4766
rect 2814 8742 2872 8754
rect 2814 4766 2826 8742
rect 2860 4766 2872 8742
rect 2814 4754 2872 4766
rect 2972 8742 3030 8754
rect 2972 4766 2984 8742
rect 3018 4766 3030 8742
rect 2972 4754 3030 4766
rect 3130 8742 3188 8754
rect 3130 4766 3142 8742
rect 3176 4766 3188 8742
rect 3130 4754 3188 4766
rect 3288 8742 3346 8754
rect 3288 4766 3300 8742
rect 3334 4766 3346 8742
rect 3288 4754 3346 4766
rect 3446 8742 3504 8754
rect 3446 4766 3458 8742
rect 3492 4766 3504 8742
rect 3446 4754 3504 4766
rect 3604 8742 3662 8754
rect 3604 4766 3616 8742
rect 3650 4766 3662 8742
rect 3604 4754 3662 4766
rect 3762 8742 3820 8754
rect 3762 4766 3774 8742
rect 3808 4766 3820 8742
rect 3762 4754 3820 4766
rect 3920 8742 3978 8754
rect 3920 4766 3932 8742
rect 3966 4766 3978 8742
rect 3920 4754 3978 4766
rect 4078 8742 4136 8754
rect 4078 4766 4090 8742
rect 4124 4766 4136 8742
rect 4078 4754 4136 4766
rect 4236 8742 4294 8754
rect 4236 4766 4248 8742
rect 4282 4766 4294 8742
rect 4236 4754 4294 4766
rect 4394 8742 4452 8754
rect 4394 4766 4406 8742
rect 4440 4766 4452 8742
rect 4394 4754 4452 4766
rect 4552 8742 4610 8754
rect 4552 4766 4564 8742
rect 4598 4766 4610 8742
rect 4552 4754 4610 4766
rect 4710 8742 4768 8754
rect 4710 4766 4722 8742
rect 4756 4766 4768 8742
rect 4710 4754 4768 4766
rect 4868 8742 4926 8754
rect 4868 4766 4880 8742
rect 4914 4766 4926 8742
rect 4868 4754 4926 4766
rect 5026 8742 5084 8754
rect 5026 4766 5038 8742
rect 5072 4766 5084 8742
rect 5026 4754 5084 4766
rect 5184 8742 5242 8754
rect 5184 4766 5196 8742
rect 5230 4766 5242 8742
rect 5184 4754 5242 4766
rect 5342 8742 5400 8754
rect 5342 4766 5354 8742
rect 5388 4766 5400 8742
rect 5342 4754 5400 4766
rect 5500 8742 5558 8754
rect 5500 4766 5512 8742
rect 5546 4766 5558 8742
rect 5500 4754 5558 4766
rect 5658 8742 5716 8754
rect 5658 4766 5670 8742
rect 5704 4766 5716 8742
rect 5658 4754 5716 4766
rect 5816 8742 5874 8754
rect 5816 4766 5828 8742
rect 5862 4766 5874 8742
rect 5816 4754 5874 4766
rect 1602 2760 1660 2772
rect 1602 2384 1614 2760
rect 1648 2384 1660 2760
rect 1602 2372 1660 2384
rect 1760 2760 1818 2772
rect 1760 2384 1772 2760
rect 1806 2384 1818 2760
rect 1760 2372 1818 2384
rect 1892 2760 1950 2772
rect 1892 2384 1904 2760
rect 1938 2384 1950 2760
rect 1892 2372 1950 2384
rect 2050 2760 2108 2772
rect 2050 2384 2062 2760
rect 2096 2384 2108 2760
rect 2050 2372 2108 2384
<< ndiffc >>
rect 563 3797 597 3973
rect 659 3797 693 3973
rect 755 3797 789 3973
rect 851 3797 885 3973
rect 947 3797 981 3973
rect 1043 3797 1077 3973
<< pdiffc >>
rect 563 3346 597 3522
rect 659 3346 693 3522
rect 755 3346 789 3522
rect 851 3346 885 3522
rect 947 3346 981 3522
rect 1043 3346 1077 3522
<< mvndiffc >>
rect 600 4332 634 6308
rect 758 4332 792 6308
rect 916 4332 950 6308
rect 1074 4332 1108 6308
rect 1232 4332 1266 6308
rect 1390 4332 1424 6308
rect 1548 4332 1582 6308
rect 1706 4332 1740 6308
rect 1864 4332 1898 6308
rect 2022 4332 2056 6308
rect 2180 4332 2214 6308
rect 1302 3144 1336 3920
rect 1460 3144 1494 3920
rect 1618 3144 1652 3920
rect 1776 3144 1810 3920
rect 1916 3144 1950 3920
rect 2074 3144 2108 3920
rect 2232 3144 2266 3920
rect 2390 3144 2424 3920
rect 2668 218 2702 4194
rect 2826 218 2860 4194
rect 2984 218 3018 4194
rect 3142 218 3176 4194
rect 3300 218 3334 4194
rect 3458 218 3492 4194
rect 3616 218 3650 4194
rect 3774 218 3808 4194
rect 3932 218 3966 4194
rect 4090 218 4124 4194
rect 4248 218 4282 4194
rect 4406 218 4440 4194
rect 4564 218 4598 4194
rect 4722 218 4756 4194
rect 4880 218 4914 4194
rect 5038 218 5072 4194
rect 5196 218 5230 4194
rect 5354 218 5388 4194
rect 5512 218 5546 4194
rect 5670 218 5704 4194
rect 5828 218 5862 4194
<< mvpdiffc >>
rect 600 6758 634 8734
rect 758 6758 792 8734
rect 916 6758 950 8734
rect 1074 6758 1108 8734
rect 1232 6758 1266 8734
rect 1390 6758 1424 8734
rect 1548 6758 1582 8734
rect 1706 6758 1740 8734
rect 1864 6758 1898 8734
rect 2022 6758 2056 8734
rect 2180 6758 2214 8734
rect 2668 4766 2702 8742
rect 2826 4766 2860 8742
rect 2984 4766 3018 8742
rect 3142 4766 3176 8742
rect 3300 4766 3334 8742
rect 3458 4766 3492 8742
rect 3616 4766 3650 8742
rect 3774 4766 3808 8742
rect 3932 4766 3966 8742
rect 4090 4766 4124 8742
rect 4248 4766 4282 8742
rect 4406 4766 4440 8742
rect 4564 4766 4598 8742
rect 4722 4766 4756 8742
rect 4880 4766 4914 8742
rect 5038 4766 5072 8742
rect 5196 4766 5230 8742
rect 5354 4766 5388 8742
rect 5512 4766 5546 8742
rect 5670 4766 5704 8742
rect 5828 4766 5862 8742
rect 1614 2384 1648 2760
rect 1772 2384 1806 2760
rect 1904 2384 1938 2760
rect 2062 2384 2096 2760
<< psubdiff >>
rect 596 4043 620 4082
rect 1035 4043 1059 4082
<< nsubdiff >>
rect 558 3227 625 3261
rect 1014 3227 1085 3261
<< mvpsubdiff >>
rect 660 4160 684 4228
rect 2122 4160 2226 4228
rect 1340 4016 1364 4106
rect 2364 4016 2388 4106
rect 2530 2746 2582 2770
rect 2530 1774 2582 1798
rect 5948 2794 6000 2818
rect 5948 1822 6000 1846
rect 2610 8 2634 114
rect 5898 8 5922 114
<< mvnsubdiff >>
rect 666 8812 696 8864
rect 2104 8812 2148 8864
rect 2732 8810 2762 8864
rect 5752 8810 5802 8864
rect 2538 7282 2592 7330
rect 2590 6334 2592 7282
rect 2538 6282 2592 6334
rect 5928 7360 5982 7412
rect 5928 6412 5930 7360
rect 5928 6364 5982 6412
rect 1634 2266 1674 2308
rect 2052 2266 2086 2308
<< psubdiffcont >>
rect 620 4043 1035 4082
<< nsubdiffcont >>
rect 625 3227 1014 3261
<< mvpsubdiffcont >>
rect 684 4160 2122 4228
rect 1364 4016 2364 4106
rect 2530 1798 2582 2746
rect 5948 1846 6000 2794
rect 2634 8 5898 114
<< mvnsubdiffcont >>
rect 696 8812 2104 8864
rect 2762 8810 5752 8864
rect 2538 6334 2590 7282
rect 5930 6412 5982 7360
rect 1674 2266 2052 2308
<< poly >>
rect 646 8746 746 8772
rect 804 8746 904 8772
rect 962 8746 1062 8772
rect 1120 8746 1220 8772
rect 1278 8746 1378 8772
rect 1436 8746 1536 8772
rect 1594 8746 1694 8772
rect 1752 8746 1852 8772
rect 1910 8746 2010 8772
rect 2068 8746 2168 8772
rect 2714 8754 2814 8780
rect 2872 8754 2972 8780
rect 3030 8754 3130 8780
rect 3188 8754 3288 8780
rect 3346 8754 3446 8780
rect 3504 8754 3604 8780
rect 3662 8754 3762 8780
rect 3820 8754 3920 8780
rect 3978 8754 4078 8780
rect 4136 8754 4236 8780
rect 4294 8754 4394 8780
rect 4452 8754 4552 8780
rect 4610 8754 4710 8780
rect 4768 8754 4868 8780
rect 4926 8754 5026 8780
rect 5084 8754 5184 8780
rect 5242 8754 5342 8780
rect 5400 8754 5500 8780
rect 5558 8754 5658 8780
rect 5716 8754 5816 8780
rect 646 6720 746 6746
rect 804 6720 904 6746
rect 962 6720 1062 6746
rect 1120 6720 1220 6746
rect 1278 6720 1378 6746
rect 1436 6720 1536 6746
rect 1594 6720 1694 6746
rect 1752 6720 1852 6746
rect 1910 6720 2010 6746
rect 2068 6720 2168 6746
rect 666 6674 726 6720
rect 824 6676 884 6720
rect 982 6676 1042 6720
rect 662 6658 728 6674
rect 662 6624 678 6658
rect 712 6624 728 6658
rect 662 6608 728 6624
rect 824 6660 1042 6676
rect 824 6626 916 6660
rect 950 6626 1042 6660
rect 824 6610 1042 6626
rect 824 6608 884 6610
rect 982 6608 1042 6610
rect 1140 6676 1200 6720
rect 1298 6676 1358 6720
rect 1140 6660 1358 6676
rect 1140 6626 1230 6660
rect 1264 6626 1358 6660
rect 1140 6610 1358 6626
rect 1140 6608 1200 6610
rect 1298 6608 1358 6610
rect 1456 6674 1516 6720
rect 1614 6674 1674 6720
rect 1456 6658 1674 6674
rect 1456 6624 1548 6658
rect 1582 6624 1674 6658
rect 1456 6608 1674 6624
rect 1772 6674 1832 6720
rect 1930 6674 1990 6720
rect 1772 6658 1990 6674
rect 1772 6624 1862 6658
rect 1896 6624 1990 6658
rect 1772 6608 1990 6624
rect 2088 6674 2148 6720
rect 2088 6658 2156 6674
rect 2088 6624 2106 6658
rect 2140 6624 2156 6658
rect 2088 6608 2156 6624
rect 666 6602 726 6608
rect 2088 6602 2148 6608
rect 666 6456 726 6462
rect 662 6440 728 6456
rect 662 6406 678 6440
rect 712 6406 728 6440
rect 662 6390 728 6406
rect 824 6442 1042 6458
rect 824 6408 916 6442
rect 950 6408 1042 6442
rect 824 6392 1042 6408
rect 666 6346 726 6390
rect 824 6346 884 6392
rect 982 6346 1042 6392
rect 1140 6442 1358 6458
rect 1140 6408 1230 6442
rect 1264 6408 1358 6442
rect 1140 6392 1358 6408
rect 1140 6346 1200 6392
rect 1298 6346 1358 6392
rect 1456 6456 1516 6458
rect 1614 6456 1674 6458
rect 1456 6440 1674 6456
rect 1456 6406 1548 6440
rect 1582 6406 1674 6440
rect 1456 6390 1674 6406
rect 1456 6346 1516 6390
rect 1614 6346 1674 6390
rect 1772 6456 1832 6458
rect 1930 6456 1990 6458
rect 1772 6440 1990 6456
rect 1772 6406 1862 6440
rect 1896 6406 1990 6440
rect 1772 6390 1990 6406
rect 1772 6346 1832 6390
rect 1930 6346 1990 6390
rect 2088 6456 2148 6462
rect 2088 6440 2156 6456
rect 2088 6406 2106 6440
rect 2140 6406 2156 6440
rect 2088 6390 2156 6406
rect 2088 6346 2148 6390
rect 646 6320 746 6346
rect 804 6320 904 6346
rect 962 6320 1062 6346
rect 1120 6320 1220 6346
rect 1278 6320 1378 6346
rect 1436 6320 1536 6346
rect 1594 6320 1694 6346
rect 1752 6320 1852 6346
rect 1910 6320 2010 6346
rect 2068 6320 2168 6346
rect 2714 4728 2814 4754
rect 2872 4728 2972 4754
rect 3030 4728 3130 4754
rect 3188 4728 3288 4754
rect 3346 4728 3446 4754
rect 3504 4728 3604 4754
rect 3662 4728 3762 4754
rect 3820 4728 3920 4754
rect 3978 4728 4078 4754
rect 4136 4728 4236 4754
rect 4294 4728 4394 4754
rect 4452 4728 4552 4754
rect 4610 4728 4710 4754
rect 4768 4728 4868 4754
rect 4926 4728 5026 4754
rect 5084 4728 5184 4754
rect 5242 4728 5342 4754
rect 5400 4728 5500 4754
rect 5558 4728 5658 4754
rect 5716 4728 5816 4754
rect 2734 4666 2794 4728
rect 2722 4650 2794 4666
rect 2722 4616 2738 4650
rect 2772 4616 2794 4650
rect 2722 4600 2794 4616
rect 646 4294 746 4320
rect 804 4294 904 4320
rect 962 4294 1062 4320
rect 1120 4294 1220 4320
rect 1278 4294 1378 4320
rect 1436 4294 1536 4320
rect 1594 4294 1694 4320
rect 1752 4294 1852 4320
rect 1910 4294 2010 4320
rect 2068 4294 2168 4320
rect 2734 4232 2794 4600
rect 2892 4666 2952 4728
rect 3050 4666 3110 4728
rect 2892 4650 3110 4666
rect 2892 4616 2982 4650
rect 3016 4616 3110 4650
rect 2892 4600 3110 4616
rect 2892 4232 2952 4600
rect 3050 4232 3110 4600
rect 3208 4666 3268 4728
rect 3366 4666 3426 4728
rect 3208 4650 3426 4666
rect 3208 4616 3298 4650
rect 3332 4616 3426 4650
rect 3208 4600 3426 4616
rect 3208 4232 3268 4600
rect 3366 4232 3426 4600
rect 3524 4666 3584 4728
rect 3682 4666 3742 4728
rect 3524 4650 3742 4666
rect 3524 4616 3614 4650
rect 3648 4616 3742 4650
rect 3524 4600 3742 4616
rect 3524 4232 3584 4600
rect 3682 4232 3742 4600
rect 3840 4666 3900 4728
rect 3998 4666 4058 4728
rect 3840 4650 4058 4666
rect 3840 4616 3930 4650
rect 3964 4616 4058 4650
rect 3840 4600 4058 4616
rect 3840 4232 3900 4600
rect 3998 4232 4058 4600
rect 4156 4666 4216 4728
rect 4314 4666 4374 4728
rect 4156 4650 4374 4666
rect 4156 4616 4248 4650
rect 4282 4616 4374 4650
rect 4156 4600 4374 4616
rect 4156 4232 4216 4600
rect 4314 4232 4374 4600
rect 4472 4666 4532 4728
rect 4630 4666 4690 4728
rect 4472 4650 4690 4666
rect 4472 4616 4564 4650
rect 4598 4616 4690 4650
rect 4472 4600 4690 4616
rect 4472 4232 4532 4600
rect 4630 4232 4690 4600
rect 4788 4666 4848 4728
rect 4946 4666 5006 4728
rect 4788 4650 5006 4666
rect 4788 4616 4878 4650
rect 4912 4616 5006 4650
rect 4788 4600 5006 4616
rect 4788 4232 4848 4600
rect 4946 4232 5006 4600
rect 5104 4666 5164 4728
rect 5262 4666 5322 4728
rect 5104 4650 5322 4666
rect 5104 4616 5194 4650
rect 5228 4616 5322 4650
rect 5104 4600 5322 4616
rect 5104 4232 5164 4600
rect 5262 4232 5322 4600
rect 5420 4666 5480 4728
rect 5578 4666 5638 4728
rect 5420 4650 5638 4666
rect 5420 4616 5512 4650
rect 5546 4616 5638 4650
rect 5420 4600 5638 4616
rect 5420 4232 5480 4600
rect 5578 4232 5638 4600
rect 5736 4666 5796 4728
rect 5736 4650 5820 4666
rect 5736 4616 5770 4650
rect 5804 4616 5820 4650
rect 5736 4600 5820 4616
rect 5736 4232 5796 4600
rect 2714 4206 2814 4232
rect 2872 4206 2972 4232
rect 3030 4206 3130 4232
rect 3188 4206 3288 4232
rect 3346 4206 3446 4232
rect 3504 4206 3604 4232
rect 3662 4206 3762 4232
rect 3820 4206 3920 4232
rect 3978 4206 4078 4232
rect 4136 4206 4236 4232
rect 4294 4206 4394 4232
rect 4452 4206 4552 4232
rect 4610 4206 4710 4232
rect 4768 4206 4868 4232
rect 4926 4206 5026 4232
rect 5084 4206 5184 4232
rect 5242 4206 5342 4232
rect 5400 4206 5500 4232
rect 5558 4206 5658 4232
rect 5716 4206 5816 4232
rect 613 3985 643 4011
rect 709 3985 739 4011
rect 805 3985 835 4011
rect 901 3985 931 4011
rect 997 3985 1027 4011
rect 1348 3932 1448 3958
rect 1506 3932 1606 3958
rect 1664 3932 1764 3958
rect 1962 3932 2062 3958
rect 2120 3932 2220 3958
rect 2278 3932 2378 3958
rect 613 3634 643 3785
rect 563 3618 643 3634
rect 563 3584 579 3618
rect 613 3584 643 3618
rect 563 3568 643 3584
rect 613 3534 643 3568
rect 709 3634 739 3785
rect 805 3634 835 3785
rect 709 3618 835 3634
rect 709 3584 755 3618
rect 789 3584 835 3618
rect 709 3568 835 3584
rect 709 3534 739 3568
rect 805 3534 835 3568
rect 901 3631 931 3785
rect 997 3631 1027 3785
rect 901 3615 1027 3631
rect 901 3581 947 3615
rect 981 3581 1027 3615
rect 901 3565 1027 3581
rect 901 3534 931 3565
rect 997 3534 1027 3565
rect 613 3308 643 3334
rect 709 3303 739 3334
rect 805 3308 835 3334
rect 901 3303 931 3334
rect 997 3308 1027 3334
rect 1348 3106 1448 3132
rect 1506 3106 1606 3132
rect 1664 3106 1764 3132
rect 1962 3106 2062 3132
rect 2120 3106 2220 3132
rect 2278 3106 2378 3132
rect 1366 3092 1432 3106
rect 1366 3058 1382 3092
rect 1416 3058 1432 3092
rect 1366 3042 1432 3058
rect 1524 3094 1590 3106
rect 1524 3060 1540 3094
rect 1574 3060 1590 3094
rect 1524 3044 1590 3060
rect 1684 3094 1750 3106
rect 1684 3060 1700 3094
rect 1734 3060 1750 3094
rect 1684 3044 1750 3060
rect 1978 3094 2044 3106
rect 1978 3060 1994 3094
rect 2028 3060 2044 3094
rect 1978 3044 2044 3060
rect 2140 3094 2206 3106
rect 2140 3060 2156 3094
rect 2190 3060 2206 3094
rect 2140 3044 2206 3060
rect 2296 3094 2362 3106
rect 2296 3060 2312 3094
rect 2346 3060 2362 3094
rect 2296 3044 2362 3060
rect 1660 2853 1760 2869
rect 1660 2819 1676 2853
rect 1744 2819 1760 2853
rect 1660 2772 1760 2819
rect 1950 2853 2050 2869
rect 1950 2819 1966 2853
rect 2034 2819 2050 2853
rect 1950 2772 2050 2819
rect 1660 2346 1760 2372
rect 1950 2346 2050 2372
rect 2714 180 2814 206
rect 2872 180 2972 206
rect 3030 180 3130 206
rect 3188 180 3288 206
rect 3346 180 3446 206
rect 3504 180 3604 206
rect 3662 180 3762 206
rect 3820 180 3920 206
rect 3978 180 4078 206
rect 4136 180 4236 206
rect 4294 180 4394 206
rect 4452 180 4552 206
rect 4610 180 4710 206
rect 4768 180 4868 206
rect 4926 180 5026 206
rect 5084 180 5184 206
rect 5242 180 5342 206
rect 5400 180 5500 206
rect 5558 180 5658 206
rect 5716 180 5816 206
<< polycont >>
rect 678 6624 712 6658
rect 916 6626 950 6660
rect 1230 6626 1264 6660
rect 1548 6624 1582 6658
rect 1862 6624 1896 6658
rect 2106 6624 2140 6658
rect 678 6406 712 6440
rect 916 6408 950 6442
rect 1230 6408 1264 6442
rect 1548 6406 1582 6440
rect 1862 6406 1896 6440
rect 2106 6406 2140 6440
rect 2738 4616 2772 4650
rect 2982 4616 3016 4650
rect 3298 4616 3332 4650
rect 3614 4616 3648 4650
rect 3930 4616 3964 4650
rect 4248 4616 4282 4650
rect 4564 4616 4598 4650
rect 4878 4616 4912 4650
rect 5194 4616 5228 4650
rect 5512 4616 5546 4650
rect 5770 4616 5804 4650
rect 579 3584 613 3618
rect 755 3584 789 3618
rect 947 3581 981 3615
rect 1382 3058 1416 3092
rect 1540 3060 1574 3094
rect 1700 3060 1734 3094
rect 1994 3060 2028 3094
rect 2156 3060 2190 3094
rect 2312 3060 2346 3094
rect 1676 2819 1744 2853
rect 1966 2819 2034 2853
<< locali >>
rect 674 8812 696 8864
rect 2104 8812 2140 8864
rect 2740 8810 2762 8864
rect 5752 8810 5794 8864
rect 600 8734 634 8750
rect 600 6742 634 6758
rect 758 8734 792 8750
rect 758 6742 792 6758
rect 916 8734 950 8750
rect 916 6742 950 6758
rect 1074 8734 1108 8750
rect 1074 6742 1108 6758
rect 1232 8734 1266 8750
rect 1232 6742 1266 6758
rect 1390 8734 1424 8750
rect 1390 6742 1424 6758
rect 1548 8734 1582 8750
rect 1548 6742 1582 6758
rect 1706 8734 1740 8750
rect 1706 6742 1740 6758
rect 1864 8734 1898 8750
rect 1864 6742 1898 6758
rect 2022 8734 2056 8750
rect 2022 6742 2056 6758
rect 2180 8734 2214 8750
rect 2668 8742 2702 8758
rect 2180 6742 2214 6758
rect 2538 7282 2592 7322
rect 662 6624 678 6658
rect 712 6624 728 6658
rect 900 6626 916 6660
rect 950 6626 966 6660
rect 1214 6626 1230 6660
rect 1264 6626 1280 6660
rect 1532 6624 1548 6658
rect 1582 6624 1598 6658
rect 1846 6624 1862 6658
rect 1896 6624 1912 6658
rect 2090 6624 2106 6658
rect 2140 6624 2156 6658
rect 662 6406 678 6440
rect 712 6406 728 6440
rect 900 6408 916 6442
rect 950 6408 966 6442
rect 1214 6408 1230 6442
rect 1264 6408 1280 6442
rect 1532 6406 1548 6440
rect 1582 6406 1598 6440
rect 1846 6406 1862 6440
rect 1896 6406 1912 6440
rect 2090 6406 2106 6440
rect 2140 6406 2156 6440
rect 2590 6334 2592 7282
rect 600 6308 634 6324
rect 600 4316 634 4332
rect 758 6308 792 6324
rect 758 4316 792 4332
rect 916 6308 950 6324
rect 916 4316 950 4332
rect 1074 6308 1108 6324
rect 1074 4316 1108 4332
rect 1232 6308 1266 6324
rect 1232 4316 1266 4332
rect 1390 6308 1424 6324
rect 1390 4316 1424 4332
rect 1548 6308 1582 6324
rect 1548 4316 1582 4332
rect 1706 6308 1740 6324
rect 1706 4316 1740 4332
rect 1864 6308 1898 6324
rect 1864 4316 1898 4332
rect 2022 6308 2056 6324
rect 2022 4316 2056 4332
rect 2180 6308 2214 6324
rect 2538 6290 2592 6334
rect 2668 4750 2702 4766
rect 2826 8742 2860 8758
rect 2826 4750 2860 4766
rect 2984 8742 3018 8758
rect 2984 4750 3018 4766
rect 3142 8742 3176 8758
rect 3142 4750 3176 4766
rect 3300 8742 3334 8758
rect 3300 4750 3334 4766
rect 3458 8742 3492 8758
rect 3458 4750 3492 4766
rect 3616 8742 3650 8758
rect 3616 4750 3650 4766
rect 3774 8742 3808 8758
rect 3774 4750 3808 4766
rect 3932 8742 3966 8758
rect 3932 4750 3966 4766
rect 4090 8742 4124 8758
rect 4090 4750 4124 4766
rect 4248 8742 4282 8758
rect 4248 4750 4282 4766
rect 4406 8742 4440 8758
rect 4406 4750 4440 4766
rect 4564 8742 4598 8758
rect 4564 4750 4598 4766
rect 4722 8742 4756 8758
rect 4722 4750 4756 4766
rect 4880 8742 4914 8758
rect 4880 4750 4914 4766
rect 5038 8742 5072 8758
rect 5038 4750 5072 4766
rect 5196 8742 5230 8758
rect 5196 4750 5230 4766
rect 5354 8742 5388 8758
rect 5354 4750 5388 4766
rect 5512 8742 5546 8758
rect 5512 4750 5546 4766
rect 5670 8742 5704 8758
rect 5670 4750 5704 4766
rect 5828 8742 5862 8758
rect 5928 7360 5982 7404
rect 5928 6412 5930 7360
rect 5928 6372 5982 6412
rect 5828 4750 5862 4766
rect 2722 4616 2738 4650
rect 2772 4616 2788 4650
rect 2966 4616 2982 4650
rect 3016 4616 3032 4650
rect 3282 4616 3298 4650
rect 3332 4616 3348 4650
rect 3598 4616 3614 4650
rect 3648 4616 3664 4650
rect 3914 4616 3930 4650
rect 3964 4616 3980 4650
rect 4232 4616 4248 4650
rect 4282 4616 4298 4650
rect 4548 4616 4564 4650
rect 4598 4616 4614 4650
rect 4862 4616 4878 4650
rect 4912 4616 4928 4650
rect 5178 4616 5194 4650
rect 5228 4616 5244 4650
rect 5496 4616 5512 4650
rect 5546 4616 5562 4650
rect 5754 4616 5770 4650
rect 5804 4616 5820 4650
rect 2180 4316 2214 4332
rect 668 4160 684 4228
rect 2122 4160 2138 4228
rect 2668 4194 2702 4210
rect 1348 4016 1364 4106
rect 2364 4016 2380 4106
rect 563 3973 597 3989
rect 563 3781 597 3797
rect 659 3973 693 3989
rect 659 3781 693 3797
rect 755 3973 789 3989
rect 755 3781 789 3797
rect 851 3973 885 3989
rect 851 3781 885 3797
rect 947 3973 981 3989
rect 947 3781 981 3797
rect 1043 3973 1077 3989
rect 1043 3781 1077 3797
rect 1302 3920 1336 3936
rect 563 3584 579 3618
rect 613 3584 629 3618
rect 739 3584 755 3618
rect 789 3584 805 3618
rect 931 3581 947 3615
rect 981 3581 997 3615
rect 563 3522 597 3538
rect 563 3330 597 3346
rect 659 3522 693 3538
rect 659 3330 693 3346
rect 755 3522 789 3538
rect 755 3330 789 3346
rect 851 3522 885 3538
rect 851 3330 885 3346
rect 947 3522 981 3538
rect 947 3330 981 3346
rect 1043 3522 1077 3538
rect 1043 3330 1077 3346
rect 1302 3128 1336 3144
rect 1460 3920 1494 3936
rect 1460 3128 1494 3144
rect 1618 3920 1652 3936
rect 1618 3128 1652 3144
rect 1776 3920 1810 3936
rect 1776 3128 1810 3144
rect 1916 3920 1950 3936
rect 1916 3128 1950 3144
rect 2074 3920 2108 3936
rect 2074 3128 2108 3144
rect 2232 3920 2266 3936
rect 2232 3128 2266 3144
rect 2390 3920 2424 3936
rect 2390 3128 2424 3144
rect 1366 3058 1382 3092
rect 1416 3058 1432 3092
rect 1524 3060 1540 3094
rect 1574 3060 1590 3094
rect 1684 3060 1700 3094
rect 1734 3060 1750 3094
rect 1978 3060 1994 3094
rect 2028 3060 2044 3094
rect 2140 3060 2156 3094
rect 2190 3060 2206 3094
rect 2296 3060 2312 3094
rect 2346 3060 2362 3094
rect 1660 2819 1676 2853
rect 1744 2819 1760 2853
rect 1950 2819 1966 2853
rect 2034 2819 2050 2853
rect 1614 2760 1648 2776
rect 1614 2368 1648 2384
rect 1772 2760 1806 2776
rect 1772 2368 1806 2384
rect 1904 2760 1938 2776
rect 1904 2368 1938 2384
rect 2062 2760 2096 2776
rect 2062 2368 2096 2384
rect 2530 2746 2582 2762
rect 1642 2266 1674 2308
rect 2052 2266 2078 2308
rect 2530 1782 2582 1798
rect 2668 202 2702 218
rect 2826 4194 2860 4210
rect 2826 202 2860 218
rect 2984 4194 3018 4210
rect 2984 202 3018 218
rect 3142 4194 3176 4210
rect 3142 202 3176 218
rect 3300 4194 3334 4210
rect 3300 202 3334 218
rect 3458 4194 3492 4210
rect 3458 202 3492 218
rect 3616 4194 3650 4210
rect 3616 202 3650 218
rect 3774 4194 3808 4210
rect 3774 202 3808 218
rect 3932 4194 3966 4210
rect 3932 202 3966 218
rect 4090 4194 4124 4210
rect 4090 202 4124 218
rect 4248 4194 4282 4210
rect 4248 202 4282 218
rect 4406 4194 4440 4210
rect 4406 202 4440 218
rect 4564 4194 4598 4210
rect 4564 202 4598 218
rect 4722 4194 4756 4210
rect 4722 202 4756 218
rect 4880 4194 4914 4210
rect 4880 202 4914 218
rect 5038 4194 5072 4210
rect 5038 202 5072 218
rect 5196 4194 5230 4210
rect 5196 202 5230 218
rect 5354 4194 5388 4210
rect 5354 202 5388 218
rect 5512 4194 5546 4210
rect 5512 202 5546 218
rect 5670 4194 5704 4210
rect 5670 202 5704 218
rect 5828 4194 5862 4210
rect 5948 2794 6000 2810
rect 5948 1830 6000 1846
rect 5828 202 5862 218
rect 2618 8 2634 114
rect 5898 8 5914 114
<< viali >>
rect 696 8812 2104 8864
rect 2762 8810 5752 8864
rect 600 6758 634 8734
rect 758 6758 792 8734
rect 916 6758 950 8734
rect 1074 6758 1108 8734
rect 1232 6758 1266 8734
rect 1390 6758 1424 8734
rect 1548 6758 1582 8734
rect 1706 6758 1740 8734
rect 1864 6758 1898 8734
rect 2022 6758 2056 8734
rect 2180 6758 2214 8734
rect 678 6624 712 6658
rect 916 6626 950 6660
rect 1230 6626 1264 6660
rect 1548 6624 1582 6658
rect 1862 6624 1896 6658
rect 2106 6624 2140 6658
rect 678 6406 712 6440
rect 916 6408 950 6442
rect 1230 6408 1264 6442
rect 1548 6406 1582 6440
rect 1862 6406 1896 6440
rect 2106 6406 2140 6440
rect 2538 6334 2590 7282
rect 600 4332 634 6308
rect 758 4332 792 6308
rect 916 4332 950 6308
rect 1074 4332 1108 6308
rect 1232 4332 1266 6308
rect 1390 4332 1424 6308
rect 1548 4332 1582 6308
rect 1706 4332 1740 6308
rect 1864 4332 1898 6308
rect 2022 4332 2056 6308
rect 2180 4332 2214 6308
rect 2668 4766 2702 8742
rect 2826 4766 2860 8742
rect 2984 4766 3018 8742
rect 3142 4766 3176 8742
rect 3300 4766 3334 8742
rect 3458 4766 3492 8742
rect 3616 4766 3650 8742
rect 3774 4766 3808 8742
rect 3932 4766 3966 8742
rect 4090 4766 4124 8742
rect 4248 4766 4282 8742
rect 4406 4766 4440 8742
rect 4564 4766 4598 8742
rect 4722 4766 4756 8742
rect 4880 4766 4914 8742
rect 5038 4766 5072 8742
rect 5196 4766 5230 8742
rect 5354 4766 5388 8742
rect 5512 4766 5546 8742
rect 5670 4766 5704 8742
rect 5828 4766 5862 8742
rect 5930 6412 5982 7360
rect 2738 4616 2772 4650
rect 2982 4616 3016 4650
rect 3298 4616 3332 4650
rect 3614 4616 3648 4650
rect 3930 4616 3964 4650
rect 4248 4616 4282 4650
rect 4564 4616 4598 4650
rect 4878 4616 4912 4650
rect 5194 4616 5228 4650
rect 5512 4616 5546 4650
rect 5770 4616 5804 4650
rect 684 4162 2122 4228
rect 555 4082 1077 4086
rect 555 4043 620 4082
rect 620 4043 1035 4082
rect 1035 4043 1077 4082
rect 555 4040 1077 4043
rect 1364 4016 2364 4106
rect 563 3797 597 3973
rect 659 3797 693 3973
rect 755 3797 789 3973
rect 851 3797 885 3973
rect 947 3797 981 3973
rect 1043 3797 1077 3973
rect 579 3584 613 3618
rect 755 3584 789 3618
rect 947 3581 981 3615
rect 563 3346 597 3522
rect 659 3346 693 3522
rect 755 3346 789 3522
rect 851 3346 885 3522
rect 947 3346 981 3522
rect 1043 3346 1077 3522
rect 552 3261 1087 3262
rect 552 3227 625 3261
rect 625 3227 1014 3261
rect 1014 3227 1087 3261
rect 552 3226 1087 3227
rect 1302 3144 1336 3920
rect 1460 3144 1494 3920
rect 1618 3144 1652 3920
rect 1776 3144 1810 3920
rect 1916 3144 1950 3920
rect 2074 3144 2108 3920
rect 2232 3144 2266 3920
rect 2390 3144 2424 3920
rect 1382 3058 1416 3092
rect 1540 3060 1574 3094
rect 1700 3060 1734 3094
rect 1994 3060 2028 3094
rect 2156 3060 2190 3094
rect 2312 3060 2346 3094
rect 1676 2819 1744 2853
rect 1966 2819 2034 2853
rect 1614 2384 1648 2760
rect 1772 2384 1806 2760
rect 1904 2384 1938 2760
rect 2062 2384 2096 2760
rect 1674 2266 2052 2308
rect 2668 218 2702 4194
rect 2826 218 2860 4194
rect 2984 218 3018 4194
rect 3142 218 3176 4194
rect 3300 218 3334 4194
rect 3458 218 3492 4194
rect 3616 218 3650 4194
rect 3774 218 3808 4194
rect 3932 218 3966 4194
rect 4090 218 4124 4194
rect 4248 218 4282 4194
rect 4406 218 4440 4194
rect 4564 218 4598 4194
rect 4722 218 4756 4194
rect 4880 218 4914 4194
rect 5038 218 5072 4194
rect 5196 218 5230 4194
rect 5354 218 5388 4194
rect 5512 218 5546 4194
rect 5670 218 5704 4194
rect 5828 218 5862 4194
rect 2634 8 5898 114
<< metal1 >>
rect 10 8898 150 8900
rect 10 8896 646 8898
rect 10 8874 5720 8896
rect 10 8864 5988 8874
rect 10 8812 696 8864
rect 2104 8812 2762 8864
rect 10 8810 2762 8812
rect 5752 8810 5988 8864
rect 10 8808 5988 8810
rect 10 7738 150 8808
rect 576 8806 5988 8808
rect 600 8746 634 8806
rect 916 8746 950 8806
rect 1232 8746 1266 8806
rect 1548 8746 1582 8806
rect 1864 8746 1898 8806
rect 2180 8746 2214 8806
rect 2532 8802 5988 8806
rect 594 8734 640 8746
rect 10 7140 152 7738
rect 12 2904 152 7140
rect 594 6758 600 8734
rect 634 6758 640 8734
rect 594 6746 640 6758
rect 752 8734 798 8746
rect 752 6758 758 8734
rect 792 6758 798 8734
rect 752 6746 798 6758
rect 910 8734 956 8746
rect 910 6758 916 8734
rect 950 6758 956 8734
rect 910 6746 956 6758
rect 1068 8734 1114 8746
rect 1068 6758 1074 8734
rect 1108 6758 1114 8734
rect 1068 6746 1114 6758
rect 1226 8734 1272 8746
rect 1226 6758 1232 8734
rect 1266 6758 1272 8734
rect 1226 6746 1272 6758
rect 1384 8734 1430 8746
rect 1384 6758 1390 8734
rect 1424 6758 1430 8734
rect 1384 6746 1430 6758
rect 1542 8734 1588 8746
rect 1542 6758 1548 8734
rect 1582 6758 1588 8734
rect 1542 6746 1588 6758
rect 1700 8734 1746 8746
rect 1700 6758 1706 8734
rect 1740 6758 1746 8734
rect 1700 6746 1746 6758
rect 1858 8734 1904 8746
rect 1858 6758 1864 8734
rect 1898 6758 1904 8734
rect 1858 6746 1904 6758
rect 2016 8734 2062 8746
rect 2016 6758 2022 8734
rect 2056 6758 2062 8734
rect 2016 6746 2062 6758
rect 2174 8734 2220 8746
rect 2174 6758 2180 8734
rect 2214 6758 2220 8734
rect 2174 6746 2220 6758
rect 2532 7284 2596 8802
rect 2666 8754 2700 8802
rect 2982 8754 3018 8802
rect 3298 8754 3334 8802
rect 3614 8754 3650 8802
rect 3930 8754 3966 8802
rect 4246 8754 4282 8802
rect 4562 8754 4598 8802
rect 4878 8754 4914 8802
rect 5194 8754 5230 8802
rect 5510 8754 5546 8802
rect 5826 8754 5862 8802
rect 2662 8742 2708 8754
rect 2662 7284 2668 8742
rect 2532 7282 2668 7284
rect 368 6694 508 6698
rect 368 6594 388 6694
rect 488 6594 508 6694
rect 658 6616 668 6668
rect 720 6616 730 6668
rect 190 6472 330 6482
rect 190 6372 208 6472
rect 308 6372 330 6472
rect 190 3652 330 6372
rect 190 3552 208 3652
rect 308 3552 330 3652
rect 190 3538 330 3552
rect 368 2998 508 6594
rect 758 6558 792 6746
rect 896 6616 906 6668
rect 958 6616 968 6668
rect 1074 6558 1108 6746
rect 1210 6616 1220 6668
rect 1272 6616 1282 6668
rect 1390 6558 1424 6746
rect 1528 6616 1538 6668
rect 1590 6616 1600 6668
rect 1706 6558 1740 6746
rect 1842 6616 1852 6668
rect 1904 6616 1914 6668
rect 2022 6558 2056 6746
rect 2086 6616 2096 6668
rect 2148 6616 2158 6668
rect 2330 6568 2340 6586
rect 738 6506 748 6558
rect 800 6506 810 6558
rect 1054 6506 1064 6558
rect 1116 6506 1126 6558
rect 1372 6506 1382 6558
rect 1434 6506 1444 6558
rect 1688 6506 1698 6558
rect 1750 6506 1760 6558
rect 2004 6506 2014 6558
rect 2066 6506 2076 6558
rect 658 6398 668 6450
rect 720 6398 730 6450
rect 758 6320 792 6506
rect 896 6398 906 6450
rect 958 6398 968 6450
rect 1074 6320 1108 6506
rect 1210 6398 1220 6450
rect 1272 6398 1282 6450
rect 1390 6320 1424 6506
rect 1528 6398 1538 6450
rect 1590 6398 1600 6450
rect 1706 6320 1740 6506
rect 1842 6398 1852 6450
rect 1904 6398 1914 6450
rect 2022 6320 2056 6506
rect 2324 6486 2340 6568
rect 2446 6568 2456 6586
rect 2446 6486 2464 6568
rect 2086 6398 2096 6450
rect 2148 6398 2158 6450
rect 594 6308 640 6320
rect 594 4332 600 6308
rect 634 4332 640 6308
rect 594 4320 640 4332
rect 752 6308 798 6320
rect 752 4332 758 6308
rect 792 4332 798 6308
rect 752 4320 798 4332
rect 910 6308 956 6320
rect 910 4332 916 6308
rect 950 4332 956 6308
rect 910 4320 956 4332
rect 1068 6308 1114 6320
rect 1068 4332 1074 6308
rect 1108 4332 1114 6308
rect 1068 4320 1114 4332
rect 1226 6308 1272 6320
rect 1226 4332 1232 6308
rect 1266 4332 1272 6308
rect 1226 4320 1272 4332
rect 1384 6308 1430 6320
rect 1384 4332 1390 6308
rect 1424 4332 1430 6308
rect 1384 4320 1430 4332
rect 1542 6308 1588 6320
rect 1542 4332 1548 6308
rect 1582 4332 1588 6308
rect 1542 4320 1588 4332
rect 1700 6308 1746 6320
rect 1700 4332 1706 6308
rect 1740 4332 1746 6308
rect 1700 4320 1746 4332
rect 1858 6308 1904 6320
rect 1858 4332 1864 6308
rect 1898 4332 1904 6308
rect 1858 4320 1904 4332
rect 2016 6308 2062 6320
rect 2016 4332 2022 6308
rect 2056 4332 2062 6308
rect 2016 4320 2062 4332
rect 2174 6308 2220 6320
rect 2174 4332 2180 6308
rect 2214 4332 2220 6308
rect 2324 4682 2464 6486
rect 2532 6334 2538 7282
rect 2590 6334 2668 7282
rect 2532 6322 2596 6334
rect 2662 4766 2668 6334
rect 2702 4766 2708 8742
rect 2662 4754 2708 4766
rect 2820 8742 2866 8754
rect 2820 4766 2826 8742
rect 2860 4766 2866 8742
rect 2820 4754 2866 4766
rect 2978 8742 3024 8754
rect 2978 4766 2984 8742
rect 3018 4766 3024 8742
rect 2978 4754 3024 4766
rect 3136 8742 3182 8754
rect 3136 4766 3142 8742
rect 3176 4766 3182 8742
rect 3136 4754 3182 4766
rect 3294 8742 3340 8754
rect 3294 4766 3300 8742
rect 3334 4766 3340 8742
rect 3294 4754 3340 4766
rect 3452 8742 3498 8754
rect 3452 4766 3458 8742
rect 3492 4766 3498 8742
rect 3452 4754 3498 4766
rect 3610 8742 3656 8754
rect 3610 4766 3616 8742
rect 3650 4766 3656 8742
rect 3610 4754 3656 4766
rect 3768 8742 3814 8754
rect 3768 4766 3774 8742
rect 3808 4766 3814 8742
rect 3768 4754 3814 4766
rect 3926 8742 3972 8754
rect 3926 4766 3932 8742
rect 3966 4766 3972 8742
rect 3926 4754 3972 4766
rect 4084 8742 4130 8754
rect 4084 4766 4090 8742
rect 4124 4766 4130 8742
rect 4084 4754 4130 4766
rect 4242 8742 4288 8754
rect 4242 4766 4248 8742
rect 4282 4766 4288 8742
rect 4242 4754 4288 4766
rect 4400 8742 4446 8754
rect 4400 4766 4406 8742
rect 4440 4766 4446 8742
rect 4400 4754 4446 4766
rect 4558 8742 4604 8754
rect 4558 4766 4564 8742
rect 4598 4766 4604 8742
rect 4558 4754 4604 4766
rect 4716 8742 4762 8754
rect 4716 4766 4722 8742
rect 4756 4766 4762 8742
rect 4716 4754 4762 4766
rect 4874 8742 4920 8754
rect 4874 4766 4880 8742
rect 4914 4766 4920 8742
rect 4874 4754 4920 4766
rect 5032 8742 5078 8754
rect 5032 4766 5038 8742
rect 5072 4766 5078 8742
rect 5032 4754 5078 4766
rect 5190 8742 5236 8754
rect 5190 4766 5196 8742
rect 5230 4766 5236 8742
rect 5190 4754 5236 4766
rect 5348 8742 5394 8754
rect 5348 4766 5354 8742
rect 5388 4766 5394 8742
rect 5348 4754 5394 4766
rect 5506 8742 5552 8754
rect 5506 4766 5512 8742
rect 5546 4766 5552 8742
rect 5506 4754 5552 4766
rect 5664 8742 5710 8754
rect 5664 4766 5670 8742
rect 5704 4766 5710 8742
rect 5664 4754 5710 4766
rect 5822 8742 5868 8754
rect 5822 4766 5828 8742
rect 5862 7360 5868 8742
rect 5924 7360 5988 8802
rect 5862 6412 5930 7360
rect 5982 6412 5988 7360
rect 5862 6410 5988 6412
rect 5862 4766 5868 6410
rect 5924 6400 5988 6410
rect 5822 4754 5868 4766
rect 2324 4582 2342 4682
rect 2448 4582 2464 4682
rect 2712 4600 2722 4666
rect 2788 4600 2798 4666
rect 2826 4554 2858 4754
rect 2956 4600 2966 4666
rect 3032 4600 3042 4666
rect 3142 4554 3174 4754
rect 3272 4600 3282 4666
rect 3348 4600 3358 4666
rect 3458 4554 3490 4754
rect 3588 4600 3598 4666
rect 3664 4600 3674 4666
rect 3774 4554 3806 4754
rect 3904 4600 3914 4666
rect 3980 4600 3990 4666
rect 4090 4554 4122 4754
rect 4222 4600 4232 4666
rect 4298 4600 4308 4666
rect 4406 4554 4438 4754
rect 4538 4600 4548 4666
rect 4614 4600 4624 4666
rect 4722 4554 4754 4754
rect 4852 4600 4862 4666
rect 4928 4600 4938 4666
rect 5038 4554 5070 4754
rect 5168 4600 5178 4666
rect 5244 4600 5254 4666
rect 5354 4554 5386 4754
rect 5486 4600 5496 4666
rect 5562 4600 5572 4666
rect 5670 4554 5702 4754
rect 5744 4600 5754 4666
rect 5820 4600 5830 4666
rect 2800 4548 6000 4554
rect 2800 4362 2806 4548
rect 2174 4320 2220 4332
rect 600 4264 634 4320
rect 916 4264 950 4320
rect 1232 4264 1266 4320
rect 1548 4264 1582 4320
rect 1864 4264 1898 4320
rect 2180 4264 2214 4320
rect 2798 4296 2806 4362
rect 572 4228 2606 4264
rect 2800 4240 2806 4296
rect 5994 4240 6000 4548
rect 2800 4234 6000 4240
rect 572 4162 684 4228
rect 2122 4162 2606 4228
rect 2826 4206 2858 4234
rect 3142 4206 3174 4234
rect 3458 4206 3490 4234
rect 3774 4206 3806 4234
rect 4090 4206 4122 4234
rect 4406 4206 4438 4234
rect 4722 4206 4754 4234
rect 5038 4206 5070 4234
rect 5354 4206 5386 4234
rect 5670 4206 5702 4234
rect 572 4106 2606 4162
rect 572 4092 1364 4106
rect 543 4086 1364 4092
rect 543 4040 555 4086
rect 1077 4040 1364 4086
rect 543 4034 1364 4040
rect 563 3985 597 4034
rect 755 3985 789 4034
rect 947 3985 981 4034
rect 1296 4016 1364 4034
rect 2364 4016 2606 4106
rect 1296 4010 2606 4016
rect 557 3973 603 3985
rect 557 3797 563 3973
rect 597 3797 603 3973
rect 557 3785 603 3797
rect 653 3973 699 3985
rect 653 3797 659 3973
rect 693 3797 699 3973
rect 653 3785 699 3797
rect 749 3973 795 3985
rect 749 3797 755 3973
rect 789 3797 795 3973
rect 749 3785 795 3797
rect 845 3973 891 3985
rect 845 3797 851 3973
rect 885 3797 891 3973
rect 845 3785 891 3797
rect 941 3973 987 3985
rect 941 3797 947 3973
rect 981 3797 987 3973
rect 941 3785 987 3797
rect 1037 3973 1083 3985
rect 1037 3797 1043 3973
rect 1077 3797 1083 3973
rect 1037 3785 1083 3797
rect 1296 3920 1342 4010
rect 661 3757 691 3785
rect 853 3757 883 3785
rect 641 3705 651 3757
rect 703 3705 713 3757
rect 833 3705 843 3757
rect 895 3705 905 3757
rect 1045 3756 1075 3785
rect 567 3618 625 3624
rect 567 3617 579 3618
rect 613 3617 625 3618
rect 560 3565 570 3617
rect 622 3565 632 3617
rect 661 3534 691 3705
rect 743 3618 801 3624
rect 743 3616 755 3618
rect 789 3616 801 3618
rect 736 3564 746 3616
rect 798 3564 808 3616
rect 853 3534 883 3705
rect 1024 3704 1034 3756
rect 1086 3704 1096 3756
rect 935 3615 993 3621
rect 935 3614 947 3615
rect 981 3614 993 3615
rect 929 3562 939 3614
rect 991 3562 1001 3614
rect 1045 3534 1075 3704
rect 557 3522 603 3534
rect 557 3346 563 3522
rect 597 3346 603 3522
rect 557 3334 603 3346
rect 653 3522 699 3534
rect 653 3346 659 3522
rect 693 3346 699 3522
rect 653 3334 699 3346
rect 749 3522 795 3534
rect 749 3346 755 3522
rect 789 3346 795 3522
rect 749 3334 795 3346
rect 845 3522 891 3534
rect 845 3346 851 3522
rect 885 3346 891 3522
rect 845 3334 891 3346
rect 941 3522 987 3534
rect 941 3346 947 3522
rect 981 3346 987 3522
rect 941 3334 987 3346
rect 1037 3522 1083 3534
rect 1037 3346 1043 3522
rect 1077 3346 1083 3522
rect 1037 3334 1083 3346
rect 563 3270 597 3334
rect 755 3270 789 3334
rect 947 3270 981 3334
rect 563 3268 1128 3270
rect 540 3262 1128 3268
rect 540 3226 552 3262
rect 1087 3226 1128 3262
rect 540 3220 1128 3226
rect 570 3184 1128 3220
rect 1296 3144 1302 3920
rect 1336 3144 1342 3920
rect 1296 3132 1342 3144
rect 1454 3920 1500 3932
rect 1454 3144 1460 3920
rect 1494 3144 1500 3920
rect 1454 3132 1500 3144
rect 1612 3920 1658 4010
rect 1792 3932 1824 3934
rect 1612 3144 1618 3920
rect 1652 3144 1658 3920
rect 1612 3132 1658 3144
rect 1770 3920 1824 3932
rect 1770 3144 1776 3920
rect 1810 3144 1824 3920
rect 1770 3132 1824 3144
rect 1910 3920 1956 4010
rect 1910 3144 1916 3920
rect 1950 3144 1956 3920
rect 1910 3132 1956 3144
rect 2068 3920 2114 3932
rect 2068 3144 2074 3920
rect 2108 3144 2114 3920
rect 2068 3132 2114 3144
rect 2226 3920 2272 4010
rect 2226 3144 2232 3920
rect 2266 3144 2272 3920
rect 2226 3132 2272 3144
rect 2384 3920 2430 3932
rect 2384 3144 2390 3920
rect 2424 3144 2430 3920
rect 2384 3132 2430 3144
rect 1364 3058 1374 3110
rect 1426 3058 1436 3110
rect 1364 3056 1436 3058
rect 1370 3052 1428 3056
rect 1464 2998 1494 3132
rect 1522 3058 1532 3110
rect 1584 3058 1594 3110
rect 1680 3058 1690 3110
rect 1742 3058 1752 3110
rect 1528 3054 1586 3058
rect 1688 3054 1746 3058
rect 1792 2998 1824 3132
rect 1974 3058 1984 3110
rect 2036 3058 2046 3110
rect 1982 3054 2040 3058
rect 368 2944 1824 2998
rect 2076 2956 2108 3132
rect 2136 3058 2146 3110
rect 2198 3058 2208 3110
rect 2292 3058 2302 3110
rect 2354 3058 2364 3110
rect 2144 3054 2202 3058
rect 2300 3054 2358 3058
rect 2066 2946 2108 2956
rect 0 2892 192 2904
rect 0 2832 12 2892
rect 72 2832 120 2892
rect 180 2832 192 2892
rect 1674 2864 1684 2916
rect 1736 2864 1746 2916
rect 1674 2859 1746 2864
rect 0 2822 192 2832
rect 1664 2853 1756 2859
rect 1664 2819 1676 2853
rect 1744 2819 1756 2853
rect 1664 2813 1756 2819
rect 1792 2854 1824 2944
rect 2056 2894 2066 2946
rect 2118 2936 2128 2946
rect 2392 2936 2430 3132
rect 2118 2902 2430 2936
rect 2118 2894 2128 2902
rect 2066 2882 2108 2894
rect 1954 2854 2046 2859
rect 1792 2853 2046 2854
rect 1792 2819 1966 2853
rect 2034 2819 2046 2853
rect 1792 2818 1974 2819
rect 1792 2772 1824 2818
rect 1954 2813 1974 2818
rect 1964 2792 1974 2813
rect 2026 2813 2046 2819
rect 2026 2792 2036 2813
rect 2076 2772 2108 2882
rect 1608 2760 1654 2772
rect 1608 2384 1614 2760
rect 1648 2384 1654 2760
rect 1608 2372 1654 2384
rect 1766 2760 1824 2772
rect 1766 2384 1772 2760
rect 1806 2384 1824 2760
rect 1766 2372 1824 2384
rect 1898 2760 1944 2772
rect 1898 2384 1904 2760
rect 1938 2384 1944 2760
rect 1898 2372 1944 2384
rect 2056 2760 2108 2772
rect 2056 2384 2062 2760
rect 2096 2384 2108 2760
rect 2056 2372 2108 2384
rect 2466 2746 2606 4010
rect 2662 4194 2708 4206
rect 2662 2746 2668 4194
rect 1614 2314 1648 2372
rect 1904 2314 1938 2372
rect 1614 2308 1680 2314
rect 1740 2308 1826 2314
rect 1886 2308 1980 2314
rect 2040 2308 2094 2314
rect 1614 2266 1674 2308
rect 2052 2266 2094 2308
rect 1614 2256 1680 2266
rect 1670 2254 1680 2256
rect 1740 2256 1826 2266
rect 1740 2254 1750 2256
rect 1816 2254 1826 2256
rect 1886 2256 1980 2266
rect 1886 2254 1896 2256
rect 1970 2254 1980 2256
rect 2040 2256 2094 2266
rect 2040 2254 2050 2256
rect 2466 1798 2668 2746
rect 2466 128 2606 1798
rect 2662 218 2668 1798
rect 2702 218 2708 4194
rect 2662 206 2708 218
rect 2820 4194 2866 4206
rect 2820 218 2826 4194
rect 2860 218 2866 4194
rect 2820 206 2866 218
rect 2978 4194 3024 4206
rect 2978 218 2984 4194
rect 3018 218 3024 4194
rect 2978 206 3024 218
rect 3136 4194 3182 4206
rect 3136 218 3142 4194
rect 3176 218 3182 4194
rect 3136 206 3182 218
rect 3294 4194 3340 4206
rect 3294 218 3300 4194
rect 3334 218 3340 4194
rect 3294 206 3340 218
rect 3452 4194 3498 4206
rect 3452 218 3458 4194
rect 3492 218 3498 4194
rect 3452 206 3498 218
rect 3610 4194 3656 4206
rect 3610 218 3616 4194
rect 3650 218 3656 4194
rect 3610 206 3656 218
rect 3768 4194 3814 4206
rect 3768 218 3774 4194
rect 3808 218 3814 4194
rect 3768 206 3814 218
rect 3926 4194 3972 4206
rect 3926 218 3932 4194
rect 3966 218 3972 4194
rect 3926 206 3972 218
rect 4084 4194 4130 4206
rect 4084 218 4090 4194
rect 4124 218 4130 4194
rect 4084 206 4130 218
rect 4242 4194 4288 4206
rect 4242 218 4248 4194
rect 4282 218 4288 4194
rect 4242 206 4288 218
rect 4400 4194 4446 4206
rect 4400 218 4406 4194
rect 4440 218 4446 4194
rect 4400 206 4446 218
rect 4558 4194 4604 4206
rect 4558 218 4564 4194
rect 4598 218 4604 4194
rect 4558 206 4604 218
rect 4716 4194 4762 4206
rect 4716 218 4722 4194
rect 4756 218 4762 4194
rect 4716 206 4762 218
rect 4874 4194 4920 4206
rect 4874 218 4880 4194
rect 4914 218 4920 4194
rect 4874 206 4920 218
rect 5032 4194 5078 4206
rect 5032 218 5038 4194
rect 5072 218 5078 4194
rect 5032 206 5078 218
rect 5190 4194 5236 4206
rect 5190 218 5196 4194
rect 5230 218 5236 4194
rect 5190 206 5236 218
rect 5348 4194 5394 4206
rect 5348 218 5354 4194
rect 5388 218 5394 4194
rect 5348 206 5394 218
rect 5506 4194 5552 4206
rect 5506 218 5512 4194
rect 5546 218 5552 4194
rect 5506 206 5552 218
rect 5664 4194 5710 4206
rect 5664 218 5670 4194
rect 5704 218 5710 4194
rect 5664 206 5710 218
rect 5822 4194 5868 4206
rect 5822 218 5828 4194
rect 5862 2796 5868 4194
rect 5862 1866 5988 2796
rect 5862 1848 6000 1866
rect 5862 218 5868 1848
rect 5822 206 5868 218
rect 2668 128 2702 206
rect 2982 128 3016 206
rect 3300 128 3334 206
rect 3614 128 3648 206
rect 3932 128 3966 206
rect 4246 128 4280 206
rect 4564 128 4598 206
rect 4878 128 4912 206
rect 5196 128 5230 206
rect 5510 128 5544 206
rect 5828 128 5862 206
rect 5946 128 6000 1848
rect 2466 114 6000 128
rect 2466 8 2634 114
rect 5898 8 6000 114
rect 2466 0 6000 8
<< via1 >>
rect 388 6594 488 6694
rect 668 6658 720 6668
rect 668 6624 678 6658
rect 678 6624 712 6658
rect 712 6624 720 6658
rect 668 6616 720 6624
rect 208 6372 308 6472
rect 208 3552 308 3652
rect 906 6660 958 6668
rect 906 6626 916 6660
rect 916 6626 950 6660
rect 950 6626 958 6660
rect 906 6616 958 6626
rect 1220 6660 1272 6668
rect 1220 6626 1230 6660
rect 1230 6626 1264 6660
rect 1264 6626 1272 6660
rect 1220 6616 1272 6626
rect 1538 6658 1590 6668
rect 1538 6624 1548 6658
rect 1548 6624 1582 6658
rect 1582 6624 1590 6658
rect 1538 6616 1590 6624
rect 1852 6658 1904 6668
rect 1852 6624 1862 6658
rect 1862 6624 1896 6658
rect 1896 6624 1904 6658
rect 1852 6616 1904 6624
rect 2096 6658 2148 6668
rect 2096 6624 2106 6658
rect 2106 6624 2140 6658
rect 2140 6624 2148 6658
rect 2096 6616 2148 6624
rect 748 6506 800 6558
rect 1064 6506 1116 6558
rect 1382 6506 1434 6558
rect 1698 6506 1750 6558
rect 2014 6506 2066 6558
rect 668 6440 720 6450
rect 668 6406 678 6440
rect 678 6406 712 6440
rect 712 6406 720 6440
rect 668 6398 720 6406
rect 906 6442 958 6450
rect 906 6408 916 6442
rect 916 6408 950 6442
rect 950 6408 958 6442
rect 906 6398 958 6408
rect 1220 6442 1272 6450
rect 1220 6408 1230 6442
rect 1230 6408 1264 6442
rect 1264 6408 1272 6442
rect 1220 6398 1272 6408
rect 1538 6440 1590 6450
rect 1538 6406 1548 6440
rect 1548 6406 1582 6440
rect 1582 6406 1590 6440
rect 1538 6398 1590 6406
rect 1852 6440 1904 6450
rect 1852 6406 1862 6440
rect 1862 6406 1896 6440
rect 1896 6406 1904 6440
rect 1852 6398 1904 6406
rect 2340 6486 2446 6586
rect 2096 6440 2148 6450
rect 2096 6406 2106 6440
rect 2106 6406 2140 6440
rect 2140 6406 2148 6440
rect 2096 6398 2148 6406
rect 2342 4582 2448 4682
rect 2722 4650 2788 4666
rect 2722 4616 2738 4650
rect 2738 4616 2772 4650
rect 2772 4616 2788 4650
rect 2722 4600 2788 4616
rect 2966 4650 3032 4666
rect 2966 4616 2982 4650
rect 2982 4616 3016 4650
rect 3016 4616 3032 4650
rect 2966 4600 3032 4616
rect 3282 4650 3348 4666
rect 3282 4616 3298 4650
rect 3298 4616 3332 4650
rect 3332 4616 3348 4650
rect 3282 4600 3348 4616
rect 3598 4650 3664 4666
rect 3598 4616 3614 4650
rect 3614 4616 3648 4650
rect 3648 4616 3664 4650
rect 3598 4600 3664 4616
rect 3914 4650 3980 4666
rect 3914 4616 3930 4650
rect 3930 4616 3964 4650
rect 3964 4616 3980 4650
rect 3914 4600 3980 4616
rect 4232 4650 4298 4666
rect 4232 4616 4248 4650
rect 4248 4616 4282 4650
rect 4282 4616 4298 4650
rect 4232 4600 4298 4616
rect 4548 4650 4614 4666
rect 4548 4616 4564 4650
rect 4564 4616 4598 4650
rect 4598 4616 4614 4650
rect 4548 4600 4614 4616
rect 4862 4650 4928 4666
rect 4862 4616 4878 4650
rect 4878 4616 4912 4650
rect 4912 4616 4928 4650
rect 4862 4600 4928 4616
rect 5178 4650 5244 4666
rect 5178 4616 5194 4650
rect 5194 4616 5228 4650
rect 5228 4616 5244 4650
rect 5178 4600 5244 4616
rect 5496 4650 5562 4666
rect 5496 4616 5512 4650
rect 5512 4616 5546 4650
rect 5546 4616 5562 4650
rect 5496 4600 5562 4616
rect 5754 4650 5820 4666
rect 5754 4616 5770 4650
rect 5770 4616 5804 4650
rect 5804 4616 5820 4650
rect 5754 4600 5820 4616
rect 2806 4240 5994 4548
rect 651 3705 703 3757
rect 843 3705 895 3757
rect 570 3584 579 3617
rect 579 3584 613 3617
rect 613 3584 622 3617
rect 570 3565 622 3584
rect 746 3584 755 3616
rect 755 3584 789 3616
rect 789 3584 798 3616
rect 746 3564 798 3584
rect 1034 3704 1086 3756
rect 939 3581 947 3614
rect 947 3581 981 3614
rect 981 3581 991 3614
rect 939 3562 991 3581
rect 1374 3092 1426 3110
rect 1374 3058 1382 3092
rect 1382 3058 1416 3092
rect 1416 3058 1426 3092
rect 1532 3094 1584 3110
rect 1532 3060 1540 3094
rect 1540 3060 1574 3094
rect 1574 3060 1584 3094
rect 1532 3058 1584 3060
rect 1690 3094 1742 3110
rect 1690 3060 1700 3094
rect 1700 3060 1734 3094
rect 1734 3060 1742 3094
rect 1690 3058 1742 3060
rect 1984 3094 2036 3110
rect 1984 3060 1994 3094
rect 1994 3060 2028 3094
rect 2028 3060 2036 3094
rect 1984 3058 2036 3060
rect 2146 3094 2198 3110
rect 2146 3060 2156 3094
rect 2156 3060 2190 3094
rect 2190 3060 2198 3094
rect 2146 3058 2198 3060
rect 2302 3094 2354 3110
rect 2302 3060 2312 3094
rect 2312 3060 2346 3094
rect 2346 3060 2354 3094
rect 2302 3058 2354 3060
rect 12 2832 72 2892
rect 120 2832 180 2892
rect 1684 2864 1736 2916
rect 2066 2894 2118 2946
rect 1974 2819 2026 2844
rect 1974 2792 2026 2819
rect 1680 2308 1740 2314
rect 1826 2308 1886 2314
rect 1980 2308 2040 2314
rect 1680 2266 1740 2308
rect 1826 2266 1886 2308
rect 1980 2266 2040 2308
rect 1680 2254 1740 2266
rect 1826 2254 1886 2266
rect 1980 2254 2040 2266
<< metal2 >>
rect 388 6694 488 6704
rect 488 6668 2290 6682
rect 488 6616 668 6668
rect 720 6616 906 6668
rect 958 6616 1220 6668
rect 1272 6616 1538 6668
rect 1590 6616 1852 6668
rect 1904 6616 2096 6668
rect 2148 6616 2290 6668
rect 488 6604 2290 6616
rect 668 6602 2290 6604
rect 388 6584 488 6594
rect 2340 6586 2446 6596
rect 518 6558 2340 6572
rect 518 6506 748 6558
rect 800 6506 1064 6558
rect 1116 6506 1382 6558
rect 1434 6506 1698 6558
rect 1750 6506 2014 6558
rect 2066 6506 2340 6558
rect 518 6492 2340 6506
rect 208 6472 308 6482
rect 2340 6476 2446 6486
rect 204 6384 208 6462
rect 308 6450 2290 6462
rect 308 6398 668 6450
rect 720 6398 906 6450
rect 958 6398 1220 6450
rect 1272 6398 1538 6450
rect 1590 6398 1852 6450
rect 1904 6398 2096 6450
rect 2148 6398 2290 6450
rect 308 6384 2290 6398
rect 208 6362 308 6372
rect 2342 4682 2448 4692
rect 2448 4666 5906 4682
rect 2448 4600 2722 4666
rect 2788 4600 2966 4666
rect 3032 4600 3282 4666
rect 3348 4600 3598 4666
rect 3664 4600 3914 4666
rect 3980 4600 4232 4666
rect 4298 4600 4548 4666
rect 4614 4600 4862 4666
rect 4928 4600 5178 4666
rect 5244 4600 5496 4666
rect 5562 4600 5754 4666
rect 5820 4600 5906 4666
rect 2448 4582 5906 4600
rect 2342 4572 2448 4582
rect 2800 4548 6000 4554
rect 2800 4378 2806 4548
rect 2616 4278 2806 4378
rect 2800 4240 2806 4278
rect 5994 4240 6000 4548
rect 2800 4234 6000 4240
rect 651 3758 703 3767
rect 843 3758 895 3767
rect 1034 3758 1086 3766
rect 549 3757 1286 3758
rect 549 3744 651 3757
rect 514 3716 651 3744
rect 549 3705 651 3716
rect 703 3705 843 3757
rect 895 3756 1286 3757
rect 895 3705 1034 3756
rect 651 3695 703 3705
rect 843 3695 895 3705
rect 1086 3705 1286 3756
rect 1034 3694 1086 3704
rect 208 3652 308 3658
rect 308 3617 1194 3628
rect 308 3568 570 3617
rect 622 3616 1194 3617
rect 622 3568 746 3616
rect 570 3555 622 3565
rect 798 3614 1194 3616
rect 798 3568 939 3614
rect 746 3554 798 3564
rect 991 3568 1194 3614
rect 939 3552 991 3562
rect 208 3538 308 3552
rect 1134 3020 1194 3568
rect 1226 3102 1286 3705
rect 1374 3110 1426 3120
rect 1226 3068 1374 3102
rect 1532 3110 1584 3120
rect 1426 3068 1532 3102
rect 1374 3048 1426 3058
rect 1690 3110 1742 3120
rect 1584 3068 1690 3102
rect 1532 3048 1584 3058
rect 1984 3110 2036 3120
rect 1742 3068 1752 3102
rect 1690 3048 1742 3058
rect 1984 3020 2036 3058
rect 2146 3110 2198 3120
rect 2146 3020 2198 3058
rect 2302 3110 2354 3120
rect 2302 3020 2354 3058
rect 1134 2986 2354 3020
rect 2066 2946 2118 2956
rect 1684 2916 2066 2936
rect 0 2892 192 2904
rect 0 2832 12 2892
rect 72 2832 120 2892
rect 180 2832 1540 2892
rect 1736 2902 2066 2916
rect 2066 2882 2118 2894
rect 1684 2854 1736 2864
rect 0 2822 192 2832
rect 1498 2312 1540 2832
rect 1950 2844 2174 2854
rect 1950 2820 1974 2844
rect 2026 2820 2174 2844
rect 1974 2760 2026 2792
rect 1680 2314 1740 2324
rect 1498 2254 1680 2312
rect 1826 2314 1886 2324
rect 1740 2254 1826 2312
rect 1980 2314 2040 2324
rect 1886 2254 1980 2312
rect 2040 2254 2124 2312
rect 1518 2252 2124 2254
rect 1680 2244 1740 2252
rect 1826 2244 1886 2252
rect 1980 2244 2040 2252
<< via2 >>
rect 2809 4243 5991 4545
<< metal3 >>
rect 2800 4548 6000 4554
rect 2800 4240 2806 4548
rect 5994 4240 6000 4548
rect 2800 4234 6000 4240
<< via3 >>
rect 2806 4545 5994 4548
rect 2806 4243 2809 4545
rect 2809 4243 5991 4545
rect 5991 4243 5994 4545
rect 2806 4240 5994 4243
<< metal4 >>
rect 2800 4548 6000 4554
rect 2800 4240 2806 4548
rect 5994 4240 6000 4548
rect 2800 4234 6000 4240
<< via4 >>
rect 2824 4258 5976 4530
<< metal5 >>
rect 2800 4530 6000 4554
rect 2800 4258 2824 4530
rect 5976 4258 6000 4530
rect 2800 4234 6000 4258
<< labels >>
rlabel metal1 570 3184 1128 3270 1 level_shifter_0/VDD
rlabel metal1 576 8806 5720 8896 1 level_shifter_0/VH
rlabel metal1 190 3648 330 6372 1 level_shifter_0/IN
rlabel metal1 2466 0 2606 4264 1 level_shifter_0/GND
rlabel space 2588 0 5942 8930 1 level_shifter_0/OUT
rlabel metal1 576 8864 2238 8870 1 level_shifter_0/stage_100_0/VH
rlabel metal2 2066 6492 2288 6572 1 level_shifter_0/stage_100_0/OUT
rlabel metal1 600 4154 2214 4160 1 level_shifter_0/stage_100_0/GND
rlabel space 520 6602 668 6682 1 level_shifter_0/stage_100_0/A
rlabel metal2 520 6384 668 6462 1 level_shifter_0/stage_100_0/B
rlabel metal2 2616 4582 2722 4682 1 level_shifter_0/inv_400_0/IN
rlabel metal1 543 4086 1089 4092 5 level_shifter_0/inv_1_8_0/GND
rlabel metal2 1086 3716 1125 3744 5 level_shifter_0/inv_1_8_0/OUT
rlabel metal2 515 3576 570 3604 5 level_shifter_0/inv_1_8_0/IN
rlabel metal1 540 3220 1099 3226 5 level_shifter_0/inv_1_8_0/VDD
rlabel metal2 2026 2820 2174 2854 5 level_shifter_0/cruzados_0/OUT
rlabel metal1 1614 2256 2094 2262 5 level_shifter_0/cruzados_0/VH
rlabel metal2 1290 3068 1374 3102 5 level_shifter_0/cruzados_0/IN1
rlabel metal2 1540 2986 1976 3020 5 level_shifter_0/cruzados_0/IN2
rlabel via2 5720 4278 5906 4378 1 level_shifter_0/OUT
rlabel via2 5720 4278 5906 4378 1 level_shifter_0/inv_400_0/OUT
<< end >>
