# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.380000 BY  4.590000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT 0.000000 0.000000 1.915000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 0.750000 ;
        RECT 0.000000 0.750000 1.915000 0.890000 ;
        RECT 0.000000 0.890000 0.330000 1.310000 ;
        RECT 0.000000 1.310000 1.915000 1.450000 ;
        RECT 0.000000 1.450000 0.330000 1.870000 ;
        RECT 0.000000 1.870000 1.915000 2.010000 ;
        RECT 0.000000 2.010000 0.330000 2.020000 ;
        RECT 0.000000 2.570000 0.330000 2.580000 ;
        RECT 0.000000 2.580000 1.915000 2.720000 ;
        RECT 0.000000 2.720000 0.330000 3.140000 ;
        RECT 0.000000 3.140000 1.915000 3.280000 ;
        RECT 0.000000 3.280000 0.330000 3.700000 ;
        RECT 0.000000 3.700000 1.915000 3.840000 ;
        RECT 0.000000 3.840000 0.330000 4.260000 ;
        RECT 0.000000 4.260000 1.915000 4.590000 ;
        RECT 2.465000 0.000000 4.380000 0.330000 ;
        RECT 2.465000 0.750000 4.380000 0.890000 ;
        RECT 2.465000 1.310000 4.380000 1.450000 ;
        RECT 2.465000 1.870000 4.380000 2.010000 ;
        RECT 2.465000 2.580000 4.380000 2.720000 ;
        RECT 2.465000 3.140000 4.380000 3.280000 ;
        RECT 2.465000 3.700000 4.380000 3.840000 ;
        RECT 2.465000 4.260000 4.380000 4.590000 ;
        RECT 4.050000 0.330000 4.380000 0.750000 ;
        RECT 4.050000 0.890000 4.380000 1.310000 ;
        RECT 4.050000 1.450000 4.380000 1.870000 ;
        RECT 4.050000 2.010000 4.380000 2.020000 ;
        RECT 4.050000 2.570000 4.380000 2.580000 ;
        RECT 4.050000 2.720000 4.380000 3.140000 ;
        RECT 4.050000 3.280000 4.380000 3.700000 ;
        RECT 4.050000 3.840000 4.380000 4.260000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT 0.000000 2.160000 4.380000 2.430000 ;
        RECT 0.470000 0.470000 3.910000 0.610000 ;
        RECT 0.470000 1.030000 3.910000 1.170000 ;
        RECT 0.470000 1.590000 3.910000 1.730000 ;
        RECT 0.470000 2.860000 3.910000 3.000000 ;
        RECT 0.470000 3.420000 3.910000 3.560000 ;
        RECT 0.470000 3.980000 3.910000 4.120000 ;
        RECT 2.055000 0.000000 2.325000 0.470000 ;
        RECT 2.055000 0.610000 2.325000 1.030000 ;
        RECT 2.055000 1.170000 2.325000 1.590000 ;
        RECT 2.055000 1.730000 2.325000 2.160000 ;
        RECT 2.055000 2.430000 2.325000 2.860000 ;
        RECT 2.055000 3.000000 2.325000 3.420000 ;
        RECT 2.055000 3.560000 2.325000 3.980000 ;
        RECT 2.055000 4.120000 2.325000 4.590000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 2.335000 1.750000 2.455000 2.005000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 4.380000 4.590000 ;
    LAYER mcon ;
      RECT 0.080000 0.410000 0.250000 0.580000 ;
      RECT 0.080000 0.770000 0.250000 0.940000 ;
      RECT 0.080000 1.130000 0.250000 1.300000 ;
      RECT 0.080000 1.490000 0.250000 1.660000 ;
      RECT 0.080000 1.850000 0.250000 2.020000 ;
      RECT 0.080000 2.210000 0.250000 2.380000 ;
      RECT 0.080000 2.570000 0.250000 2.740000 ;
      RECT 0.080000 2.930000 0.250000 3.100000 ;
      RECT 0.080000 3.290000 0.250000 3.460000 ;
      RECT 0.080000 3.650000 0.250000 3.820000 ;
      RECT 0.080000 4.010000 0.250000 4.180000 ;
      RECT 0.485000 0.080000 0.655000 0.250000 ;
      RECT 0.485000 4.340000 0.655000 4.510000 ;
      RECT 0.845000 0.080000 1.015000 0.250000 ;
      RECT 0.845000 4.340000 1.015000 4.510000 ;
      RECT 1.205000 0.080000 1.375000 0.250000 ;
      RECT 1.205000 4.340000 1.375000 4.510000 ;
      RECT 1.565000 0.080000 1.735000 0.250000 ;
      RECT 1.565000 4.340000 1.735000 4.510000 ;
      RECT 1.925000 0.080000 2.095000 0.250000 ;
      RECT 1.925000 4.340000 2.095000 4.510000 ;
      RECT 2.285000 0.080000 2.455000 0.250000 ;
      RECT 2.285000 4.340000 2.455000 4.510000 ;
      RECT 2.645000 0.080000 2.815000 0.250000 ;
      RECT 2.645000 4.340000 2.815000 4.510000 ;
      RECT 3.005000 0.080000 3.175000 0.250000 ;
      RECT 3.005000 4.340000 3.175000 4.510000 ;
      RECT 3.365000 0.080000 3.535000 0.250000 ;
      RECT 3.365000 4.340000 3.535000 4.510000 ;
      RECT 3.725000 0.080000 3.895000 0.250000 ;
      RECT 3.725000 4.340000 3.895000 4.510000 ;
      RECT 4.130000 0.410000 4.300000 0.580000 ;
      RECT 4.130000 0.770000 4.300000 0.940000 ;
      RECT 4.130000 1.130000 4.300000 1.300000 ;
      RECT 4.130000 1.490000 4.300000 1.660000 ;
      RECT 4.130000 1.850000 4.300000 2.020000 ;
      RECT 4.130000 2.210000 4.300000 2.380000 ;
      RECT 4.130000 2.570000 4.300000 2.740000 ;
      RECT 4.130000 2.930000 4.300000 3.100000 ;
      RECT 4.130000 3.290000 4.300000 3.460000 ;
      RECT 4.130000 3.650000 4.300000 3.820000 ;
      RECT 4.130000 4.010000 4.300000 4.180000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 4.380000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 4.260000 ;
      RECT 0.000000 4.260000 4.380000 4.590000 ;
      RECT 0.565000 0.470000 0.705000 2.135000 ;
      RECT 0.565000 2.135000 3.815000 2.455000 ;
      RECT 0.565000 2.455000 0.705000 4.120000 ;
      RECT 0.845000 0.330000 0.985000 1.995000 ;
      RECT 0.845000 2.595000 0.985000 4.260000 ;
      RECT 1.125000 0.470000 1.265000 2.135000 ;
      RECT 1.125000 2.455000 1.265000 4.120000 ;
      RECT 1.405000 0.330000 1.545000 1.995000 ;
      RECT 1.405000 2.595000 1.545000 4.260000 ;
      RECT 1.685000 0.470000 1.825000 2.135000 ;
      RECT 1.685000 2.455000 1.825000 4.120000 ;
      RECT 2.055000 0.470000 2.325000 2.135000 ;
      RECT 2.055000 2.455000 2.325000 4.120000 ;
      RECT 2.555000 0.470000 2.695000 2.135000 ;
      RECT 2.555000 2.455000 2.695000 4.120000 ;
      RECT 2.835000 0.330000 2.975000 1.995000 ;
      RECT 2.835000 2.595000 2.975000 4.260000 ;
      RECT 3.115000 0.470000 3.255000 2.135000 ;
      RECT 3.115000 2.455000 3.255000 4.120000 ;
      RECT 3.395000 0.330000 3.535000 1.995000 ;
      RECT 3.395000 2.595000 3.535000 4.260000 ;
      RECT 3.675000 0.470000 3.815000 2.135000 ;
      RECT 3.675000 2.455000 3.815000 4.120000 ;
      RECT 4.050000 0.330000 4.380000 4.260000 ;
    LAYER via ;
      RECT 0.035000 0.380000 0.295000 0.640000 ;
      RECT 0.035000 0.700000 0.295000 0.960000 ;
      RECT 0.035000 1.020000 0.295000 1.280000 ;
      RECT 0.035000 1.340000 0.295000 1.600000 ;
      RECT 0.035000 1.660000 0.295000 1.920000 ;
      RECT 0.035000 2.670000 0.295000 2.930000 ;
      RECT 0.035000 2.990000 0.295000 3.250000 ;
      RECT 0.035000 3.310000 0.295000 3.570000 ;
      RECT 0.035000 3.630000 0.295000 3.890000 ;
      RECT 0.035000 3.950000 0.295000 4.210000 ;
      RECT 0.260000 0.035000 0.520000 0.295000 ;
      RECT 0.260000 4.295000 0.520000 4.555000 ;
      RECT 0.580000 0.035000 0.840000 0.295000 ;
      RECT 0.580000 4.295000 0.840000 4.555000 ;
      RECT 0.595000 2.165000 0.855000 2.425000 ;
      RECT 0.900000 0.035000 1.160000 0.295000 ;
      RECT 0.900000 4.295000 1.160000 4.555000 ;
      RECT 0.915000 2.165000 1.175000 2.425000 ;
      RECT 1.220000 0.035000 1.480000 0.295000 ;
      RECT 1.220000 4.295000 1.480000 4.555000 ;
      RECT 1.235000 2.165000 1.495000 2.425000 ;
      RECT 1.540000 0.035000 1.800000 0.295000 ;
      RECT 1.540000 4.295000 1.800000 4.555000 ;
      RECT 1.555000 2.165000 1.815000 2.425000 ;
      RECT 2.060000 0.500000 2.320000 0.760000 ;
      RECT 2.060000 0.820000 2.320000 1.080000 ;
      RECT 2.060000 1.140000 2.320000 1.400000 ;
      RECT 2.060000 1.460000 2.320000 1.720000 ;
      RECT 2.060000 1.780000 2.320000 2.040000 ;
      RECT 2.060000 2.550000 2.320000 2.810000 ;
      RECT 2.060000 2.870000 2.320000 3.130000 ;
      RECT 2.060000 3.190000 2.320000 3.450000 ;
      RECT 2.060000 3.510000 2.320000 3.770000 ;
      RECT 2.060000 3.830000 2.320000 4.090000 ;
      RECT 2.565000 2.165000 2.825000 2.425000 ;
      RECT 2.580000 0.035000 2.840000 0.295000 ;
      RECT 2.580000 4.295000 2.840000 4.555000 ;
      RECT 2.885000 2.165000 3.145000 2.425000 ;
      RECT 2.900000 0.035000 3.160000 0.295000 ;
      RECT 2.900000 4.295000 3.160000 4.555000 ;
      RECT 3.205000 2.165000 3.465000 2.425000 ;
      RECT 3.220000 0.035000 3.480000 0.295000 ;
      RECT 3.220000 4.295000 3.480000 4.555000 ;
      RECT 3.525000 2.165000 3.785000 2.425000 ;
      RECT 3.540000 0.035000 3.800000 0.295000 ;
      RECT 3.540000 4.295000 3.800000 4.555000 ;
      RECT 3.860000 0.035000 4.120000 0.295000 ;
      RECT 3.860000 4.295000 4.120000 4.555000 ;
      RECT 4.085000 0.380000 4.345000 0.640000 ;
      RECT 4.085000 0.700000 4.345000 0.960000 ;
      RECT 4.085000 1.020000 4.345000 1.280000 ;
      RECT 4.085000 1.340000 4.345000 1.600000 ;
      RECT 4.085000 1.660000 4.345000 1.920000 ;
      RECT 4.085000 2.670000 4.345000 2.930000 ;
      RECT 4.085000 2.990000 4.345000 3.250000 ;
      RECT 4.085000 3.310000 4.345000 3.570000 ;
      RECT 4.085000 3.630000 4.345000 3.890000 ;
      RECT 4.085000 3.950000 4.345000 4.210000 ;
  END
END sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1
END LIBRARY
