* NGSPICE file created from Unnamed_e9e9e382.ext - technology: sky130A

.subckt ota AVSS AVDD INM INP VOUT NBC_10U NB_10U
X0 AVDD a_n14196_2392# a_n14196_2392# AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=49.1712 ps=283.36 w=1.88 l=3 M=4
X2 a_7567_n7591# a_7567_n7591# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X3 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=102.063 ps=586.58 w=4 l=2 M=23.235
X4 VOUT a_n793_n4248# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1 M=2
X5 a_7567_n7591# NB_10U a_4567_n7591# AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X6 a_n793_n4248# a_n3478_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X7 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=0 ps=0 w=3 l=4 M=4
X8 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0 ps=0 w=0.5 l=4 M=4
X9 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=1 M=5.63636
X10 a_4567_n7591# NBC_10U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X11 a_n8111_n7591# NB_10U a_n14196_2392# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X12 NBC_10U NB_10U a_n2123_n7595# AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X13 a_n7071_n377# INM a_n14274_2810# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X14 AVSS NBC_10U a_n2123_n7595# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X15 AVSS NBC_10U a_n8111_n7591# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X16 a_n3478_1981# a_n2600_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X17 a_n2600_1981# AVSS a_n3478_1981# AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=4
X18 a_n511_n10433# NB_10U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=2
X19 a_n2600_1981# AVDD a_n3478_1981# AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0.195 ps=1.78 w=0.5 l=4
X20 a_4636_n502# a_7567_n7591# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X21 VOUT a_n331_9295# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X22 a_n511_n10433# NB_10U NB_10U AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X23 AVSS a_n14274_2810# a_n7071_n377# AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=1.0725 ps=6.28 w=2.75 l=1
X24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1 M=4
X25 a_n331_9295# a_n2600_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X26 AVDD a_n14196_2392# a_n14274_2810# AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X27 a_n331_9295# AVSS a_n2600_1981# AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=4
X28 a_n331_9295# INP a_n7071_n377# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X29 a_n331_9295# AVDD a_n2600_1981# AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0.195 ps=1.78 w=0.5 l=4
X30 a_n1678_n502# a_4636_n502# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=1.0725 ps=6.28 w=2.75 l=1
X31 a_n793_n4248# a_n793_n4248# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1 M=2
X32 a_n3478_1981# INM a_n1678_n502# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X33 a_4636_n502# INP a_n1678_n502# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
C0 VOUT a_7567_n7591# 0.030081f
C1 AVDD a_n7071_n377# 0.312363f
C2 a_n2123_n7595# NBC_10U 1.86424f
C3 a_4636_n502# a_n7071_n377# 0.01349f
C4 a_n7071_n377# a_n3478_1981# 0.154388f
C5 VOUT INP 0.624677f
C6 a_n7071_n377# a_n14274_2810# 0.770148f
C7 a_n8111_n7591# NBC_10U 0.688699f
C8 a_4567_n7591# a_7567_n7591# 0.908378f
C9 VOUT INM 1.70571f
C10 a_n1678_n502# a_n331_9295# 0.145287f
C11 NB_10U NBC_10U 4.04866f
C12 a_n14196_2392# a_n793_n4248# 0.030081f
C13 a_n14196_2392# a_n8111_n7591# 0.905992f
C14 AVDD a_n14196_2392# 13.6909f
C15 AVDD a_n1678_n502# 0.002776f
C16 INP a_n331_9295# 0.33566f
C17 a_4636_n502# a_n1678_n502# 0.77567f
C18 a_n14196_2392# a_n14274_2810# 0.81726f
C19 AVDD a_7567_n7591# 13.691f
C20 a_n14196_2392# NB_10U 0.68562f
C21 a_n1678_n502# a_n3478_1981# 0.702961f
C22 a_n2600_1981# a_n331_9295# 2.40293f
C23 a_4636_n502# a_7567_n7591# 0.81726f
C24 a_n1678_n502# a_n14274_2810# 0.014407f
C25 AVDD INP 1.02e-19
C26 a_7567_n7591# NB_10U 0.693f
C27 a_n7071_n377# a_n1678_n502# 0.673655f
C28 a_4636_n502# INP 1.00579f
C29 AVDD a_n2600_1981# 11.861799f
C30 a_n2600_1981# a_n3478_1981# 2.43658f
C31 INM a_n793_n4248# 0.402672f
C32 VOUT a_n331_9295# 0.546473f
C33 a_n7071_n377# INP 0.454012f
C34 AVDD INM 1.02e-19
C35 a_n7071_n377# a_n2600_1981# 1.51e-19
C36 VOUT a_n793_n4248# 1.67238f
C37 INM a_n3478_1981# 0.318063f
C38 VOUT AVDD 6.07543f
C39 INM a_n14274_2810# 1.01091f
C40 a_7567_n7591# NBC_10U 0.2407f
C41 a_4636_n502# VOUT 0.412229f
C42 VOUT a_n3478_1981# 0.019931f
C43 a_n7071_n377# INM 0.443361f
C44 VOUT a_n14274_2810# 0.042473f
C45 a_n511_n10433# NB_10U 2.43324f
C46 a_n2123_n7595# a_n793_n4248# 5.78e-19
C47 a_n793_n4248# a_n331_9295# 0.008459f
C48 a_4567_n7591# NB_10U 0.884825f
C49 a_n1678_n502# INP 0.444433f
C50 AVDD a_n331_9295# 10.589099f
C51 a_7567_n7591# INP 0.111898f
C52 a_4636_n502# a_n331_9295# 0.003411f
C53 a_n2123_n7595# NB_10U 0.884326f
C54 a_n1678_n502# a_n2600_1981# 5.52e-20
C55 a_n3478_1981# a_n331_9295# 0.926096f
C56 a_n511_n10433# NBC_10U 0.225304f
C57 AVDD a_n793_n4248# 6.57186f
C58 a_n14196_2392# INM 0.111898f
C59 a_n793_n4248# a_n3478_1981# 0.579778f
C60 a_n1678_n502# INM 0.472144f
C61 a_n7071_n377# a_n331_9295# 0.753404f
C62 a_4636_n502# AVDD 5.27562f
C63 a_n793_n4248# a_n14274_2810# 0.328962f
C64 AVDD a_n3478_1981# 11.1099f
C65 VOUT a_n14196_2392# 0.3024f
C66 a_n8111_n7591# NB_10U 0.884326f
C67 AVDD a_n14274_2810# 5.27646f
C68 a_4567_n7591# NBC_10U 0.886164f
C69 VOUT a_n1678_n502# 3.66e-19
C70 a_n14274_2810# a_n3478_1981# 0.002492f
C71 NBC_10U AVSS 30.1985f
C72 NB_10U AVSS 30.492498f
C73 INP AVSS 11.368901f
C74 INM AVSS 10.2179f
C75 VOUT AVSS 31.356201f
C76 AVDD AVSS 0.198435p
C77 a_n511_n10433# AVSS 3.93212f
C78 a_4567_n7591# AVSS 3.97159f
C79 a_n2123_n7595# AVSS 4.51136f
C80 a_n8111_n7591# AVSS 4.02475f
C81 a_n1678_n502# AVSS 8.590281f
C82 a_n7071_n377# AVSS 8.062799f
C83 a_4636_n502# AVSS 10.5205f
C84 a_7567_n7591# AVSS 8.656019f
C85 a_n14274_2810# AVSS 10.512199f
C86 a_n14196_2392# AVSS 8.488259f
C87 a_n2600_1981# AVSS 5.51582f
C88 a_n793_n4248# AVSS 26.0236f
C89 a_n331_9295# AVSS 7.30627f
C90 a_n3478_1981# AVSS 7.09573f
.ends

