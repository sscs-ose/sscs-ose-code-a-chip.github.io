.param VDD=1.8 VG=1.397 VCM=1.097 I_B=50u vi=0.6 fi=10000000 WMB=22 LMB=0.5 WM4=22 LM4=0.5 WM1=7 LM1=0.5 WM3=14 LM3=0.5 RL=2k I_CM=250u
