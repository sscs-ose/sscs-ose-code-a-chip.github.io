.param w1_2=$W1-2
.param w3_4=$W3-4
.param w5_6=$W5-6
.param w7_8=$W7-8
.param w9_10=$W9-10
.param beta=1
.param nf1_2=1
.param nf3_4=1
.param nf5_6=1
.param nf7_8=1
.param nf9_10=1

.param iref_ideal=65u
.param iref_post_layout=70u
