** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/tb_cm_ota_working_v2_extracted_ac.sch
**.subckt tb_cm_ota_working_v2_extracted_ac
V1 vdd GND 1.8
C1 out GND 500f m=1
V3 inn GND DC 1
V4 inp GND DC 1 AC 1
X1 vdd out inp inn itail GND cm_ota
I3 itail GND 73.87u
**** begin user architecture code

** opencircuitdesign pdks isntsall
.lib /opt/pdk/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.temp 27
.option savecurrents
.save all
.control
	ac dec 100 1 1e15
	plot vdb(out) vs frequency
	plot (180*cph(out)/pi) vs frequency
.endc


**** end user architecture code
**.ends

* expanding   symbol:  cm_ota.sym # of pins=6
** sym_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sym
** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sch
.subckt cm_ota vdd out inp inn itail vss
X0 AVSS li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 AVSS li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 AVSS li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3 AVSS li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 li_4275_2335# li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 AVSS li_4275_2335# li_4275_2335# AVSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 li_4275_2335# li_4275_2335# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7 AVSS li_4275_2335# li_4275_2335# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 m1_914_2324# INP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.235 pd=2.8 as=7.22 ps=86.4 w=0.42 l=0.15
X9 AVSS INP m1_914_2324# AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10 m1_914_2324# INP AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11 AVSS INP m1_914_2324# AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12 m1_7138_2408# INN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.235 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X13 AVSS INN m1_7138_2408# AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X14 m1_7138_2408# INN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X15 AVSS INN m1_7138_2408# AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X16 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X25 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X27 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X31 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X40 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X41 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X42 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X43 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X44 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X45 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X46 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X48 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X49 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X50 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X51 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X52 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X54 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X55 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X56 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X57 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X58 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X59 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X60 m1_4042_560# m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X61 AVSS m1_4042_560# m1_4042_560# AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X62 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X63 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X64 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X65 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X66 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X67 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X68 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X69 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X70 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X71 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X72 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X73 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X75 AVDD_1V8 m1_914_2324# OUT AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X76 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X77 OUT m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X78 m1_914_2324# m1_914_2324# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X79 AVDD_1V8 m1_914_2324# m1_914_2324# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X80 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=2.54 pd=30.6 as=0.941 ps=11.2 w=0.42 l=0.15
X81 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X82 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X83 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X84 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X85 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X86 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X87 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X88 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X89 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X90 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X91 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X92 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X93 AVDD_1V8 m1_7138_2408# m1_4042_560# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X94 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X95 m1_4042_560# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X96 m1_7138_2408# m1_7138_2408# AVDD_1V8 AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X97 AVDD_1V8 m1_7138_2408# m1_7138_2408# AVDD_1V8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X98 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X99 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X100 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X101 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X102 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X103 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X104 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X105 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X106 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X107 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X108 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X109 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X110 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X112 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X113 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X114 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X115 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X116 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X117 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X118 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X119 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X120 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X121 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X122 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X123 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X124 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X125 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X126 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X127 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X128 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X129 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X130 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X131 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X132 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X133 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X134 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X135 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X136 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X137 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X139 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X140 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X141 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X142 OUT m1_4042_560# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X143 AVSS m1_4042_560# OUT AVSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 m1_914_2324# m1_4042_560# 0.0195f
C1 OUT m1_914_2324# 1.1f
C2 INP m1_4042_560# 0.00381f
C3 li_4275_2335# m1_7138_2408# 1.51e-19
C4 AVDD_1V8 m1_7138_2408# 7.73f
C5 li_4275_2335# AVDD_1V8 0.0109f
C6 INN m1_7138_2408# 0.254f
C7 li_4275_2335# INN 0.0413f
C8 AVDD_1V8 INN 0.0333f
C9 OUT INP 8.6e-19
C10 li_4275_2335# m1_914_2324# 0.00535f
C11 m1_914_2324# AVDD_1V8 7.68f
C12 OUT m1_4042_560# 2.34f
C13 li_4275_2335# INP 0.0442f
C14 INP AVDD_1V8 0.033f
C15 m1_4042_560# m1_7138_2408# 1.11f
C16 li_4275_2335# m1_4042_560# 0.0091f
C17 m1_4042_560# AVDD_1V8 8.37f
C18 m1_4042_560# INN 0.00467f
C19 m1_914_2324# INP 0.254f
C20 li_4275_2335# OUT 0.0189f
C21 OUT AVDD_1V8 6.79f
C22 OUT AVSS 18.5f
C23 m1_4042_560# AVSS 48.3f
C24 m1_914_2324# AVSS 2.8f
C25 AVDD_1V8 AVSS 31.3f
C26 m1_7138_2408# AVSS 2.8f
C27 INN AVSS 1.47f
C28 INP AVSS 1.46f
C29 li_4275_2335# AVSS 5.94f
.ends
.GLOBAL GND
.end
