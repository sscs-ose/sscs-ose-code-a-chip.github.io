# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o2subcell
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o2subcell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.380000 BY  4.590000 ;
  OBS
    LAYER li1 ;
      RECT 0.000000 0.320000 0.270000 0.460000 ;
      RECT 0.000000 0.460000 3.940000 0.630000 ;
      RECT 0.000000 0.630000 0.270000 1.160000 ;
      RECT 0.000000 1.160000 3.940000 1.330000 ;
      RECT 0.000000 1.330000 0.270000 1.860000 ;
      RECT 0.000000 1.860000 3.940000 2.030000 ;
      RECT 0.000000 2.030000 0.270000 2.560000 ;
      RECT 0.000000 2.560000 3.940000 2.730000 ;
      RECT 0.000000 2.730000 0.270000 3.260000 ;
      RECT 0.000000 3.260000 3.940000 3.430000 ;
      RECT 0.000000 3.430000 0.270000 3.960000 ;
      RECT 0.000000 3.960000 3.940000 4.130000 ;
      RECT 0.440000 0.810000 4.380000 0.980000 ;
      RECT 0.440000 1.510000 4.380000 1.680000 ;
      RECT 0.440000 2.210000 4.380000 2.380000 ;
      RECT 0.440000 2.910000 4.380000 3.080000 ;
      RECT 0.440000 3.610000 4.380000 3.780000 ;
      RECT 4.110000 0.460000 4.380000 0.810000 ;
      RECT 4.110000 0.980000 4.380000 1.510000 ;
      RECT 4.110000 1.680000 4.380000 2.210000 ;
      RECT 4.110000 2.380000 4.380000 2.910000 ;
      RECT 4.110000 3.080000 4.380000 3.610000 ;
      RECT 4.110000 3.780000 4.380000 4.130000 ;
    LAYER mcon ;
      RECT 0.050000 0.450000 0.220000 0.620000 ;
      RECT 0.050000 0.810000 0.220000 0.980000 ;
      RECT 0.050000 1.170000 0.220000 1.340000 ;
      RECT 0.050000 1.530000 0.220000 1.700000 ;
      RECT 0.050000 1.890000 0.220000 2.060000 ;
      RECT 0.050000 2.250000 0.220000 2.420000 ;
      RECT 0.050000 2.610000 0.220000 2.780000 ;
      RECT 0.050000 2.970000 0.220000 3.140000 ;
      RECT 0.050000 3.330000 0.220000 3.500000 ;
      RECT 0.050000 3.690000 0.220000 3.860000 ;
      RECT 4.160000 0.575000 4.330000 0.745000 ;
      RECT 4.160000 0.935000 4.330000 1.105000 ;
      RECT 4.160000 1.295000 4.330000 1.465000 ;
      RECT 4.160000 1.655000 4.330000 1.825000 ;
      RECT 4.160000 2.015000 4.330000 2.185000 ;
      RECT 4.160000 2.375000 4.330000 2.545000 ;
      RECT 4.160000 2.735000 4.330000 2.905000 ;
      RECT 4.160000 3.095000 4.330000 3.265000 ;
      RECT 4.160000 3.455000 4.330000 3.625000 ;
      RECT 4.160000 3.815000 4.330000 3.985000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 4.380000 0.320000 ;
      RECT 0.000000 0.320000 0.270000 4.130000 ;
      RECT 0.000000 4.270000 4.380000 4.590000 ;
      RECT 0.440000 0.320000 0.580000 4.130000 ;
      RECT 0.720000 0.460000 0.860000 4.270000 ;
      RECT 1.000000 0.320000 1.140000 4.130000 ;
      RECT 1.280000 0.460000 1.420000 4.270000 ;
      RECT 1.560000 0.320000 1.700000 4.130000 ;
      RECT 1.840000 0.460000 1.980000 4.270000 ;
      RECT 2.120000 0.320000 2.260000 4.130000 ;
      RECT 2.400000 0.460000 2.540000 4.270000 ;
      RECT 2.680000 0.320000 2.820000 4.130000 ;
      RECT 2.960000 0.460000 3.100000 4.270000 ;
      RECT 3.240000 0.320000 3.380000 4.130000 ;
      RECT 3.520000 0.460000 3.660000 4.270000 ;
      RECT 3.800000 0.320000 3.940000 4.130000 ;
      RECT 4.110000 0.460000 4.380000 4.270000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 4.380000 0.320000 ;
      RECT 0.000000 0.320000 0.270000 4.130000 ;
      RECT 0.000000 4.270000 4.380000 4.590000 ;
      RECT 0.440000 0.460000 0.580000 4.270000 ;
      RECT 0.720000 0.320000 0.860000 4.130000 ;
      RECT 1.000000 0.460000 1.140000 4.270000 ;
      RECT 1.280000 0.320000 1.420000 4.130000 ;
      RECT 1.560000 0.460000 1.700000 4.270000 ;
      RECT 1.840000 0.320000 1.980000 4.130000 ;
      RECT 2.120000 0.460000 2.260000 4.270000 ;
      RECT 2.400000 0.320000 2.540000 4.130000 ;
      RECT 2.680000 0.460000 2.820000 4.270000 ;
      RECT 2.960000 0.320000 3.100000 4.130000 ;
      RECT 3.240000 0.460000 3.380000 4.270000 ;
      RECT 3.520000 0.320000 3.660000 4.130000 ;
      RECT 3.800000 0.460000 3.940000 4.270000 ;
      RECT 4.110000 0.460000 4.380000 4.270000 ;
    LAYER via ;
      RECT 0.005000 0.265000 0.265000 0.525000 ;
      RECT 0.005000 0.585000 0.265000 0.845000 ;
      RECT 0.005000 0.905000 0.265000 1.165000 ;
      RECT 0.005000 1.225000 0.265000 1.485000 ;
      RECT 0.005000 1.545000 0.265000 1.805000 ;
      RECT 0.005000 1.865000 0.265000 2.125000 ;
      RECT 0.005000 2.185000 0.265000 2.445000 ;
      RECT 0.005000 2.505000 0.265000 2.765000 ;
      RECT 0.005000 2.825000 0.265000 3.085000 ;
      RECT 0.005000 3.145000 0.265000 3.405000 ;
      RECT 0.005000 3.465000 0.265000 3.725000 ;
      RECT 0.005000 3.785000 0.265000 4.045000 ;
      RECT 0.380000 0.030000 0.640000 0.290000 ;
      RECT 0.380000 4.300000 0.640000 4.560000 ;
      RECT 0.700000 0.030000 0.960000 0.290000 ;
      RECT 0.700000 4.300000 0.960000 4.560000 ;
      RECT 1.020000 0.030000 1.280000 0.290000 ;
      RECT 1.020000 4.300000 1.280000 4.560000 ;
      RECT 1.340000 0.030000 1.600000 0.290000 ;
      RECT 1.340000 4.300000 1.600000 4.560000 ;
      RECT 1.660000 0.030000 1.920000 0.290000 ;
      RECT 1.660000 4.300000 1.920000 4.560000 ;
      RECT 1.980000 0.030000 2.240000 0.290000 ;
      RECT 1.980000 4.300000 2.240000 4.560000 ;
      RECT 2.300000 0.030000 2.560000 0.290000 ;
      RECT 2.300000 4.300000 2.560000 4.560000 ;
      RECT 2.620000 0.030000 2.880000 0.290000 ;
      RECT 2.620000 4.300000 2.880000 4.560000 ;
      RECT 2.940000 0.030000 3.200000 0.290000 ;
      RECT 2.940000 4.300000 3.200000 4.560000 ;
      RECT 3.260000 0.030000 3.520000 0.290000 ;
      RECT 3.260000 4.300000 3.520000 4.560000 ;
      RECT 3.580000 0.030000 3.840000 0.290000 ;
      RECT 3.580000 4.300000 3.840000 4.560000 ;
      RECT 4.115000 0.490000 4.375000 0.750000 ;
      RECT 4.115000 0.810000 4.375000 1.070000 ;
      RECT 4.115000 1.130000 4.375000 1.390000 ;
      RECT 4.115000 1.450000 4.375000 1.710000 ;
      RECT 4.115000 1.770000 4.375000 2.030000 ;
      RECT 4.115000 2.090000 4.375000 2.350000 ;
      RECT 4.115000 2.410000 4.375000 2.670000 ;
      RECT 4.115000 2.730000 4.375000 2.990000 ;
      RECT 4.115000 3.050000 4.375000 3.310000 ;
      RECT 4.115000 3.370000 4.375000 3.630000 ;
      RECT 4.115000 3.690000 4.375000 3.950000 ;
  END
END sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o2subcell
END LIBRARY
