# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF04W0p84L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF04W0p84L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  2.360000 BY  1.960000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.470400 ;
    PORT
      LAYER met3 ;
        RECT 0.600000 0.215000 0.930000 0.655000 ;
        RECT 0.600000 0.655000 1.790000 0.985000 ;
        RECT 1.460000 0.215000 1.790000 0.655000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.504000 ;
    PORT
      LAYER met1 ;
        RECT 0.510000 1.205000 1.880000 1.495000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.680400 ;
    PORT
      LAYER met1 ;
        RECT 0.220000 -0.445000 2.170000 -0.145000 ;
        RECT 0.220000 -0.145000 0.450000  0.945000 ;
        RECT 1.080000 -0.145000 1.310000  0.945000 ;
        RECT 1.940000 -0.145000 2.170000  0.945000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.250000 0.255000 0.420000 0.945000 ;
      RECT 0.520000 1.175000 1.870000 1.515000 ;
      RECT 0.680000 0.255000 0.850000 0.945000 ;
      RECT 1.110000 0.255000 1.280000 0.945000 ;
      RECT 1.540000 0.255000 1.710000 0.945000 ;
      RECT 1.970000 0.255000 2.140000 0.945000 ;
    LAYER mcon ;
      RECT 0.250000 0.335000 0.420000 0.505000 ;
      RECT 0.250000 0.695000 0.420000 0.865000 ;
      RECT 0.570000 1.265000 0.740000 1.435000 ;
      RECT 0.680000 0.335000 0.850000 0.505000 ;
      RECT 0.680000 0.695000 0.850000 0.865000 ;
      RECT 0.930000 1.265000 1.100000 1.435000 ;
      RECT 1.110000 0.335000 1.280000 0.505000 ;
      RECT 1.110000 0.695000 1.280000 0.865000 ;
      RECT 1.290000 1.265000 1.460000 1.435000 ;
      RECT 1.540000 0.335000 1.710000 0.505000 ;
      RECT 1.540000 0.695000 1.710000 0.865000 ;
      RECT 1.650000 1.265000 1.820000 1.435000 ;
      RECT 1.970000 0.335000 2.140000 0.505000 ;
      RECT 1.970000 0.695000 2.140000 0.865000 ;
    LAYER met1 ;
      RECT 0.635000 0.255000 0.895000 0.945000 ;
      RECT 1.495000 0.255000 1.755000 0.945000 ;
    LAYER met2 ;
      RECT 0.600000 0.215000 0.930000 0.985000 ;
      RECT 1.460000 0.215000 1.790000 0.985000 ;
    LAYER via ;
      RECT 0.635000 0.310000 0.895000 0.570000 ;
      RECT 0.635000 0.630000 0.895000 0.890000 ;
      RECT 1.495000 0.310000 1.755000 0.570000 ;
      RECT 1.495000 0.630000 1.755000 0.890000 ;
    LAYER via2 ;
      RECT 0.625000 0.260000 0.905000 0.540000 ;
      RECT 0.625000 0.660000 0.905000 0.940000 ;
      RECT 1.485000 0.260000 1.765000 0.540000 ;
      RECT 1.485000 0.660000 1.765000 0.940000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF04W0p84L0p15
END LIBRARY
