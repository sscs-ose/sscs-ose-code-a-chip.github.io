# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50 ;
  ORIGIN -0.050000  0.000000 ;
  SIZE  5.020000 BY  8.010000 ;
  PIN DRAIN
    ANTENNADIFFAREA  3.970400 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.405000 5.070000 5.605000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  14.179999 ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.100000 4.085000 0.270000 ;
        RECT 1.035000 7.740000 4.085000 7.910000 ;
      LAYER mcon ;
        RECT 1.215000 0.100000 1.385000 0.270000 ;
        RECT 1.215000 7.740000 1.385000 7.910000 ;
        RECT 1.575000 0.100000 1.745000 0.270000 ;
        RECT 1.575000 7.740000 1.745000 7.910000 ;
        RECT 1.935000 0.100000 2.105000 0.270000 ;
        RECT 1.935000 7.740000 2.105000 7.910000 ;
        RECT 2.295000 0.100000 2.465000 0.270000 ;
        RECT 2.295000 7.740000 2.465000 7.910000 ;
        RECT 2.655000 0.100000 2.825000 0.270000 ;
        RECT 2.655000 7.740000 2.825000 7.910000 ;
        RECT 3.015000 0.100000 3.185000 0.270000 ;
        RECT 3.015000 7.740000 3.185000 7.910000 ;
        RECT 3.375000 0.100000 3.545000 0.270000 ;
        RECT 3.375000 7.740000 3.545000 7.910000 ;
        RECT 3.735000 0.100000 3.905000 0.270000 ;
        RECT 3.735000 7.740000 3.905000 7.910000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.155000 0.000000 3.965000 0.330000 ;
        RECT 1.155000 7.680000 3.965000 8.010000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  5.955600 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.525000 5.070000 2.125000 ;
        RECT 0.050000 5.885000 5.070000 7.485000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  2.056100 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.525000 0.470000 7.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.650000 0.525000 4.940000 7.485000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.440000 0.410000 7.570000 ;
      RECT 0.915000 0.440000 1.085000 7.570000 ;
      RECT 1.695000 0.440000 1.865000 7.570000 ;
      RECT 2.475000 0.440000 2.645000 7.570000 ;
      RECT 3.255000 0.440000 3.425000 7.570000 ;
      RECT 4.035000 0.440000 4.205000 7.570000 ;
      RECT 4.710000 0.610000 4.880000 7.400000 ;
    LAYER mcon ;
      RECT 0.240000 0.680000 0.410000 0.850000 ;
      RECT 0.240000 1.040000 0.410000 1.210000 ;
      RECT 0.240000 1.400000 0.410000 1.570000 ;
      RECT 0.240000 1.760000 0.410000 1.930000 ;
      RECT 0.240000 2.120000 0.410000 2.290000 ;
      RECT 0.240000 2.480000 0.410000 2.650000 ;
      RECT 0.240000 2.840000 0.410000 3.010000 ;
      RECT 0.240000 3.200000 0.410000 3.370000 ;
      RECT 0.240000 3.560000 0.410000 3.730000 ;
      RECT 0.240000 3.920000 0.410000 4.090000 ;
      RECT 0.240000 4.280000 0.410000 4.450000 ;
      RECT 0.240000 4.640000 0.410000 4.810000 ;
      RECT 0.240000 5.000000 0.410000 5.170000 ;
      RECT 0.240000 5.360000 0.410000 5.530000 ;
      RECT 0.240000 5.720000 0.410000 5.890000 ;
      RECT 0.240000 6.080000 0.410000 6.250000 ;
      RECT 0.240000 6.440000 0.410000 6.610000 ;
      RECT 0.240000 6.800000 0.410000 6.970000 ;
      RECT 0.240000 7.160000 0.410000 7.330000 ;
      RECT 0.915000 0.680000 1.085000 0.850000 ;
      RECT 0.915000 1.040000 1.085000 1.210000 ;
      RECT 0.915000 1.400000 1.085000 1.570000 ;
      RECT 0.915000 1.760000 1.085000 1.930000 ;
      RECT 0.915000 2.120000 1.085000 2.290000 ;
      RECT 0.915000 2.480000 1.085000 2.650000 ;
      RECT 0.915000 2.840000 1.085000 3.010000 ;
      RECT 0.915000 3.200000 1.085000 3.370000 ;
      RECT 0.915000 3.560000 1.085000 3.730000 ;
      RECT 0.915000 3.920000 1.085000 4.090000 ;
      RECT 0.915000 4.280000 1.085000 4.450000 ;
      RECT 0.915000 4.640000 1.085000 4.810000 ;
      RECT 0.915000 5.000000 1.085000 5.170000 ;
      RECT 0.915000 5.360000 1.085000 5.530000 ;
      RECT 0.915000 5.720000 1.085000 5.890000 ;
      RECT 0.915000 6.080000 1.085000 6.250000 ;
      RECT 0.915000 6.440000 1.085000 6.610000 ;
      RECT 0.915000 6.800000 1.085000 6.970000 ;
      RECT 0.915000 7.160000 1.085000 7.330000 ;
      RECT 1.695000 0.680000 1.865000 0.850000 ;
      RECT 1.695000 1.040000 1.865000 1.210000 ;
      RECT 1.695000 1.400000 1.865000 1.570000 ;
      RECT 1.695000 1.760000 1.865000 1.930000 ;
      RECT 1.695000 2.120000 1.865000 2.290000 ;
      RECT 1.695000 2.480000 1.865000 2.650000 ;
      RECT 1.695000 2.840000 1.865000 3.010000 ;
      RECT 1.695000 3.200000 1.865000 3.370000 ;
      RECT 1.695000 3.560000 1.865000 3.730000 ;
      RECT 1.695000 3.920000 1.865000 4.090000 ;
      RECT 1.695000 4.280000 1.865000 4.450000 ;
      RECT 1.695000 4.640000 1.865000 4.810000 ;
      RECT 1.695000 5.000000 1.865000 5.170000 ;
      RECT 1.695000 5.360000 1.865000 5.530000 ;
      RECT 1.695000 5.720000 1.865000 5.890000 ;
      RECT 1.695000 6.080000 1.865000 6.250000 ;
      RECT 1.695000 6.440000 1.865000 6.610000 ;
      RECT 1.695000 6.800000 1.865000 6.970000 ;
      RECT 1.695000 7.160000 1.865000 7.330000 ;
      RECT 2.475000 0.680000 2.645000 0.850000 ;
      RECT 2.475000 1.040000 2.645000 1.210000 ;
      RECT 2.475000 1.400000 2.645000 1.570000 ;
      RECT 2.475000 1.760000 2.645000 1.930000 ;
      RECT 2.475000 2.120000 2.645000 2.290000 ;
      RECT 2.475000 2.480000 2.645000 2.650000 ;
      RECT 2.475000 2.840000 2.645000 3.010000 ;
      RECT 2.475000 3.200000 2.645000 3.370000 ;
      RECT 2.475000 3.560000 2.645000 3.730000 ;
      RECT 2.475000 3.920000 2.645000 4.090000 ;
      RECT 2.475000 4.280000 2.645000 4.450000 ;
      RECT 2.475000 4.640000 2.645000 4.810000 ;
      RECT 2.475000 5.000000 2.645000 5.170000 ;
      RECT 2.475000 5.360000 2.645000 5.530000 ;
      RECT 2.475000 5.720000 2.645000 5.890000 ;
      RECT 2.475000 6.080000 2.645000 6.250000 ;
      RECT 2.475000 6.440000 2.645000 6.610000 ;
      RECT 2.475000 6.800000 2.645000 6.970000 ;
      RECT 2.475000 7.160000 2.645000 7.330000 ;
      RECT 3.255000 0.680000 3.425000 0.850000 ;
      RECT 3.255000 1.040000 3.425000 1.210000 ;
      RECT 3.255000 1.400000 3.425000 1.570000 ;
      RECT 3.255000 1.760000 3.425000 1.930000 ;
      RECT 3.255000 2.120000 3.425000 2.290000 ;
      RECT 3.255000 2.480000 3.425000 2.650000 ;
      RECT 3.255000 2.840000 3.425000 3.010000 ;
      RECT 3.255000 3.200000 3.425000 3.370000 ;
      RECT 3.255000 3.560000 3.425000 3.730000 ;
      RECT 3.255000 3.920000 3.425000 4.090000 ;
      RECT 3.255000 4.280000 3.425000 4.450000 ;
      RECT 3.255000 4.640000 3.425000 4.810000 ;
      RECT 3.255000 5.000000 3.425000 5.170000 ;
      RECT 3.255000 5.360000 3.425000 5.530000 ;
      RECT 3.255000 5.720000 3.425000 5.890000 ;
      RECT 3.255000 6.080000 3.425000 6.250000 ;
      RECT 3.255000 6.440000 3.425000 6.610000 ;
      RECT 3.255000 6.800000 3.425000 6.970000 ;
      RECT 3.255000 7.160000 3.425000 7.330000 ;
      RECT 4.035000 0.680000 4.205000 0.850000 ;
      RECT 4.035000 1.040000 4.205000 1.210000 ;
      RECT 4.035000 1.400000 4.205000 1.570000 ;
      RECT 4.035000 1.760000 4.205000 1.930000 ;
      RECT 4.035000 2.120000 4.205000 2.290000 ;
      RECT 4.035000 2.480000 4.205000 2.650000 ;
      RECT 4.035000 2.840000 4.205000 3.010000 ;
      RECT 4.035000 3.200000 4.205000 3.370000 ;
      RECT 4.035000 3.560000 4.205000 3.730000 ;
      RECT 4.035000 3.920000 4.205000 4.090000 ;
      RECT 4.035000 4.280000 4.205000 4.450000 ;
      RECT 4.035000 4.640000 4.205000 4.810000 ;
      RECT 4.035000 5.000000 4.205000 5.170000 ;
      RECT 4.035000 5.360000 4.205000 5.530000 ;
      RECT 4.035000 5.720000 4.205000 5.890000 ;
      RECT 4.035000 6.080000 4.205000 6.250000 ;
      RECT 4.035000 6.440000 4.205000 6.610000 ;
      RECT 4.035000 6.800000 4.205000 6.970000 ;
      RECT 4.035000 7.160000 4.205000 7.330000 ;
      RECT 4.710000 0.680000 4.880000 0.850000 ;
      RECT 4.710000 1.040000 4.880000 1.210000 ;
      RECT 4.710000 1.400000 4.880000 1.570000 ;
      RECT 4.710000 1.760000 4.880000 1.930000 ;
      RECT 4.710000 2.120000 4.880000 2.290000 ;
      RECT 4.710000 2.480000 4.880000 2.650000 ;
      RECT 4.710000 2.840000 4.880000 3.010000 ;
      RECT 4.710000 3.200000 4.880000 3.370000 ;
      RECT 4.710000 3.560000 4.880000 3.730000 ;
      RECT 4.710000 3.920000 4.880000 4.090000 ;
      RECT 4.710000 4.280000 4.880000 4.450000 ;
      RECT 4.710000 4.640000 4.880000 4.810000 ;
      RECT 4.710000 5.000000 4.880000 5.170000 ;
      RECT 4.710000 5.360000 4.880000 5.530000 ;
      RECT 4.710000 5.720000 4.880000 5.890000 ;
      RECT 4.710000 6.080000 4.880000 6.250000 ;
      RECT 4.710000 6.440000 4.880000 6.610000 ;
      RECT 4.710000 6.800000 4.880000 6.970000 ;
      RECT 4.710000 7.160000 4.880000 7.330000 ;
    LAYER met1 ;
      RECT 0.870000 0.525000 1.130000 7.485000 ;
      RECT 1.650000 0.525000 1.910000 7.485000 ;
      RECT 2.430000 0.525000 2.690000 7.485000 ;
      RECT 3.210000 0.525000 3.470000 7.485000 ;
      RECT 3.990000 0.525000 4.250000 7.485000 ;
    LAYER via ;
      RECT 0.870000 0.555000 1.130000 0.815000 ;
      RECT 0.870000 0.875000 1.130000 1.135000 ;
      RECT 0.870000 1.195000 1.130000 1.455000 ;
      RECT 0.870000 1.515000 1.130000 1.775000 ;
      RECT 0.870000 1.835000 1.130000 2.095000 ;
      RECT 0.870000 5.915000 1.130000 6.175000 ;
      RECT 0.870000 6.235000 1.130000 6.495000 ;
      RECT 0.870000 6.555000 1.130000 6.815000 ;
      RECT 0.870000 6.875000 1.130000 7.135000 ;
      RECT 0.870000 7.195000 1.130000 7.455000 ;
      RECT 1.650000 2.435000 1.910000 2.695000 ;
      RECT 1.650000 2.755000 1.910000 3.015000 ;
      RECT 1.650000 3.075000 1.910000 3.335000 ;
      RECT 1.650000 3.395000 1.910000 3.655000 ;
      RECT 1.650000 3.715000 1.910000 3.975000 ;
      RECT 1.650000 4.035000 1.910000 4.295000 ;
      RECT 1.650000 4.355000 1.910000 4.615000 ;
      RECT 1.650000 4.675000 1.910000 4.935000 ;
      RECT 1.650000 4.995000 1.910000 5.255000 ;
      RECT 1.650000 5.315000 1.910000 5.575000 ;
      RECT 2.430000 0.555000 2.690000 0.815000 ;
      RECT 2.430000 0.875000 2.690000 1.135000 ;
      RECT 2.430000 1.195000 2.690000 1.455000 ;
      RECT 2.430000 1.515000 2.690000 1.775000 ;
      RECT 2.430000 1.835000 2.690000 2.095000 ;
      RECT 2.430000 5.915000 2.690000 6.175000 ;
      RECT 2.430000 6.235000 2.690000 6.495000 ;
      RECT 2.430000 6.555000 2.690000 6.815000 ;
      RECT 2.430000 6.875000 2.690000 7.135000 ;
      RECT 2.430000 7.195000 2.690000 7.455000 ;
      RECT 3.210000 2.435000 3.470000 2.695000 ;
      RECT 3.210000 2.755000 3.470000 3.015000 ;
      RECT 3.210000 3.075000 3.470000 3.335000 ;
      RECT 3.210000 3.395000 3.470000 3.655000 ;
      RECT 3.210000 3.715000 3.470000 3.975000 ;
      RECT 3.210000 4.035000 3.470000 4.295000 ;
      RECT 3.210000 4.355000 3.470000 4.615000 ;
      RECT 3.210000 4.675000 3.470000 4.935000 ;
      RECT 3.210000 4.995000 3.470000 5.255000 ;
      RECT 3.210000 5.315000 3.470000 5.575000 ;
      RECT 3.990000 0.555000 4.250000 0.815000 ;
      RECT 3.990000 0.875000 4.250000 1.135000 ;
      RECT 3.990000 1.195000 4.250000 1.455000 ;
      RECT 3.990000 1.515000 4.250000 1.775000 ;
      RECT 3.990000 1.835000 4.250000 2.095000 ;
      RECT 3.990000 5.915000 4.250000 6.175000 ;
      RECT 3.990000 6.235000 4.250000 6.495000 ;
      RECT 3.990000 6.555000 4.250000 6.815000 ;
      RECT 3.990000 6.875000 4.250000 7.135000 ;
      RECT 3.990000 7.195000 4.250000 7.455000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50
END LIBRARY
