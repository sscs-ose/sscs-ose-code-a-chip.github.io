# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.800000 BY  6.090000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT 0.000000 0.000000 6.800000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 5.760000 ;
        RECT 0.000000 5.760000 6.800000 6.090000 ;
        RECT 1.270000 0.330000 1.610000 2.580000 ;
        RECT 1.270000 3.510000 1.610000 5.760000 ;
        RECT 2.550000 0.330000 2.890000 2.580000 ;
        RECT 2.550000 3.510000 2.890000 5.760000 ;
        RECT 3.910000 0.330000 4.250000 2.580000 ;
        RECT 3.910000 3.510000 4.250000 5.760000 ;
        RECT 5.190000 0.330000 5.530000 2.580000 ;
        RECT 5.190000 3.510000 5.530000 5.760000 ;
        RECT 6.470000 0.330000 6.800000 5.760000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT 0.630000 0.630000 0.970000 2.880000 ;
        RECT 0.630000 2.880000 6.170000 3.210000 ;
        RECT 0.630000 3.210000 0.970000 5.460000 ;
        RECT 1.910000 0.630000 2.250000 2.880000 ;
        RECT 1.910000 3.210000 2.250000 5.460000 ;
        RECT 3.190000 0.630000 3.610000 2.880000 ;
        RECT 3.190000 3.210000 3.610000 5.460000 ;
        RECT 4.550000 0.630000 4.890000 2.880000 ;
        RECT 4.550000 3.210000 4.890000 5.460000 ;
        RECT 5.830000 0.630000 6.170000 2.880000 ;
        RECT 5.830000 3.210000 6.170000 5.460000 ;
    END
  END C1
  PIN MET4
    PORT
      LAYER met4 ;
        RECT 0.000000 0.000000 6.800000 6.090000 ;
    END
  END MET4
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 2.735000 4.370000 2.840000 4.615000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 6.800000 6.090000 ;
    LAYER mcon ;
      RECT 0.080000 0.440000 0.250000 0.610000 ;
      RECT 0.080000 0.800000 0.250000 0.970000 ;
      RECT 0.080000 1.160000 0.250000 1.330000 ;
      RECT 0.080000 1.520000 0.250000 1.690000 ;
      RECT 0.080000 1.880000 0.250000 2.050000 ;
      RECT 0.080000 2.240000 0.250000 2.410000 ;
      RECT 0.080000 2.600000 0.250000 2.770000 ;
      RECT 0.080000 2.960000 0.250000 3.130000 ;
      RECT 0.080000 3.320000 0.250000 3.490000 ;
      RECT 0.080000 3.680000 0.250000 3.850000 ;
      RECT 0.080000 4.040000 0.250000 4.210000 ;
      RECT 0.080000 4.400000 0.250000 4.570000 ;
      RECT 0.080000 4.760000 0.250000 4.930000 ;
      RECT 0.080000 5.120000 0.250000 5.290000 ;
      RECT 0.080000 5.480000 0.250000 5.650000 ;
      RECT 0.410000 0.080000 0.580000 0.250000 ;
      RECT 0.410000 5.840000 0.580000 6.010000 ;
      RECT 0.770000 0.080000 0.940000 0.250000 ;
      RECT 0.770000 5.840000 0.940000 6.010000 ;
      RECT 1.130000 0.080000 1.300000 0.250000 ;
      RECT 1.130000 5.840000 1.300000 6.010000 ;
      RECT 1.490000 0.080000 1.660000 0.250000 ;
      RECT 1.490000 5.840000 1.660000 6.010000 ;
      RECT 1.850000 0.080000 2.020000 0.250000 ;
      RECT 1.850000 5.840000 2.020000 6.010000 ;
      RECT 2.210000 0.080000 2.380000 0.250000 ;
      RECT 2.210000 5.840000 2.380000 6.010000 ;
      RECT 2.570000 0.080000 2.740000 0.250000 ;
      RECT 2.570000 5.840000 2.740000 6.010000 ;
      RECT 2.930000 0.080000 3.100000 0.250000 ;
      RECT 2.930000 5.840000 3.100000 6.010000 ;
      RECT 3.315000 0.080000 3.485000 0.250000 ;
      RECT 3.315000 5.840000 3.485000 6.010000 ;
      RECT 3.700000 0.080000 3.870000 0.250000 ;
      RECT 3.700000 5.840000 3.870000 6.010000 ;
      RECT 4.060000 0.080000 4.230000 0.250000 ;
      RECT 4.060000 5.840000 4.230000 6.010000 ;
      RECT 4.420000 0.080000 4.590000 0.250000 ;
      RECT 4.420000 5.840000 4.590000 6.010000 ;
      RECT 4.780000 0.080000 4.950000 0.250000 ;
      RECT 4.780000 5.840000 4.950000 6.010000 ;
      RECT 5.140000 0.080000 5.310000 0.250000 ;
      RECT 5.140000 5.840000 5.310000 6.010000 ;
      RECT 5.500000 0.080000 5.670000 0.250000 ;
      RECT 5.500000 5.840000 5.670000 6.010000 ;
      RECT 5.860000 0.080000 6.030000 0.250000 ;
      RECT 5.860000 5.840000 6.030000 6.010000 ;
      RECT 6.220000 0.080000 6.390000 0.250000 ;
      RECT 6.220000 5.840000 6.390000 6.010000 ;
      RECT 6.550000 0.440000 6.720000 0.610000 ;
      RECT 6.550000 0.800000 6.720000 0.970000 ;
      RECT 6.550000 1.160000 6.720000 1.330000 ;
      RECT 6.550000 1.520000 6.720000 1.690000 ;
      RECT 6.550000 1.880000 6.720000 2.050000 ;
      RECT 6.550000 2.240000 6.720000 2.410000 ;
      RECT 6.550000 2.600000 6.720000 2.770000 ;
      RECT 6.550000 2.960000 6.720000 3.130000 ;
      RECT 6.550000 3.320000 6.720000 3.490000 ;
      RECT 6.550000 3.680000 6.720000 3.850000 ;
      RECT 6.550000 4.040000 6.720000 4.210000 ;
      RECT 6.550000 4.400000 6.720000 4.570000 ;
      RECT 6.550000 4.760000 6.720000 4.930000 ;
      RECT 6.550000 5.120000 6.720000 5.290000 ;
      RECT 6.550000 5.480000 6.720000 5.650000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 6.800000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 5.760000 ;
      RECT 0.000000 5.760000 6.800000 6.090000 ;
      RECT 0.470000 0.470000 0.610000 2.885000 ;
      RECT 0.470000 2.885000 6.330000 3.205000 ;
      RECT 0.470000 3.205000 0.610000 5.620000 ;
      RECT 0.750000 0.330000 0.890000 2.745000 ;
      RECT 0.750000 3.345000 0.890000 5.760000 ;
      RECT 1.030000 0.470000 1.170000 2.885000 ;
      RECT 1.030000 3.205000 1.170000 5.620000 ;
      RECT 1.310000 0.330000 1.450000 2.745000 ;
      RECT 1.310000 3.345000 1.450000 5.760000 ;
      RECT 1.590000 0.470000 1.730000 2.885000 ;
      RECT 1.590000 3.205000 1.730000 5.620000 ;
      RECT 1.870000 0.330000 2.010000 2.745000 ;
      RECT 1.870000 3.345000 2.010000 5.760000 ;
      RECT 2.150000 0.470000 2.290000 2.885000 ;
      RECT 2.150000 3.205000 2.290000 5.620000 ;
      RECT 2.430000 0.330000 2.570000 2.745000 ;
      RECT 2.430000 3.345000 2.570000 5.760000 ;
      RECT 2.710000 0.470000 2.850000 2.885000 ;
      RECT 2.710000 3.205000 2.850000 5.620000 ;
      RECT 2.990000 0.330000 3.130000 2.745000 ;
      RECT 2.990000 3.345000 3.130000 5.760000 ;
      RECT 3.270000 0.470000 3.530000 2.885000 ;
      RECT 3.270000 3.205000 3.530000 5.620000 ;
      RECT 3.670000 0.330000 3.810000 2.745000 ;
      RECT 3.670000 3.345000 3.810000 5.760000 ;
      RECT 3.950000 0.470000 4.090000 2.885000 ;
      RECT 3.950000 3.205000 4.090000 5.620000 ;
      RECT 4.230000 0.330000 4.370000 2.745000 ;
      RECT 4.230000 3.345000 4.370000 5.760000 ;
      RECT 4.510000 0.470000 4.650000 2.885000 ;
      RECT 4.510000 3.205000 4.650000 5.620000 ;
      RECT 4.790000 0.330000 4.930000 2.745000 ;
      RECT 4.790000 3.345000 4.930000 5.760000 ;
      RECT 5.070000 0.470000 5.210000 2.885000 ;
      RECT 5.070000 3.205000 5.210000 5.620000 ;
      RECT 5.350000 0.330000 5.490000 2.745000 ;
      RECT 5.350000 3.345000 5.490000 5.760000 ;
      RECT 5.630000 0.470000 5.770000 2.885000 ;
      RECT 5.630000 3.205000 5.770000 5.620000 ;
      RECT 5.910000 0.330000 6.050000 2.745000 ;
      RECT 5.910000 3.345000 6.050000 5.760000 ;
      RECT 6.190000 0.470000 6.330000 2.885000 ;
      RECT 6.190000 3.205000 6.330000 5.620000 ;
      RECT 6.470000 0.330000 6.800000 5.760000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 3.095000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 0.750000 ;
      RECT 0.000000 0.750000 3.095000 0.890000 ;
      RECT 0.000000 0.890000 0.330000 1.310000 ;
      RECT 0.000000 1.310000 3.095000 1.450000 ;
      RECT 0.000000 1.450000 0.330000 1.870000 ;
      RECT 0.000000 1.870000 3.095000 2.010000 ;
      RECT 0.000000 2.010000 0.330000 2.430000 ;
      RECT 0.000000 2.430000 3.095000 2.765000 ;
      RECT 0.000000 2.905000 6.800000 3.185000 ;
      RECT 0.000000 3.325000 3.095000 3.660000 ;
      RECT 0.000000 3.660000 0.330000 4.080000 ;
      RECT 0.000000 4.080000 3.095000 4.220000 ;
      RECT 0.000000 4.220000 0.330000 4.640000 ;
      RECT 0.000000 4.640000 3.095000 4.780000 ;
      RECT 0.000000 4.780000 0.330000 5.200000 ;
      RECT 0.000000 5.200000 3.095000 5.340000 ;
      RECT 0.000000 5.340000 0.330000 5.760000 ;
      RECT 0.000000 5.760000 3.095000 6.090000 ;
      RECT 0.470000 0.470000 6.330000 0.610000 ;
      RECT 0.470000 1.030000 6.330000 1.170000 ;
      RECT 0.470000 1.590000 6.330000 1.730000 ;
      RECT 0.470000 2.150000 6.330000 2.290000 ;
      RECT 0.470000 3.800000 6.330000 3.940000 ;
      RECT 0.470000 4.360000 6.330000 4.500000 ;
      RECT 0.470000 4.920000 6.330000 5.060000 ;
      RECT 0.470000 5.480000 6.330000 5.620000 ;
      RECT 3.235000 0.000000 3.565000 0.470000 ;
      RECT 3.235000 0.610000 3.565000 1.030000 ;
      RECT 3.235000 1.170000 3.565000 1.590000 ;
      RECT 3.235000 1.730000 3.565000 2.150000 ;
      RECT 3.235000 2.290000 3.565000 2.905000 ;
      RECT 3.235000 3.185000 3.565000 3.800000 ;
      RECT 3.235000 3.940000 3.565000 4.360000 ;
      RECT 3.235000 4.500000 3.565000 4.920000 ;
      RECT 3.235000 5.060000 3.565000 5.480000 ;
      RECT 3.235000 5.620000 3.565000 6.090000 ;
      RECT 3.705000 0.000000 6.800000 0.330000 ;
      RECT 3.705000 0.750000 6.800000 0.890000 ;
      RECT 3.705000 1.310000 6.800000 1.450000 ;
      RECT 3.705000 1.870000 6.800000 2.010000 ;
      RECT 3.705000 2.430000 6.800000 2.765000 ;
      RECT 3.705000 3.325000 6.800000 3.660000 ;
      RECT 3.705000 4.080000 6.800000 4.220000 ;
      RECT 3.705000 4.640000 6.800000 4.780000 ;
      RECT 3.705000 5.200000 6.800000 5.340000 ;
      RECT 3.705000 5.760000 6.800000 6.090000 ;
      RECT 6.470000 0.330000 6.800000 0.750000 ;
      RECT 6.470000 0.890000 6.800000 1.310000 ;
      RECT 6.470000 1.450000 6.800000 1.870000 ;
      RECT 6.470000 2.010000 6.800000 2.430000 ;
      RECT 6.470000 3.660000 6.800000 4.080000 ;
      RECT 6.470000 4.220000 6.800000 4.640000 ;
      RECT 6.470000 4.780000 6.800000 5.200000 ;
      RECT 6.470000 5.340000 6.800000 5.760000 ;
    LAYER via ;
      RECT 0.035000 0.355000 0.295000 0.615000 ;
      RECT 0.035000 0.675000 0.295000 0.935000 ;
      RECT 0.035000 0.995000 0.295000 1.255000 ;
      RECT 0.035000 1.315000 0.295000 1.575000 ;
      RECT 0.035000 1.635000 0.295000 1.895000 ;
      RECT 0.035000 1.955000 0.295000 2.215000 ;
      RECT 0.035000 2.275000 0.295000 2.535000 ;
      RECT 0.035000 3.555000 0.295000 3.815000 ;
      RECT 0.035000 3.875000 0.295000 4.135000 ;
      RECT 0.035000 4.195000 0.295000 4.455000 ;
      RECT 0.035000 4.515000 0.295000 4.775000 ;
      RECT 0.035000 4.835000 0.295000 5.095000 ;
      RECT 0.035000 5.155000 0.295000 5.415000 ;
      RECT 0.035000 5.475000 0.295000 5.735000 ;
      RECT 0.365000 0.035000 0.625000 0.295000 ;
      RECT 0.365000 5.795000 0.625000 6.055000 ;
      RECT 0.525000 2.915000 0.785000 3.175000 ;
      RECT 0.685000 0.035000 0.945000 0.295000 ;
      RECT 0.685000 5.795000 0.945000 6.055000 ;
      RECT 0.845000 2.915000 1.105000 3.175000 ;
      RECT 1.005000 0.035000 1.265000 0.295000 ;
      RECT 1.005000 5.795000 1.265000 6.055000 ;
      RECT 1.165000 2.915000 1.425000 3.175000 ;
      RECT 1.325000 0.035000 1.585000 0.295000 ;
      RECT 1.325000 5.795000 1.585000 6.055000 ;
      RECT 1.485000 2.915000 1.745000 3.175000 ;
      RECT 1.645000 0.035000 1.905000 0.295000 ;
      RECT 1.645000 5.795000 1.905000 6.055000 ;
      RECT 1.805000 2.915000 2.065000 3.175000 ;
      RECT 1.965000 0.035000 2.225000 0.295000 ;
      RECT 1.965000 5.795000 2.225000 6.055000 ;
      RECT 2.125000 2.915000 2.385000 3.175000 ;
      RECT 2.285000 0.035000 2.545000 0.295000 ;
      RECT 2.285000 5.795000 2.545000 6.055000 ;
      RECT 2.445000 2.915000 2.705000 3.175000 ;
      RECT 2.605000 0.035000 2.865000 0.295000 ;
      RECT 2.605000 5.795000 2.865000 6.055000 ;
      RECT 2.765000 2.915000 3.025000 3.175000 ;
      RECT 3.085000 2.915000 3.345000 3.175000 ;
      RECT 3.270000 0.515000 3.530000 0.775000 ;
      RECT 3.270000 0.835000 3.530000 1.095000 ;
      RECT 3.270000 1.155000 3.530000 1.415000 ;
      RECT 3.270000 1.475000 3.530000 1.735000 ;
      RECT 3.270000 1.795000 3.530000 2.055000 ;
      RECT 3.270000 2.115000 3.530000 2.375000 ;
      RECT 3.270000 2.435000 3.530000 2.695000 ;
      RECT 3.270000 3.395000 3.530000 3.655000 ;
      RECT 3.270000 3.715000 3.530000 3.975000 ;
      RECT 3.270000 4.035000 3.530000 4.295000 ;
      RECT 3.270000 4.355000 3.530000 4.615000 ;
      RECT 3.270000 4.675000 3.530000 4.935000 ;
      RECT 3.270000 4.995000 3.530000 5.255000 ;
      RECT 3.270000 5.315000 3.530000 5.575000 ;
      RECT 3.455000 2.915000 3.715000 3.175000 ;
      RECT 3.775000 2.915000 4.035000 3.175000 ;
      RECT 3.935000 0.035000 4.195000 0.295000 ;
      RECT 3.935000 5.795000 4.195000 6.055000 ;
      RECT 4.095000 2.915000 4.355000 3.175000 ;
      RECT 4.255000 0.035000 4.515000 0.295000 ;
      RECT 4.255000 5.795000 4.515000 6.055000 ;
      RECT 4.415000 2.915000 4.675000 3.175000 ;
      RECT 4.575000 0.035000 4.835000 0.295000 ;
      RECT 4.575000 5.795000 4.835000 6.055000 ;
      RECT 4.735000 2.915000 4.995000 3.175000 ;
      RECT 4.895000 0.035000 5.155000 0.295000 ;
      RECT 4.895000 5.795000 5.155000 6.055000 ;
      RECT 5.055000 2.915000 5.315000 3.175000 ;
      RECT 5.215000 0.035000 5.475000 0.295000 ;
      RECT 5.215000 5.795000 5.475000 6.055000 ;
      RECT 5.375000 2.915000 5.635000 3.175000 ;
      RECT 5.535000 0.035000 5.795000 0.295000 ;
      RECT 5.535000 5.795000 5.795000 6.055000 ;
      RECT 5.695000 2.915000 5.955000 3.175000 ;
      RECT 5.855000 0.035000 6.115000 0.295000 ;
      RECT 5.855000 5.795000 6.115000 6.055000 ;
      RECT 6.015000 2.915000 6.275000 3.175000 ;
      RECT 6.175000 0.035000 6.435000 0.295000 ;
      RECT 6.175000 5.795000 6.435000 6.055000 ;
      RECT 6.505000 0.355000 6.765000 0.615000 ;
      RECT 6.505000 0.675000 6.765000 0.935000 ;
      RECT 6.505000 0.995000 6.765000 1.255000 ;
      RECT 6.505000 1.315000 6.765000 1.575000 ;
      RECT 6.505000 1.635000 6.765000 1.895000 ;
      RECT 6.505000 1.955000 6.765000 2.215000 ;
      RECT 6.505000 2.275000 6.765000 2.535000 ;
      RECT 6.505000 3.555000 6.765000 3.815000 ;
      RECT 6.505000 3.875000 6.765000 4.135000 ;
      RECT 6.505000 4.195000 6.765000 4.455000 ;
      RECT 6.505000 4.515000 6.765000 4.775000 ;
      RECT 6.505000 4.835000 6.765000 5.095000 ;
      RECT 6.505000 5.155000 6.765000 5.415000 ;
      RECT 6.505000 5.475000 6.765000 5.735000 ;
    LAYER via2 ;
      RECT 0.025000 0.400000 0.305000 0.680000 ;
      RECT 0.025000 0.800000 0.305000 1.080000 ;
      RECT 0.025000 1.200000 0.305000 1.480000 ;
      RECT 0.025000 1.600000 0.305000 1.880000 ;
      RECT 0.025000 2.000000 0.305000 2.280000 ;
      RECT 0.025000 2.400000 0.305000 2.680000 ;
      RECT 0.025000 3.410000 0.305000 3.690000 ;
      RECT 0.025000 3.810000 0.305000 4.090000 ;
      RECT 0.025000 4.210000 0.305000 4.490000 ;
      RECT 0.025000 4.610000 0.305000 4.890000 ;
      RECT 0.025000 5.010000 0.305000 5.290000 ;
      RECT 0.025000 5.410000 0.305000 5.690000 ;
      RECT 0.440000 0.025000 0.720000 0.305000 ;
      RECT 0.440000 5.785000 0.720000 6.065000 ;
      RECT 0.835000 2.905000 1.115000 3.185000 ;
      RECT 0.840000 0.025000 1.120000 0.305000 ;
      RECT 0.840000 5.785000 1.120000 6.065000 ;
      RECT 1.235000 2.905000 1.515000 3.185000 ;
      RECT 1.240000 0.025000 1.520000 0.305000 ;
      RECT 1.240000 5.785000 1.520000 6.065000 ;
      RECT 1.635000 2.905000 1.915000 3.185000 ;
      RECT 1.640000 0.025000 1.920000 0.305000 ;
      RECT 1.640000 5.785000 1.920000 6.065000 ;
      RECT 2.035000 2.905000 2.315000 3.185000 ;
      RECT 2.040000 0.025000 2.320000 0.305000 ;
      RECT 2.040000 5.785000 2.320000 6.065000 ;
      RECT 2.435000 2.905000 2.715000 3.185000 ;
      RECT 2.440000 0.025000 2.720000 0.305000 ;
      RECT 2.440000 5.785000 2.720000 6.065000 ;
      RECT 2.835000 2.905000 3.115000 3.185000 ;
      RECT 3.255000 0.705000 3.535000 0.985000 ;
      RECT 3.255000 1.105000 3.535000 1.385000 ;
      RECT 3.255000 1.505000 3.535000 1.785000 ;
      RECT 3.255000 1.905000 3.535000 2.185000 ;
      RECT 3.255000 2.305000 3.535000 2.585000 ;
      RECT 3.255000 3.505000 3.535000 3.785000 ;
      RECT 3.255000 3.905000 3.535000 4.185000 ;
      RECT 3.255000 4.305000 3.535000 4.585000 ;
      RECT 3.255000 4.705000 3.535000 4.985000 ;
      RECT 3.255000 5.105000 3.535000 5.385000 ;
      RECT 3.260000 2.905000 3.540000 3.185000 ;
      RECT 3.685000 2.905000 3.965000 3.185000 ;
      RECT 4.085000 2.905000 4.365000 3.185000 ;
      RECT 4.090000 0.025000 4.370000 0.305000 ;
      RECT 4.090000 5.785000 4.370000 6.065000 ;
      RECT 4.485000 2.905000 4.765000 3.185000 ;
      RECT 4.490000 0.025000 4.770000 0.305000 ;
      RECT 4.490000 5.785000 4.770000 6.065000 ;
      RECT 4.885000 2.905000 5.165000 3.185000 ;
      RECT 4.890000 0.025000 5.170000 0.305000 ;
      RECT 4.890000 5.785000 5.170000 6.065000 ;
      RECT 5.285000 2.905000 5.565000 3.185000 ;
      RECT 5.290000 0.025000 5.570000 0.305000 ;
      RECT 5.290000 5.785000 5.570000 6.065000 ;
      RECT 5.685000 2.905000 5.965000 3.185000 ;
      RECT 5.690000 0.025000 5.970000 0.305000 ;
      RECT 5.690000 5.785000 5.970000 6.065000 ;
      RECT 6.090000 0.025000 6.370000 0.305000 ;
      RECT 6.090000 5.785000 6.370000 6.065000 ;
      RECT 6.495000 0.400000 6.775000 0.680000 ;
      RECT 6.495000 0.800000 6.775000 1.080000 ;
      RECT 6.495000 1.200000 6.775000 1.480000 ;
      RECT 6.495000 1.600000 6.775000 1.880000 ;
      RECT 6.495000 2.000000 6.775000 2.280000 ;
      RECT 6.495000 2.400000 6.775000 2.680000 ;
      RECT 6.495000 3.410000 6.775000 3.690000 ;
      RECT 6.495000 3.810000 6.775000 4.090000 ;
      RECT 6.495000 4.210000 6.775000 4.490000 ;
      RECT 6.495000 4.610000 6.775000 4.890000 ;
      RECT 6.495000 5.010000 6.775000 5.290000 ;
      RECT 6.495000 5.410000 6.775000 5.690000 ;
  END
END sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4
END LIBRARY
