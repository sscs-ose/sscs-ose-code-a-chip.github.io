# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  9.660000 BY  5.970000 ;
  PIN DRAIN
    ANTENNADIFFAREA  7.070000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 3.110000 9.730000 5.470000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  25.25000 ;
    PORT
      LAYER met1 ;
        RECT 0.975000 0.000000 8.825000 0.330000 ;
        RECT 0.975000 5.640000 8.825000 5.970000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  8.484000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 0.500000 9.730000 2.860000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.464500 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.500000 0.475000 5.470000 ;
    END
    PORT
      LAYER met1 ;
        RECT 9.330000 0.500000 9.625000 5.470000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.560000 0.410000 5.410000 ;
      RECT 0.915000 0.440000 1.085000 5.530000 ;
      RECT 0.995000 0.100000 8.805000 0.270000 ;
      RECT 0.995000 5.700000 8.805000 5.870000 ;
      RECT 1.695000 0.440000 1.865000 5.530000 ;
      RECT 2.475000 0.440000 2.645000 5.530000 ;
      RECT 3.255000 0.440000 3.425000 5.530000 ;
      RECT 4.035000 0.440000 4.205000 5.530000 ;
      RECT 4.815000 0.440000 4.985000 5.530000 ;
      RECT 5.595000 0.440000 5.765000 5.530000 ;
      RECT 6.375000 0.440000 6.545000 5.530000 ;
      RECT 7.155000 0.440000 7.325000 5.530000 ;
      RECT 7.935000 0.440000 8.105000 5.530000 ;
      RECT 8.715000 0.440000 8.885000 5.530000 ;
      RECT 9.390000 0.560000 9.560000 5.410000 ;
    LAYER mcon ;
      RECT 0.240000 0.920000 0.410000 1.090000 ;
      RECT 0.240000 1.280000 0.410000 1.450000 ;
      RECT 0.240000 1.640000 0.410000 1.810000 ;
      RECT 0.240000 2.000000 0.410000 2.170000 ;
      RECT 0.240000 2.360000 0.410000 2.530000 ;
      RECT 0.240000 2.720000 0.410000 2.890000 ;
      RECT 0.240000 3.080000 0.410000 3.250000 ;
      RECT 0.240000 3.440000 0.410000 3.610000 ;
      RECT 0.240000 3.800000 0.410000 3.970000 ;
      RECT 0.240000 4.160000 0.410000 4.330000 ;
      RECT 0.240000 4.520000 0.410000 4.690000 ;
      RECT 0.240000 4.880000 0.410000 5.050000 ;
      RECT 0.240000 5.240000 0.410000 5.410000 ;
      RECT 0.915000 0.560000 1.085000 0.730000 ;
      RECT 0.915000 0.920000 1.085000 1.090000 ;
      RECT 0.915000 1.280000 1.085000 1.450000 ;
      RECT 0.915000 1.640000 1.085000 1.810000 ;
      RECT 0.915000 2.000000 1.085000 2.170000 ;
      RECT 0.915000 2.360000 1.085000 2.530000 ;
      RECT 0.915000 2.720000 1.085000 2.890000 ;
      RECT 0.915000 3.080000 1.085000 3.250000 ;
      RECT 0.915000 3.440000 1.085000 3.610000 ;
      RECT 0.915000 3.800000 1.085000 3.970000 ;
      RECT 0.915000 4.160000 1.085000 4.330000 ;
      RECT 0.915000 4.520000 1.085000 4.690000 ;
      RECT 0.915000 4.880000 1.085000 5.050000 ;
      RECT 0.915000 5.240000 1.085000 5.410000 ;
      RECT 1.035000 0.100000 1.205000 0.270000 ;
      RECT 1.035000 5.700000 1.205000 5.870000 ;
      RECT 1.395000 0.100000 1.565000 0.270000 ;
      RECT 1.395000 5.700000 1.565000 5.870000 ;
      RECT 1.695000 0.560000 1.865000 0.730000 ;
      RECT 1.695000 0.920000 1.865000 1.090000 ;
      RECT 1.695000 1.280000 1.865000 1.450000 ;
      RECT 1.695000 1.640000 1.865000 1.810000 ;
      RECT 1.695000 2.000000 1.865000 2.170000 ;
      RECT 1.695000 2.360000 1.865000 2.530000 ;
      RECT 1.695000 2.720000 1.865000 2.890000 ;
      RECT 1.695000 3.080000 1.865000 3.250000 ;
      RECT 1.695000 3.440000 1.865000 3.610000 ;
      RECT 1.695000 3.800000 1.865000 3.970000 ;
      RECT 1.695000 4.160000 1.865000 4.330000 ;
      RECT 1.695000 4.520000 1.865000 4.690000 ;
      RECT 1.695000 4.880000 1.865000 5.050000 ;
      RECT 1.695000 5.240000 1.865000 5.410000 ;
      RECT 1.755000 0.100000 1.925000 0.270000 ;
      RECT 1.755000 5.700000 1.925000 5.870000 ;
      RECT 2.115000 0.100000 2.285000 0.270000 ;
      RECT 2.115000 5.700000 2.285000 5.870000 ;
      RECT 2.475000 0.100000 2.645000 0.270000 ;
      RECT 2.475000 0.560000 2.645000 0.730000 ;
      RECT 2.475000 0.920000 2.645000 1.090000 ;
      RECT 2.475000 1.280000 2.645000 1.450000 ;
      RECT 2.475000 1.640000 2.645000 1.810000 ;
      RECT 2.475000 2.000000 2.645000 2.170000 ;
      RECT 2.475000 2.360000 2.645000 2.530000 ;
      RECT 2.475000 2.720000 2.645000 2.890000 ;
      RECT 2.475000 3.080000 2.645000 3.250000 ;
      RECT 2.475000 3.440000 2.645000 3.610000 ;
      RECT 2.475000 3.800000 2.645000 3.970000 ;
      RECT 2.475000 4.160000 2.645000 4.330000 ;
      RECT 2.475000 4.520000 2.645000 4.690000 ;
      RECT 2.475000 4.880000 2.645000 5.050000 ;
      RECT 2.475000 5.240000 2.645000 5.410000 ;
      RECT 2.475000 5.700000 2.645000 5.870000 ;
      RECT 2.835000 0.100000 3.005000 0.270000 ;
      RECT 2.835000 5.700000 3.005000 5.870000 ;
      RECT 3.195000 0.100000 3.365000 0.270000 ;
      RECT 3.195000 5.700000 3.365000 5.870000 ;
      RECT 3.255000 0.560000 3.425000 0.730000 ;
      RECT 3.255000 0.920000 3.425000 1.090000 ;
      RECT 3.255000 1.280000 3.425000 1.450000 ;
      RECT 3.255000 1.640000 3.425000 1.810000 ;
      RECT 3.255000 2.000000 3.425000 2.170000 ;
      RECT 3.255000 2.360000 3.425000 2.530000 ;
      RECT 3.255000 2.720000 3.425000 2.890000 ;
      RECT 3.255000 3.080000 3.425000 3.250000 ;
      RECT 3.255000 3.440000 3.425000 3.610000 ;
      RECT 3.255000 3.800000 3.425000 3.970000 ;
      RECT 3.255000 4.160000 3.425000 4.330000 ;
      RECT 3.255000 4.520000 3.425000 4.690000 ;
      RECT 3.255000 4.880000 3.425000 5.050000 ;
      RECT 3.255000 5.240000 3.425000 5.410000 ;
      RECT 3.555000 0.100000 3.725000 0.270000 ;
      RECT 3.555000 5.700000 3.725000 5.870000 ;
      RECT 3.915000 0.100000 4.085000 0.270000 ;
      RECT 3.915000 5.700000 4.085000 5.870000 ;
      RECT 4.035000 0.560000 4.205000 0.730000 ;
      RECT 4.035000 0.920000 4.205000 1.090000 ;
      RECT 4.035000 1.280000 4.205000 1.450000 ;
      RECT 4.035000 1.640000 4.205000 1.810000 ;
      RECT 4.035000 2.000000 4.205000 2.170000 ;
      RECT 4.035000 2.360000 4.205000 2.530000 ;
      RECT 4.035000 2.720000 4.205000 2.890000 ;
      RECT 4.035000 3.080000 4.205000 3.250000 ;
      RECT 4.035000 3.440000 4.205000 3.610000 ;
      RECT 4.035000 3.800000 4.205000 3.970000 ;
      RECT 4.035000 4.160000 4.205000 4.330000 ;
      RECT 4.035000 4.520000 4.205000 4.690000 ;
      RECT 4.035000 4.880000 4.205000 5.050000 ;
      RECT 4.035000 5.240000 4.205000 5.410000 ;
      RECT 4.275000 0.100000 4.445000 0.270000 ;
      RECT 4.275000 5.700000 4.445000 5.870000 ;
      RECT 4.635000 0.100000 4.805000 0.270000 ;
      RECT 4.635000 5.700000 4.805000 5.870000 ;
      RECT 4.815000 0.560000 4.985000 0.730000 ;
      RECT 4.815000 0.920000 4.985000 1.090000 ;
      RECT 4.815000 1.280000 4.985000 1.450000 ;
      RECT 4.815000 1.640000 4.985000 1.810000 ;
      RECT 4.815000 2.000000 4.985000 2.170000 ;
      RECT 4.815000 2.360000 4.985000 2.530000 ;
      RECT 4.815000 2.720000 4.985000 2.890000 ;
      RECT 4.815000 3.080000 4.985000 3.250000 ;
      RECT 4.815000 3.440000 4.985000 3.610000 ;
      RECT 4.815000 3.800000 4.985000 3.970000 ;
      RECT 4.815000 4.160000 4.985000 4.330000 ;
      RECT 4.815000 4.520000 4.985000 4.690000 ;
      RECT 4.815000 4.880000 4.985000 5.050000 ;
      RECT 4.815000 5.240000 4.985000 5.410000 ;
      RECT 4.995000 0.100000 5.165000 0.270000 ;
      RECT 4.995000 5.700000 5.165000 5.870000 ;
      RECT 5.355000 0.100000 5.525000 0.270000 ;
      RECT 5.355000 5.700000 5.525000 5.870000 ;
      RECT 5.595000 0.560000 5.765000 0.730000 ;
      RECT 5.595000 0.920000 5.765000 1.090000 ;
      RECT 5.595000 1.280000 5.765000 1.450000 ;
      RECT 5.595000 1.640000 5.765000 1.810000 ;
      RECT 5.595000 2.000000 5.765000 2.170000 ;
      RECT 5.595000 2.360000 5.765000 2.530000 ;
      RECT 5.595000 2.720000 5.765000 2.890000 ;
      RECT 5.595000 3.080000 5.765000 3.250000 ;
      RECT 5.595000 3.440000 5.765000 3.610000 ;
      RECT 5.595000 3.800000 5.765000 3.970000 ;
      RECT 5.595000 4.160000 5.765000 4.330000 ;
      RECT 5.595000 4.520000 5.765000 4.690000 ;
      RECT 5.595000 4.880000 5.765000 5.050000 ;
      RECT 5.595000 5.240000 5.765000 5.410000 ;
      RECT 5.715000 0.100000 5.885000 0.270000 ;
      RECT 5.715000 5.700000 5.885000 5.870000 ;
      RECT 6.075000 0.100000 6.245000 0.270000 ;
      RECT 6.075000 5.700000 6.245000 5.870000 ;
      RECT 6.375000 0.560000 6.545000 0.730000 ;
      RECT 6.375000 0.920000 6.545000 1.090000 ;
      RECT 6.375000 1.280000 6.545000 1.450000 ;
      RECT 6.375000 1.640000 6.545000 1.810000 ;
      RECT 6.375000 2.000000 6.545000 2.170000 ;
      RECT 6.375000 2.360000 6.545000 2.530000 ;
      RECT 6.375000 2.720000 6.545000 2.890000 ;
      RECT 6.375000 3.080000 6.545000 3.250000 ;
      RECT 6.375000 3.440000 6.545000 3.610000 ;
      RECT 6.375000 3.800000 6.545000 3.970000 ;
      RECT 6.375000 4.160000 6.545000 4.330000 ;
      RECT 6.375000 4.520000 6.545000 4.690000 ;
      RECT 6.375000 4.880000 6.545000 5.050000 ;
      RECT 6.375000 5.240000 6.545000 5.410000 ;
      RECT 6.435000 0.100000 6.605000 0.270000 ;
      RECT 6.435000 5.700000 6.605000 5.870000 ;
      RECT 6.795000 0.100000 6.965000 0.270000 ;
      RECT 6.795000 5.700000 6.965000 5.870000 ;
      RECT 7.155000 0.100000 7.325000 0.270000 ;
      RECT 7.155000 0.560000 7.325000 0.730000 ;
      RECT 7.155000 0.920000 7.325000 1.090000 ;
      RECT 7.155000 1.280000 7.325000 1.450000 ;
      RECT 7.155000 1.640000 7.325000 1.810000 ;
      RECT 7.155000 2.000000 7.325000 2.170000 ;
      RECT 7.155000 2.360000 7.325000 2.530000 ;
      RECT 7.155000 2.720000 7.325000 2.890000 ;
      RECT 7.155000 3.080000 7.325000 3.250000 ;
      RECT 7.155000 3.440000 7.325000 3.610000 ;
      RECT 7.155000 3.800000 7.325000 3.970000 ;
      RECT 7.155000 4.160000 7.325000 4.330000 ;
      RECT 7.155000 4.520000 7.325000 4.690000 ;
      RECT 7.155000 4.880000 7.325000 5.050000 ;
      RECT 7.155000 5.240000 7.325000 5.410000 ;
      RECT 7.155000 5.700000 7.325000 5.870000 ;
      RECT 7.515000 0.100000 7.685000 0.270000 ;
      RECT 7.515000 5.700000 7.685000 5.870000 ;
      RECT 7.875000 0.100000 8.045000 0.270000 ;
      RECT 7.875000 5.700000 8.045000 5.870000 ;
      RECT 7.935000 0.560000 8.105000 0.730000 ;
      RECT 7.935000 0.920000 8.105000 1.090000 ;
      RECT 7.935000 1.280000 8.105000 1.450000 ;
      RECT 7.935000 1.640000 8.105000 1.810000 ;
      RECT 7.935000 2.000000 8.105000 2.170000 ;
      RECT 7.935000 2.360000 8.105000 2.530000 ;
      RECT 7.935000 2.720000 8.105000 2.890000 ;
      RECT 7.935000 3.080000 8.105000 3.250000 ;
      RECT 7.935000 3.440000 8.105000 3.610000 ;
      RECT 7.935000 3.800000 8.105000 3.970000 ;
      RECT 7.935000 4.160000 8.105000 4.330000 ;
      RECT 7.935000 4.520000 8.105000 4.690000 ;
      RECT 7.935000 4.880000 8.105000 5.050000 ;
      RECT 7.935000 5.240000 8.105000 5.410000 ;
      RECT 8.235000 0.100000 8.405000 0.270000 ;
      RECT 8.235000 5.700000 8.405000 5.870000 ;
      RECT 8.595000 0.100000 8.765000 0.270000 ;
      RECT 8.595000 5.700000 8.765000 5.870000 ;
      RECT 8.715000 0.560000 8.885000 0.730000 ;
      RECT 8.715000 0.920000 8.885000 1.090000 ;
      RECT 8.715000 1.280000 8.885000 1.450000 ;
      RECT 8.715000 1.640000 8.885000 1.810000 ;
      RECT 8.715000 2.000000 8.885000 2.170000 ;
      RECT 8.715000 2.360000 8.885000 2.530000 ;
      RECT 8.715000 2.720000 8.885000 2.890000 ;
      RECT 8.715000 3.080000 8.885000 3.250000 ;
      RECT 8.715000 3.440000 8.885000 3.610000 ;
      RECT 8.715000 3.800000 8.885000 3.970000 ;
      RECT 8.715000 4.160000 8.885000 4.330000 ;
      RECT 8.715000 4.520000 8.885000 4.690000 ;
      RECT 8.715000 4.880000 8.885000 5.050000 ;
      RECT 8.715000 5.240000 8.885000 5.410000 ;
      RECT 9.390000 0.920000 9.560000 1.090000 ;
      RECT 9.390000 1.280000 9.560000 1.450000 ;
      RECT 9.390000 1.640000 9.560000 1.810000 ;
      RECT 9.390000 2.000000 9.560000 2.170000 ;
      RECT 9.390000 2.360000 9.560000 2.530000 ;
      RECT 9.390000 2.720000 9.560000 2.890000 ;
      RECT 9.390000 3.080000 9.560000 3.250000 ;
      RECT 9.390000 3.440000 9.560000 3.610000 ;
      RECT 9.390000 3.800000 9.560000 3.970000 ;
      RECT 9.390000 4.160000 9.560000 4.330000 ;
      RECT 9.390000 4.520000 9.560000 4.690000 ;
      RECT 9.390000 4.880000 9.560000 5.050000 ;
      RECT 9.390000 5.240000 9.560000 5.410000 ;
    LAYER met1 ;
      RECT 0.870000 0.500000 1.130000 5.470000 ;
      RECT 1.650000 0.500000 1.910000 5.470000 ;
      RECT 2.430000 0.500000 2.690000 5.470000 ;
      RECT 3.210000 0.500000 3.470000 5.470000 ;
      RECT 3.990000 0.500000 4.250000 5.470000 ;
      RECT 4.770000 0.500000 5.030000 5.470000 ;
      RECT 5.550000 0.500000 5.810000 5.470000 ;
      RECT 6.330000 0.500000 6.590000 5.470000 ;
      RECT 7.110000 0.500000 7.370000 5.470000 ;
      RECT 7.890000 0.500000 8.150000 5.470000 ;
      RECT 8.670000 0.500000 8.930000 5.470000 ;
    LAYER via ;
      RECT 0.870000 0.530000 1.130000 0.790000 ;
      RECT 0.870000 0.850000 1.130000 1.110000 ;
      RECT 0.870000 1.170000 1.130000 1.430000 ;
      RECT 0.870000 1.490000 1.130000 1.750000 ;
      RECT 0.870000 1.810000 1.130000 2.070000 ;
      RECT 0.870000 2.130000 1.130000 2.390000 ;
      RECT 0.870000 2.450000 1.130000 2.710000 ;
      RECT 1.650000 3.260000 1.910000 3.520000 ;
      RECT 1.650000 3.580000 1.910000 3.840000 ;
      RECT 1.650000 3.900000 1.910000 4.160000 ;
      RECT 1.650000 4.220000 1.910000 4.480000 ;
      RECT 1.650000 4.540000 1.910000 4.800000 ;
      RECT 1.650000 4.860000 1.910000 5.120000 ;
      RECT 1.650000 5.180000 1.910000 5.440000 ;
      RECT 2.430000 0.530000 2.690000 0.790000 ;
      RECT 2.430000 0.850000 2.690000 1.110000 ;
      RECT 2.430000 1.170000 2.690000 1.430000 ;
      RECT 2.430000 1.490000 2.690000 1.750000 ;
      RECT 2.430000 1.810000 2.690000 2.070000 ;
      RECT 2.430000 2.130000 2.690000 2.390000 ;
      RECT 2.430000 2.450000 2.690000 2.710000 ;
      RECT 3.210000 3.260000 3.470000 3.520000 ;
      RECT 3.210000 3.580000 3.470000 3.840000 ;
      RECT 3.210000 3.900000 3.470000 4.160000 ;
      RECT 3.210000 4.220000 3.470000 4.480000 ;
      RECT 3.210000 4.540000 3.470000 4.800000 ;
      RECT 3.210000 4.860000 3.470000 5.120000 ;
      RECT 3.210000 5.180000 3.470000 5.440000 ;
      RECT 3.990000 0.530000 4.250000 0.790000 ;
      RECT 3.990000 0.850000 4.250000 1.110000 ;
      RECT 3.990000 1.170000 4.250000 1.430000 ;
      RECT 3.990000 1.490000 4.250000 1.750000 ;
      RECT 3.990000 1.810000 4.250000 2.070000 ;
      RECT 3.990000 2.130000 4.250000 2.390000 ;
      RECT 3.990000 2.450000 4.250000 2.710000 ;
      RECT 4.770000 3.260000 5.030000 3.520000 ;
      RECT 4.770000 3.580000 5.030000 3.840000 ;
      RECT 4.770000 3.900000 5.030000 4.160000 ;
      RECT 4.770000 4.220000 5.030000 4.480000 ;
      RECT 4.770000 4.540000 5.030000 4.800000 ;
      RECT 4.770000 4.860000 5.030000 5.120000 ;
      RECT 4.770000 5.180000 5.030000 5.440000 ;
      RECT 5.550000 0.530000 5.810000 0.790000 ;
      RECT 5.550000 0.850000 5.810000 1.110000 ;
      RECT 5.550000 1.170000 5.810000 1.430000 ;
      RECT 5.550000 1.490000 5.810000 1.750000 ;
      RECT 5.550000 1.810000 5.810000 2.070000 ;
      RECT 5.550000 2.130000 5.810000 2.390000 ;
      RECT 5.550000 2.450000 5.810000 2.710000 ;
      RECT 6.330000 3.260000 6.590000 3.520000 ;
      RECT 6.330000 3.580000 6.590000 3.840000 ;
      RECT 6.330000 3.900000 6.590000 4.160000 ;
      RECT 6.330000 4.220000 6.590000 4.480000 ;
      RECT 6.330000 4.540000 6.590000 4.800000 ;
      RECT 6.330000 4.860000 6.590000 5.120000 ;
      RECT 6.330000 5.180000 6.590000 5.440000 ;
      RECT 7.110000 0.530000 7.370000 0.790000 ;
      RECT 7.110000 0.850000 7.370000 1.110000 ;
      RECT 7.110000 1.170000 7.370000 1.430000 ;
      RECT 7.110000 1.490000 7.370000 1.750000 ;
      RECT 7.110000 1.810000 7.370000 2.070000 ;
      RECT 7.110000 2.130000 7.370000 2.390000 ;
      RECT 7.110000 2.450000 7.370000 2.710000 ;
      RECT 7.890000 3.260000 8.150000 3.520000 ;
      RECT 7.890000 3.580000 8.150000 3.840000 ;
      RECT 7.890000 3.900000 8.150000 4.160000 ;
      RECT 7.890000 4.220000 8.150000 4.480000 ;
      RECT 7.890000 4.540000 8.150000 4.800000 ;
      RECT 7.890000 4.860000 8.150000 5.120000 ;
      RECT 7.890000 5.180000 8.150000 5.440000 ;
      RECT 8.670000 0.530000 8.930000 0.790000 ;
      RECT 8.670000 0.850000 8.930000 1.110000 ;
      RECT 8.670000 1.170000 8.930000 1.430000 ;
      RECT 8.670000 1.490000 8.930000 1.750000 ;
      RECT 8.670000 1.810000 8.930000 2.070000 ;
      RECT 8.670000 2.130000 8.930000 2.390000 ;
      RECT 8.670000 2.450000 8.930000 2.710000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50
END LIBRARY
