# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_aura_blocking
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_aura_blocking ;
  ORIGIN  0.000000  213.9700 ;
  SIZE  1555.530 BY  412.1700 ;
  PIN B_P
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 -205.320000 11.985000 -202.345000 ;
    END
  END B_P
  PIN D_N2
    ANTENNADIFFAREA  3.360000 ;
    PORT
      LAYER met3 ;
        RECT 102.420000 102.075000 102.750000 102.515000 ;
        RECT 102.420000 102.515000 109.180000 102.845000 ;
        RECT 103.280000 102.075000 103.610000 102.515000 ;
        RECT 104.140000 102.075000 104.470000 102.515000 ;
        RECT 105.000000 102.075000 109.180000 102.515000 ;
    END
  END D_N2
  PIN D_P
    ANTENNADIFFAREA  0.235200 ;
    PORT
      LAYER met2 ;
        RECT 68.470000 -125.230000 68.730000 -124.590000 ;
    END
  END D_P
  PIN D_P2
    ANTENNADIFFAREA  0.840000 ;
    PORT
      LAYER met2 ;
        RECT 100.600000 -123.070000 103.420000 -122.430000 ;
    END
  END D_P2
  PIN G
    ANTENNAGATEAREA  0.126000 ;
    PORT
      LAYER met1 ;
        RECT 69.265000 100.485000 69.915000 100.775000 ;
    END
  END G
  PIN G_N2
    ANTENNAGATEAREA  3.600000 ;
    PORT
      LAYER met1 ;
        RECT 102.470000 103.065000 105.280000 111.830000 ;
    END
  END G_N2
  PIN G_P
    ANTENNAGATEAREA  0.252000 ;
    PORT
      LAYER met1 ;
        RECT 68.275000 -124.305000 68.925000 -124.015000 ;
    END
  END G_P
  PIN G_P2
    ANTENNAGATEAREA  0.900000 ;
    PORT
      LAYER met1 ;
        RECT 102.965000 -122.145000 103.615000 -120.555000 ;
    END
  END G_P2
  PIN NWELL
    ANTENNADIFFAREA  43.51075 ;
    PORT
      LAYER li1 ;
        RECT 9.175000 8.650000 11.985000 11.625000 ;
    END
  END NWELL
  PIN S
    ANTENNADIFFAREA  0.235200 ;
    PORT
      LAYER met1 ;
        RECT 69.045000 99.265000 70.135000  99.565000 ;
        RECT 69.045000 99.565000 69.275000 100.310000 ;
        RECT 69.905000 99.565000 70.135000 100.310000 ;
    END
  END S
  PIN S_N2
    ANTENNADIFFAREA  4.200000 ;
    PORT
      LAYER met1 ;
        RECT 102.040000 88.255000 105.710000  99.565000 ;
        RECT 102.040000 99.565000 102.270000 102.815000 ;
        RECT 102.900000 99.565000 103.130000 102.815000 ;
        RECT 103.760000 99.565000 103.990000 102.815000 ;
        RECT 104.620000 99.565000 104.850000 102.815000 ;
        RECT 105.480000 99.565000 105.710000 102.815000 ;
    END
  END S_N2
  PIN S_P
    ANTENNADIFFAREA  0.445200 ;
    PORT
      LAYER met1 ;
        RECT 68.055000 -125.955000 69.145000 -125.655000 ;
        RECT 68.055000 -125.655000 68.285000 -124.565000 ;
        RECT 68.915000 -125.655000 69.145000 -124.565000 ;
    END
  END S_P
  PIN S_P2
    ANTENNADIFFAREA  1.590000 ;
    PORT
      LAYER met1 ;
        RECT 102.745000 -127.045000 103.835000 -125.655000 ;
        RECT 102.745000 -125.655000 102.975000 -122.405000 ;
        RECT 103.605000 -125.655000 103.835000 -122.405000 ;
    END
  END S_P2
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 60.140000 90.690000 62.950000 93.665000 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 69.460000 99.965000 69.720000 100.310000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  68.085000 -125.255000  68.255000 -124.565000 ;
      RECT  68.265000 -124.335000  68.935000 -123.995000 ;
      RECT  68.515000 -125.255000  68.685000 -124.565000 ;
      RECT  68.945000 -125.255000  69.115000 -124.565000 ;
      RECT  69.075000   99.965000  69.245000  100.295000 ;
      RECT  69.255000  100.465000  69.925000  100.795000 ;
      RECT  69.505000   99.965000  69.675000  100.295000 ;
      RECT  69.935000   99.965000  70.105000  100.295000 ;
      RECT 102.070000   99.965000 102.240000  102.815000 ;
      RECT 102.500000   99.965000 102.670000  102.815000 ;
      RECT 102.520000  103.045000 105.230000  103.375000 ;
      RECT 102.775000 -125.275000 102.945000 -122.405000 ;
      RECT 102.930000   99.965000 103.100000  102.815000 ;
      RECT 102.955000 -122.175000 103.625000 -121.835000 ;
      RECT 103.205000 -125.255000 103.375000 -122.405000 ;
      RECT 103.360000   99.965000 103.530000  102.815000 ;
      RECT 103.635000 -125.255000 103.805000 -122.405000 ;
      RECT 103.790000   99.965000 103.960000  102.815000 ;
      RECT 104.220000   99.965000 104.390000  102.815000 ;
      RECT 104.650000   99.965000 104.820000  102.815000 ;
      RECT 105.080000   99.965000 105.250000  102.815000 ;
      RECT 105.510000   99.965000 105.680000  102.815000 ;
    LAYER mcon ;
      RECT  68.085000 -125.175000  68.255000 -125.005000 ;
      RECT  68.085000 -124.815000  68.255000 -124.645000 ;
      RECT  68.335000 -124.245000  68.505000 -124.075000 ;
      RECT  68.515000 -125.175000  68.685000 -125.005000 ;
      RECT  68.515000 -124.815000  68.685000 -124.645000 ;
      RECT  68.695000 -124.245000  68.865000 -124.075000 ;
      RECT  68.945000 -125.175000  69.115000 -125.005000 ;
      RECT  68.945000 -124.815000  69.115000 -124.645000 ;
      RECT  69.075000  100.045000  69.245000  100.215000 ;
      RECT  69.325000  100.545000  69.495000  100.715000 ;
      RECT  69.505000  100.045000  69.675000  100.215000 ;
      RECT  69.685000  100.545000  69.855000  100.715000 ;
      RECT  69.935000  100.045000  70.105000  100.215000 ;
      RECT 102.070000  100.045000 102.240000  100.215000 ;
      RECT 102.070000  100.405000 102.240000  100.575000 ;
      RECT 102.070000  100.765000 102.240000  100.935000 ;
      RECT 102.070000  101.125000 102.240000  101.295000 ;
      RECT 102.070000  101.485000 102.240000  101.655000 ;
      RECT 102.070000  101.845000 102.240000  102.015000 ;
      RECT 102.070000  102.205000 102.240000  102.375000 ;
      RECT 102.070000  102.565000 102.240000  102.735000 ;
      RECT 102.500000  100.045000 102.670000  100.215000 ;
      RECT 102.500000  100.405000 102.670000  100.575000 ;
      RECT 102.500000  100.765000 102.670000  100.935000 ;
      RECT 102.500000  101.125000 102.670000  101.295000 ;
      RECT 102.500000  101.485000 102.670000  101.655000 ;
      RECT 102.500000  101.845000 102.670000  102.015000 ;
      RECT 102.500000  102.205000 102.670000  102.375000 ;
      RECT 102.500000  102.565000 102.670000  102.735000 ;
      RECT 102.530000  103.125000 102.700000  103.295000 ;
      RECT 102.775000 -125.175000 102.945000 -125.005000 ;
      RECT 102.775000 -124.815000 102.945000 -124.645000 ;
      RECT 102.775000 -124.455000 102.945000 -124.285000 ;
      RECT 102.775000 -124.095000 102.945000 -123.925000 ;
      RECT 102.775000 -123.735000 102.945000 -123.565000 ;
      RECT 102.775000 -123.375000 102.945000 -123.205000 ;
      RECT 102.775000 -123.015000 102.945000 -122.845000 ;
      RECT 102.775000 -122.655000 102.945000 -122.485000 ;
      RECT 102.890000  103.125000 103.060000  103.295000 ;
      RECT 102.930000  100.045000 103.100000  100.215000 ;
      RECT 102.930000  100.405000 103.100000  100.575000 ;
      RECT 102.930000  100.765000 103.100000  100.935000 ;
      RECT 102.930000  101.125000 103.100000  101.295000 ;
      RECT 102.930000  101.485000 103.100000  101.655000 ;
      RECT 102.930000  101.845000 103.100000  102.015000 ;
      RECT 102.930000  102.205000 103.100000  102.375000 ;
      RECT 102.930000  102.565000 103.100000  102.735000 ;
      RECT 103.025000 -122.085000 103.195000 -121.915000 ;
      RECT 103.205000 -125.175000 103.375000 -125.005000 ;
      RECT 103.205000 -124.815000 103.375000 -124.645000 ;
      RECT 103.205000 -124.455000 103.375000 -124.285000 ;
      RECT 103.205000 -124.095000 103.375000 -123.925000 ;
      RECT 103.205000 -123.735000 103.375000 -123.565000 ;
      RECT 103.205000 -123.375000 103.375000 -123.205000 ;
      RECT 103.205000 -123.015000 103.375000 -122.845000 ;
      RECT 103.205000 -122.655000 103.375000 -122.485000 ;
      RECT 103.250000  103.125000 103.420000  103.295000 ;
      RECT 103.360000  100.045000 103.530000  100.215000 ;
      RECT 103.360000  100.405000 103.530000  100.575000 ;
      RECT 103.360000  100.765000 103.530000  100.935000 ;
      RECT 103.360000  101.125000 103.530000  101.295000 ;
      RECT 103.360000  101.485000 103.530000  101.655000 ;
      RECT 103.360000  101.845000 103.530000  102.015000 ;
      RECT 103.360000  102.205000 103.530000  102.375000 ;
      RECT 103.360000  102.565000 103.530000  102.735000 ;
      RECT 103.385000 -122.085000 103.555000 -121.915000 ;
      RECT 103.610000  103.125000 103.780000  103.295000 ;
      RECT 103.635000 -125.175000 103.805000 -125.005000 ;
      RECT 103.635000 -124.815000 103.805000 -124.645000 ;
      RECT 103.635000 -124.455000 103.805000 -124.285000 ;
      RECT 103.635000 -124.095000 103.805000 -123.925000 ;
      RECT 103.635000 -123.735000 103.805000 -123.565000 ;
      RECT 103.635000 -123.375000 103.805000 -123.205000 ;
      RECT 103.635000 -123.015000 103.805000 -122.845000 ;
      RECT 103.635000 -122.655000 103.805000 -122.485000 ;
      RECT 103.790000  100.045000 103.960000  100.215000 ;
      RECT 103.790000  100.405000 103.960000  100.575000 ;
      RECT 103.790000  100.765000 103.960000  100.935000 ;
      RECT 103.790000  101.125000 103.960000  101.295000 ;
      RECT 103.790000  101.485000 103.960000  101.655000 ;
      RECT 103.790000  101.845000 103.960000  102.015000 ;
      RECT 103.790000  102.205000 103.960000  102.375000 ;
      RECT 103.790000  102.565000 103.960000  102.735000 ;
      RECT 103.970000  103.125000 104.140000  103.295000 ;
      RECT 104.220000  100.045000 104.390000  100.215000 ;
      RECT 104.220000  100.405000 104.390000  100.575000 ;
      RECT 104.220000  100.765000 104.390000  100.935000 ;
      RECT 104.220000  101.125000 104.390000  101.295000 ;
      RECT 104.220000  101.485000 104.390000  101.655000 ;
      RECT 104.220000  101.845000 104.390000  102.015000 ;
      RECT 104.220000  102.205000 104.390000  102.375000 ;
      RECT 104.220000  102.565000 104.390000  102.735000 ;
      RECT 104.330000  103.125000 104.500000  103.295000 ;
      RECT 104.650000  100.045000 104.820000  100.215000 ;
      RECT 104.650000  100.405000 104.820000  100.575000 ;
      RECT 104.650000  100.765000 104.820000  100.935000 ;
      RECT 104.650000  101.125000 104.820000  101.295000 ;
      RECT 104.650000  101.485000 104.820000  101.655000 ;
      RECT 104.650000  101.845000 104.820000  102.015000 ;
      RECT 104.650000  102.205000 104.820000  102.375000 ;
      RECT 104.650000  102.565000 104.820000  102.735000 ;
      RECT 104.690000  103.125000 104.860000  103.295000 ;
      RECT 105.050000  103.125000 105.220000  103.295000 ;
      RECT 105.080000  100.045000 105.250000  100.215000 ;
      RECT 105.080000  100.405000 105.250000  100.575000 ;
      RECT 105.080000  100.765000 105.250000  100.935000 ;
      RECT 105.080000  101.125000 105.250000  101.295000 ;
      RECT 105.080000  101.485000 105.250000  101.655000 ;
      RECT 105.080000  101.845000 105.250000  102.015000 ;
      RECT 105.080000  102.205000 105.250000  102.375000 ;
      RECT 105.080000  102.565000 105.250000  102.735000 ;
      RECT 105.510000  100.045000 105.680000  100.215000 ;
      RECT 105.510000  100.405000 105.680000  100.575000 ;
      RECT 105.510000  100.765000 105.680000  100.935000 ;
      RECT 105.510000  101.125000 105.680000  101.295000 ;
      RECT 105.510000  101.485000 105.680000  101.655000 ;
      RECT 105.510000  101.845000 105.680000  102.015000 ;
      RECT 105.510000  102.205000 105.680000  102.375000 ;
      RECT 105.510000  102.565000 105.680000  102.735000 ;
    LAYER met1 ;
      RECT  68.470000 -125.255000  68.730000 -124.565000 ;
      RECT  69.460000   99.965000  69.720000  100.310000 ;
      RECT 102.455000   99.965000 102.715000  102.815000 ;
      RECT 103.160000 -125.255000 103.420000 -122.405000 ;
      RECT 103.315000   99.965000 103.575000  102.815000 ;
      RECT 104.175000   99.965000 104.435000  102.815000 ;
      RECT 105.035000   99.965000 105.295000  102.815000 ;
    LAYER met2 ;
      RECT 102.420000 102.075000 102.750000 102.845000 ;
      RECT 103.280000 102.075000 103.610000 102.845000 ;
      RECT 104.140000 102.075000 104.470000 102.845000 ;
      RECT 105.000000 102.075000 105.330000 102.845000 ;
    LAYER via ;
      RECT  68.470000 -125.200000  68.730000 -124.940000 ;
      RECT  68.470000 -124.880000  68.730000 -124.620000 ;
      RECT  69.460000  100.020000  69.720000  100.280000 ;
      RECT 102.455000  102.170000 102.715000  102.430000 ;
      RECT 102.455000  102.490000 102.715000  102.750000 ;
      RECT 103.160000 -123.040000 103.420000 -122.780000 ;
      RECT 103.160000 -122.720000 103.420000 -122.460000 ;
      RECT 103.315000  102.170000 103.575000  102.430000 ;
      RECT 103.315000  102.490000 103.575000  102.750000 ;
      RECT 104.175000  102.170000 104.435000  102.430000 ;
      RECT 104.175000  102.490000 104.435000  102.750000 ;
      RECT 105.035000  102.170000 105.295000  102.430000 ;
      RECT 105.035000  102.490000 105.295000  102.750000 ;
    LAYER via2 ;
      RECT 102.445000 102.120000 102.725000 102.400000 ;
      RECT 102.445000 102.520000 102.725000 102.800000 ;
      RECT 103.305000 102.120000 103.585000 102.400000 ;
      RECT 103.305000 102.520000 103.585000 102.800000 ;
      RECT 104.165000 102.120000 104.445000 102.400000 ;
      RECT 104.165000 102.520000 104.445000 102.800000 ;
      RECT 105.025000 102.120000 105.305000 102.400000 ;
      RECT 105.025000 102.520000 105.305000 102.800000 ;
  END
END sky130_fd_pr__rf_aura_blocking
END LIBRARY
