* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 49
.param
+ sky130_fd_pr__pfet_g5v0d10v5__toxe_mult = 0.958
+ sky130_fd_pr__pfet_g5v0d10v5__rshp_mult = 1.0
+ sky130_fd_pr__pfet_g5v0d10v5__overlap_mult = 0.7713
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = 9.5405e-1
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = 9.6374e-1
+ sky130_fd_pr__pfet_g5v0d10v5__lint_diff = 1.21275e-8
+ sky130_fd_pr__pfet_g5v0d10v5__wint_diff = -2.252e-8
+ sky130_fd_pr__pfet_g5v0d10v5__dlc_diff = 1.21275e-8
+ sky130_fd_pr__pfet_g5v0d10v5__dwc_diff = -2.252e-8
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 000, W = 10.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0 = -7.0417e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0 = -1.6969e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0 = 0.017499
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0 = 0.79042
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0 = -0.0014907
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0 = 0.01176
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0 = -2299.9
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 001, W = 15.0, L = 1.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1 = -2.4145e-20
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1 = 4.9447e-13
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1 = -0.01331
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1 = 0.0098739
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1 = 0.25894
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1 = -0.00028675
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1 = 0.010985
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1 = -0.021704
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 002, W = 15.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2 = -5.9283e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2 = -1.0976e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2 = 0.018416
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2 = 0.43209
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2 = -0.0013484
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2 = 0.020609
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2 = -1462.8
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 003, W = 1.5, L = 1.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3 = -0.044965
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3 = -2.763e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3 = -8.0117e-13
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3 = 0.016875
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3 = 0.0038857
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3 = 0.45247
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3 = -0.00043468
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3 = 0.030589
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 004, W = 1.5, L = 2.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4 = 0.49257
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4 = -0.0003094
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4 = 0.016822
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4 = -0.018182
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4 = -2.5531e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4 = -1.0749e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4 = 0.0041275
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4 = 0.0031794
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 005, W = 1.5, L = 4.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5 = 0.0052484
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5 = 0.58054
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5 = -0.0012815
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5 = 0.020192
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5 = 0.0086062
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5 = -4.572e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5 = -6.5592e-13
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5 = -0.0015263
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 006, W = 1.5, L = 0.5
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6 = 0.016254
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6 = 0.49885
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6 = -0.0025251
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6 = 0.047372
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6 = -6661.1
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6 = -1.0982e-18
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6 = -3.2409e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 007, W = 1.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7 = -0.0021467
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7 = 0.0084703
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7 = 0.030318
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7 = 0.43788
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7 = -0.00066807
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7 = -0.0030899
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7 = -3.5624e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7 = -1.2741e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 008, W = 1.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8 = -0.016142
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8 = 0.0067645
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8 = 0.030752
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8 = 0.4547
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8 = -0.00077831
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8 = -0.026222
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8 = -4.4393e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8 = -1.4493e-12
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 009, W = 1.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9 = 0.0029481
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9 = 0.0027432
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9 = 0.015539
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9 = 0.71845
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9 = -0.00042336
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9 = -0.014773
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9 = -2.0157e-19
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9 = -7.4139e-13
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 010, W = 1.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10 = 0.70361
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10 = -0.00042053
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10 = 0.022196
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10 = -0.0067387
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10 = 0.0036563
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10 = -5.2664e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10 = -1.3846e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10 = 0.00089972
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 011, W = 1.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11 = -14172.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11 = 0.64218
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11 = -0.00092434
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11 = 0.0053489
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11 = 0.016056
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11 = -6.2109e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11 = -3.4177e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 012, W = 1.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12 = -6394.2
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12 = 0.33479
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12 = -0.0022874
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12 = 0.042948
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12 = 0.0099952
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12 = -1.7117e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12 = -7.9172e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 013, W = 1.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13 = -6.2641e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13 = -2070.7
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13 = 0.24106
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13 = -0.0012391
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13 = 0.017619
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13 = 0.011885
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13 = -2.2611e-12
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 014, W = 20.0, L = 1.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14 = -2.2339e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14 = -3.4748e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14 = -0.0027677
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14 = 0.2613
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14 = -0.0010173
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14 = 0.0089301
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14 = -0.0046561
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14 = 0.0098286
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 015, W = 20.0, L = 0.5
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15 = 0.016758
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15 = -7.6331e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15 = -6.7478e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15 = -2345.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15 = 0.71112
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15 = -0.0017943
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15 = 0.0086003
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 016, W = 3.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16 = 0.023953
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16 = -0.0019796
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16 = 0.0096476
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16 = -4.2162e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16 = -6.0752e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16 = -0.0013042
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16 = 0.43547
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16 = -0.0019407
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 017, W = 3.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17 = 0.097301
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17 = -0.00011849
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17 = 0.0077129
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17 = -0.0022265
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17 = 0.0026014
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17 = 5.6809e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17 = 6.4174e-20
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17 = 0.00023435
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 018, W = 3.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18 = 0.98097
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18 = -0.0016199
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18 = 0.027082
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18 = -0.0013044
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18 = 0.0039521
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18 = -2.8525e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18 = -5.257e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18 = 0.00079995
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 019, W = 3.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19 = 0.69159
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19 = -0.00098827
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19 = 0.020715
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19 = 0.0027349
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19 = 0.001832
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19 = -6.8749e-14
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19 = -2.8016e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19 = -0.0005243
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 020, W = 3.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20 = 0.7433
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20 = -0.0010358
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20 = 0.0030566
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20 = 0.018187
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20 = -1.1077e-15
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20 = -3.469e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20 = -17641.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 021, W = 3.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21 = -5271.6
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21 = 0.42889
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21 = -0.0023822
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21 = 0.035099
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21 = 0.014984
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21 = -1.5233e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21 = -8.2984e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 022, W = 5.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22 = -0.011727
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22 = -0.022708
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22 = 0.22792
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22 = 0.00011294
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22 = -0.0065197
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22 = -0.019475
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22 = 0.0070962
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22 = 8.3705e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22 = 1.2248e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 023, W = 5.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23 = -0.0011748
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23 = -0.00064682
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23 = 0.0034225
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23 = 0.0069922
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23 = 0.0019484
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23 = 1.6171e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23 = -1.9654e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 024, W = 5.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24 = -5.9401e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24 = -7.8837e-5
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24 = 1.0085
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24 = -0.0020126
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24 = 0.022537
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24 = 0.0044239
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24 = 0.0045906
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24 = 1.9223e-13
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 025, W = 5.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25 = 1.7394e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25 = -4.7403e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25 = -0.0019895
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25 = 0.69602
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25 = -0.0016361
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25 = 0.02005
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25 = 0.011231
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25 = 0.0019101
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 026, W = 5.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26 = 0.014594
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26 = 1.8778e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26 = -4.0807e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26 = -3166.3
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26 = -0.0014253
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26 = 0.0029841
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 027, W = 5.0, L = 0.6
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27 = 0.0097998
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27 = 0.01485
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27 = -2.5143e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27 = -1.3084e-18
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27 = -1532.4
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27 = 0.39658
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27 = -0.0037304
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 028, W = 5.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28 = 0.26345
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28 = -0.0026196
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28 = 0.007018
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28 = 0.0081963
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28 = -1.4739e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28 = -9.7683e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28 = -1594.3
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 029, W = 7.0, L = 1.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29 = 0.41794
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29 = -0.0013974
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29 = 0.019167
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29 = -0.024678
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29 = 0.0098388
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29 = 1.5999e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29 = -3.925e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29 = -0.015175
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 030, W = 7.0, L = 2.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30 = 0.089816
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30 = -0.00060514
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30 = 0.0016094
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30 = 0.014146
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30 = 0.0023551
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30 = 2.0301e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30 = -1.7954e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30 = -0.0021302
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 031, W = 7.0, L = 4.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31 = 0.95786
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31 = -0.0019727
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31 = 0.021836
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31 = 0.015705
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31 = 0.0042542
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31 = 5.7956e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31 = -5.0534e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31 = -0.0026549
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 032, W = 7.0, L = 8.0
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32 = 0.68072
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32 = -0.0015217
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32 = 0.020982
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32 = 0.013747
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32 = 0.0019231
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32 = 3.8882e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32 = -4.1047e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32 = -0.0026026
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 033, W = 7.0, L = 0.5
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33 = -2670.2
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33 = 0.75873
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33 = -0.002097
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33 = 0.0039967
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33 = 0.017705
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33 = -8.0619e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33 = -7.3071e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 034, W = 7.0, L = 0.8
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34 = -1248.7
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34 = 0.28977
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34 = -0.0029381
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34 = 0.014786
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34 = 0.0087393
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34 = -6.1221e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34 = -9.5744e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 035, W = 0.42, L = 1.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35 = 6.7839e-20
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35 = -0.022763
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35 = 2.1877e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35 = -2.8156e-10
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35 = 0.35049
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35 = 0.0015076
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35 = 0.0056123
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35 = 0.0024959
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35 = -2.5118e-12
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 036, W = 0.42, L = 20.0
* --------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36 = -1.3292e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36 = 1.5957e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36 = 6.5479e-9
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36 = 1.0621e-8
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36 = 0.934
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36 = 0.00087945
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36 = 0.0086474
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36 = 0.0018058
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 037, W = 0.42, L = 2.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37 = -0.0010027
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37 = -2.3745e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37 = 2.8046e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37 = -0.040574
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37 = 3.8102e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37 = 6.352e-9
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37 = 0.27454
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37 = 0.0020631
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37 = 0.020372
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 038, W = 0.42, L = 4.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38 = 0.016159
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38 = 0.00074828
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38 = -1.5443e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38 = 2.6851e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38 = -0.037654
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38 = 4.723e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38 = 4.1672e-9
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38 = 0.22795
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38 = 0.0016924
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 039, W = 0.42, L = 8.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39 = 0.5609
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39 = 0.00064671
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39 = 0.027561
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39 = 0.0021797
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39 = -1.5173e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39 = 7.7269e-21
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39 = 3.7175e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39 = 9.268e-9
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 040, W = 0.42, L = 0.5
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40 = 0.50613
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40 = -0.0028309
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40 = 0.10585
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40 = 0.024914
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40 = -7.3558e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40 = -1.7838e-18
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40 = -12133.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 041, W = 0.42, L = 0.6
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41 = 0.0013149
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41 = 0.030622
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41 = 0.010608
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41 = -2.8842e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41 = -9.3118e-20
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41 = -6371.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 042, W = 0.42, L = 0.8
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42 = 0.61881
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42 = -2.936e-5
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42 = 0.056572
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42 = 0.011445
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42 = 4.9203e-15
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42 = -2.4879e-20
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42 = -3762.9
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 043, W = 0.75, L = 1.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43 = 1.6542e-7
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43 = 2.2364e-10
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43 = 0.3228
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43 = -0.00118
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43 = 0.027713
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43 = 0.0079579
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43 = -3.5343e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43 = -8.1028e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 044, W = 0.75, L = 2.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44 = 9.4635e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44 = 6.4018e-11
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44 = 0.38632
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44 = -0.0016524
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44 = 0.022555
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44 = 0.0084984
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44 = -3.2465e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44 = -9.0123e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44 = 0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 045, W = 0.75, L = 4.0
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45 = 6.3575e-8
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45 = 2.0655e-10
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45 = 0.68349
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45 = -0.00047153
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45 = 0.024269
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45 = 0.0051778
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45 = -9.9452e-13
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45 = -2.6577e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 046, W = 0.75, L = 0.5
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46 = -1.2351e-18
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46 = -6817.7
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46 = 0.44635
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46 = -0.0022504
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46 = 0.061329
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46 = 0.019348
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46 = -4.7537e-12
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 047, W = 0.75, L = 0.8
* -------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47 = -2.9185e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47 = -9.5406e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47 = -7552.8
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47 = 0.33372
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47 = -0.0021664
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47 = 0.028491
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47 = 0.01126
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 048, W = 0.7, L = 0.6
* ------------------------------
+ sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48 = 0.010007
+ sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48 = -1.83e-12
+ sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48 = -1.195e-19
+ sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48 = -5655.8
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48 = 0.00048052
+ sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48 = 0.0
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48 = 0.0044283
.include "sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"
