# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.500000 BY  5.970000 ;
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 3.110000 3.500000 5.470000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.636000 ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.100000 2.595000 0.270000 ;
        RECT 0.905000 5.700000 2.595000 5.870000 ;
      LAYER mcon ;
        RECT 0.945000 0.100000 1.115000 0.270000 ;
        RECT 0.945000 5.700000 1.115000 5.870000 ;
        RECT 1.305000 0.100000 1.475000 0.270000 ;
        RECT 1.305000 5.700000 1.475000 5.870000 ;
        RECT 1.665000 0.100000 1.835000 0.270000 ;
        RECT 1.665000 5.700000 1.835000 5.870000 ;
        RECT 2.025000 0.100000 2.195000 0.270000 ;
        RECT 2.025000 5.700000 2.195000 5.870000 ;
        RECT 2.385000 0.100000 2.555000 0.270000 ;
        RECT 2.385000 5.700000 2.555000 5.870000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.885000 0.000000 2.615000 0.330000 ;
        RECT 0.885000 5.640000 2.615000 5.970000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.500000 3.500000 2.860000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.464500 ;
    PORT
      LAYER met1 ;
        RECT 0.130000 0.500000 0.420000 5.470000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.080000 0.500000 3.370000 5.470000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.190000 0.560000 0.360000 5.410000 ;
      RECT 0.745000 0.440000 0.915000 5.530000 ;
      RECT 1.205000 0.440000 1.375000 5.530000 ;
      RECT 1.665000 0.440000 1.835000 5.530000 ;
      RECT 2.125000 0.440000 2.295000 5.530000 ;
      RECT 2.585000 0.440000 2.755000 5.530000 ;
      RECT 3.140000 0.560000 3.310000 5.410000 ;
    LAYER mcon ;
      RECT 0.190000 0.920000 0.360000 1.090000 ;
      RECT 0.190000 1.280000 0.360000 1.450000 ;
      RECT 0.190000 1.640000 0.360000 1.810000 ;
      RECT 0.190000 2.000000 0.360000 2.170000 ;
      RECT 0.190000 2.360000 0.360000 2.530000 ;
      RECT 0.190000 2.720000 0.360000 2.890000 ;
      RECT 0.190000 3.080000 0.360000 3.250000 ;
      RECT 0.190000 3.440000 0.360000 3.610000 ;
      RECT 0.190000 3.800000 0.360000 3.970000 ;
      RECT 0.190000 4.160000 0.360000 4.330000 ;
      RECT 0.190000 4.520000 0.360000 4.690000 ;
      RECT 0.190000 4.880000 0.360000 5.050000 ;
      RECT 0.190000 5.240000 0.360000 5.410000 ;
      RECT 0.745000 0.560000 0.915000 0.730000 ;
      RECT 0.745000 0.920000 0.915000 1.090000 ;
      RECT 0.745000 1.280000 0.915000 1.450000 ;
      RECT 0.745000 1.640000 0.915000 1.810000 ;
      RECT 0.745000 2.000000 0.915000 2.170000 ;
      RECT 0.745000 2.360000 0.915000 2.530000 ;
      RECT 0.745000 2.720000 0.915000 2.890000 ;
      RECT 0.745000 3.080000 0.915000 3.250000 ;
      RECT 0.745000 3.440000 0.915000 3.610000 ;
      RECT 0.745000 3.800000 0.915000 3.970000 ;
      RECT 0.745000 4.160000 0.915000 4.330000 ;
      RECT 0.745000 4.520000 0.915000 4.690000 ;
      RECT 0.745000 4.880000 0.915000 5.050000 ;
      RECT 0.745000 5.240000 0.915000 5.410000 ;
      RECT 1.205000 0.560000 1.375000 0.730000 ;
      RECT 1.205000 0.920000 1.375000 1.090000 ;
      RECT 1.205000 1.280000 1.375000 1.450000 ;
      RECT 1.205000 1.640000 1.375000 1.810000 ;
      RECT 1.205000 2.000000 1.375000 2.170000 ;
      RECT 1.205000 2.360000 1.375000 2.530000 ;
      RECT 1.205000 2.720000 1.375000 2.890000 ;
      RECT 1.205000 3.080000 1.375000 3.250000 ;
      RECT 1.205000 3.440000 1.375000 3.610000 ;
      RECT 1.205000 3.800000 1.375000 3.970000 ;
      RECT 1.205000 4.160000 1.375000 4.330000 ;
      RECT 1.205000 4.520000 1.375000 4.690000 ;
      RECT 1.205000 4.880000 1.375000 5.050000 ;
      RECT 1.205000 5.240000 1.375000 5.410000 ;
      RECT 1.665000 0.560000 1.835000 0.730000 ;
      RECT 1.665000 0.920000 1.835000 1.090000 ;
      RECT 1.665000 1.280000 1.835000 1.450000 ;
      RECT 1.665000 1.640000 1.835000 1.810000 ;
      RECT 1.665000 2.000000 1.835000 2.170000 ;
      RECT 1.665000 2.360000 1.835000 2.530000 ;
      RECT 1.665000 2.720000 1.835000 2.890000 ;
      RECT 1.665000 3.080000 1.835000 3.250000 ;
      RECT 1.665000 3.440000 1.835000 3.610000 ;
      RECT 1.665000 3.800000 1.835000 3.970000 ;
      RECT 1.665000 4.160000 1.835000 4.330000 ;
      RECT 1.665000 4.520000 1.835000 4.690000 ;
      RECT 1.665000 4.880000 1.835000 5.050000 ;
      RECT 1.665000 5.240000 1.835000 5.410000 ;
      RECT 2.125000 0.560000 2.295000 0.730000 ;
      RECT 2.125000 0.920000 2.295000 1.090000 ;
      RECT 2.125000 1.280000 2.295000 1.450000 ;
      RECT 2.125000 1.640000 2.295000 1.810000 ;
      RECT 2.125000 2.000000 2.295000 2.170000 ;
      RECT 2.125000 2.360000 2.295000 2.530000 ;
      RECT 2.125000 2.720000 2.295000 2.890000 ;
      RECT 2.125000 3.080000 2.295000 3.250000 ;
      RECT 2.125000 3.440000 2.295000 3.610000 ;
      RECT 2.125000 3.800000 2.295000 3.970000 ;
      RECT 2.125000 4.160000 2.295000 4.330000 ;
      RECT 2.125000 4.520000 2.295000 4.690000 ;
      RECT 2.125000 4.880000 2.295000 5.050000 ;
      RECT 2.125000 5.240000 2.295000 5.410000 ;
      RECT 2.585000 0.560000 2.755000 0.730000 ;
      RECT 2.585000 0.920000 2.755000 1.090000 ;
      RECT 2.585000 1.280000 2.755000 1.450000 ;
      RECT 2.585000 1.640000 2.755000 1.810000 ;
      RECT 2.585000 2.000000 2.755000 2.170000 ;
      RECT 2.585000 2.360000 2.755000 2.530000 ;
      RECT 2.585000 2.720000 2.755000 2.890000 ;
      RECT 2.585000 3.080000 2.755000 3.250000 ;
      RECT 2.585000 3.440000 2.755000 3.610000 ;
      RECT 2.585000 3.800000 2.755000 3.970000 ;
      RECT 2.585000 4.160000 2.755000 4.330000 ;
      RECT 2.585000 4.520000 2.755000 4.690000 ;
      RECT 2.585000 4.880000 2.755000 5.050000 ;
      RECT 2.585000 5.240000 2.755000 5.410000 ;
      RECT 3.140000 0.920000 3.310000 1.090000 ;
      RECT 3.140000 1.280000 3.310000 1.450000 ;
      RECT 3.140000 1.640000 3.310000 1.810000 ;
      RECT 3.140000 2.000000 3.310000 2.170000 ;
      RECT 3.140000 2.360000 3.310000 2.530000 ;
      RECT 3.140000 2.720000 3.310000 2.890000 ;
      RECT 3.140000 3.080000 3.310000 3.250000 ;
      RECT 3.140000 3.440000 3.310000 3.610000 ;
      RECT 3.140000 3.800000 3.310000 3.970000 ;
      RECT 3.140000 4.160000 3.310000 4.330000 ;
      RECT 3.140000 4.520000 3.310000 4.690000 ;
      RECT 3.140000 4.880000 3.310000 5.050000 ;
      RECT 3.140000 5.240000 3.310000 5.410000 ;
    LAYER met1 ;
      RECT 0.700000 0.500000 0.960000 5.470000 ;
      RECT 1.160000 0.500000 1.420000 5.470000 ;
      RECT 1.620000 0.500000 1.880000 5.470000 ;
      RECT 2.080000 0.500000 2.340000 5.470000 ;
      RECT 2.540000 0.500000 2.800000 5.470000 ;
    LAYER via ;
      RECT 0.700000 0.530000 0.960000 0.790000 ;
      RECT 0.700000 0.850000 0.960000 1.110000 ;
      RECT 0.700000 1.170000 0.960000 1.430000 ;
      RECT 0.700000 1.490000 0.960000 1.750000 ;
      RECT 0.700000 1.810000 0.960000 2.070000 ;
      RECT 0.700000 2.130000 0.960000 2.390000 ;
      RECT 0.700000 2.450000 0.960000 2.710000 ;
      RECT 1.160000 3.260000 1.420000 3.520000 ;
      RECT 1.160000 3.580000 1.420000 3.840000 ;
      RECT 1.160000 3.900000 1.420000 4.160000 ;
      RECT 1.160000 4.220000 1.420000 4.480000 ;
      RECT 1.160000 4.540000 1.420000 4.800000 ;
      RECT 1.160000 4.860000 1.420000 5.120000 ;
      RECT 1.160000 5.180000 1.420000 5.440000 ;
      RECT 1.620000 0.530000 1.880000 0.790000 ;
      RECT 1.620000 0.850000 1.880000 1.110000 ;
      RECT 1.620000 1.170000 1.880000 1.430000 ;
      RECT 1.620000 1.490000 1.880000 1.750000 ;
      RECT 1.620000 1.810000 1.880000 2.070000 ;
      RECT 1.620000 2.130000 1.880000 2.390000 ;
      RECT 1.620000 2.450000 1.880000 2.710000 ;
      RECT 2.080000 3.260000 2.340000 3.520000 ;
      RECT 2.080000 3.580000 2.340000 3.840000 ;
      RECT 2.080000 3.900000 2.340000 4.160000 ;
      RECT 2.080000 4.220000 2.340000 4.480000 ;
      RECT 2.080000 4.540000 2.340000 4.800000 ;
      RECT 2.080000 4.860000 2.340000 5.120000 ;
      RECT 2.080000 5.180000 2.340000 5.440000 ;
      RECT 2.540000 0.530000 2.800000 0.790000 ;
      RECT 2.540000 0.850000 2.800000 1.110000 ;
      RECT 2.540000 1.170000 2.800000 1.430000 ;
      RECT 2.540000 1.490000 2.800000 1.750000 ;
      RECT 2.540000 1.810000 2.800000 2.070000 ;
      RECT 2.540000 2.130000 2.800000 2.390000 ;
      RECT 2.540000 2.450000 2.800000 2.710000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18
END LIBRARY
