# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_55p8x11p7_pol1m1m2m3m4m5_noshield_m5pullin
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_55p8x11p7_pol1m1m2m3m4m5_noshield_m5pullin ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  55.73000 BY  11.69000 ;
  OBS
    LAYER li1 ;
      RECT  0.000000  0.000000 55.730000  0.330000 ;
      RECT  0.000000  0.330000  0.140000 11.220000 ;
      RECT  0.000000 11.360000 55.730000 11.690000 ;
      RECT  0.280000  0.470000  0.420000 11.360000 ;
      RECT  0.560000  0.330000  0.700000 11.220000 ;
      RECT  0.840000  0.470000  0.980000 11.360000 ;
      RECT  1.120000  0.330000  1.260000 11.220000 ;
      RECT  1.400000  0.470000  1.540000 11.360000 ;
      RECT  1.680000  0.330000  1.820000 11.220000 ;
      RECT  1.960000  0.470000  2.100000 11.360000 ;
      RECT  2.240000  0.330000  2.380000 11.220000 ;
      RECT  2.520000  0.470000  2.660000 11.360000 ;
      RECT  2.800000  0.330000  2.940000 11.220000 ;
      RECT  3.080000  0.470000  3.220000 11.360000 ;
      RECT  3.360000  0.330000  3.500000 11.220000 ;
      RECT  3.640000  0.470000  3.780000 11.360000 ;
      RECT  3.920000  0.330000  4.060000 11.220000 ;
      RECT  4.200000  0.470000  4.340000 11.360000 ;
      RECT  4.480000  0.330000  4.620000 11.220000 ;
      RECT  4.760000  0.470000  4.900000 11.360000 ;
      RECT  5.040000  0.330000  5.180000 11.220000 ;
      RECT  5.320000  0.470000  5.460000 11.360000 ;
      RECT  5.600000  0.330000  5.740000 11.220000 ;
      RECT  5.880000  0.470000  6.020000 11.360000 ;
      RECT  6.160000  0.330000  6.300000 11.220000 ;
      RECT  6.440000  0.470000  6.580000 11.360000 ;
      RECT  6.720000  0.330000  6.860000 11.220000 ;
      RECT  7.000000  0.470000  7.140000 11.360000 ;
      RECT  7.280000  0.330000  7.420000 11.220000 ;
      RECT  7.560000  0.470000  7.700000 11.360000 ;
      RECT  7.840000  0.330000  7.980000 11.220000 ;
      RECT  8.120000  0.470000  8.260000 11.360000 ;
      RECT  8.400000  0.330000  8.540000 11.220000 ;
      RECT  8.680000  0.470000  8.820000 11.360000 ;
      RECT  8.960000  0.330000  9.100000 11.220000 ;
      RECT  9.240000  0.470000  9.380000 11.360000 ;
      RECT  9.520000  0.330000  9.660000 11.220000 ;
      RECT  9.800000  0.470000  9.940000 11.360000 ;
      RECT 10.080000  0.330000 10.220000 11.220000 ;
      RECT 10.360000  0.470000 10.500000 11.360000 ;
      RECT 10.640000  0.330000 10.780000 11.220000 ;
      RECT 10.920000  0.470000 11.060000 11.360000 ;
      RECT 11.200000  0.330000 11.340000 11.220000 ;
      RECT 11.480000  0.470000 11.620000 11.360000 ;
      RECT 11.760000  0.330000 11.900000 11.220000 ;
      RECT 12.040000  0.470000 12.180000 11.360000 ;
      RECT 12.320000  0.330000 12.460000 11.220000 ;
      RECT 12.600000  0.470000 12.740000 11.360000 ;
      RECT 12.880000  0.330000 13.020000 11.220000 ;
      RECT 13.160000  0.470000 13.300000 11.360000 ;
      RECT 13.440000  0.330000 13.580000 11.220000 ;
      RECT 13.720000  0.470000 13.860000 11.360000 ;
      RECT 14.000000  0.330000 14.140000 11.220000 ;
      RECT 14.280000  0.470000 14.420000 11.360000 ;
      RECT 14.560000  0.330000 14.700000 11.220000 ;
      RECT 14.840000  0.470000 14.980000 11.360000 ;
      RECT 15.120000  0.330000 15.260000 11.220000 ;
      RECT 15.400000  0.470000 15.540000 11.360000 ;
      RECT 15.680000  0.330000 15.820000 11.220000 ;
      RECT 15.960000  0.470000 16.100000 11.360000 ;
      RECT 16.240000  0.330000 16.380000 11.220000 ;
      RECT 16.520000  0.470000 16.660000 11.360000 ;
      RECT 16.800000  0.330000 16.940000 11.220000 ;
      RECT 17.080000  0.470000 17.220000 11.360000 ;
      RECT 17.360000  0.330000 17.500000 11.220000 ;
      RECT 17.640000  0.470000 17.780000 11.360000 ;
      RECT 17.920000  0.330000 18.060000 11.220000 ;
      RECT 18.200000  0.470000 18.340000 11.360000 ;
      RECT 18.480000  0.330000 18.620000 11.220000 ;
      RECT 18.760000  0.470000 18.900000 11.360000 ;
      RECT 19.040000  0.330000 19.180000 11.220000 ;
      RECT 19.320000  0.470000 19.460000 11.360000 ;
      RECT 19.600000  0.330000 19.740000 11.220000 ;
      RECT 19.880000  0.470000 20.020000 11.360000 ;
      RECT 20.160000  0.330000 20.300000 11.220000 ;
      RECT 20.440000  0.470000 20.580000 11.360000 ;
      RECT 20.720000  0.330000 20.860000 11.220000 ;
      RECT 21.000000  0.470000 21.140000 11.360000 ;
      RECT 21.280000  0.330000 21.420000 11.220000 ;
      RECT 21.560000  0.470000 21.700000 11.360000 ;
      RECT 21.840000  0.330000 21.980000 11.220000 ;
      RECT 22.120000  0.470000 22.260000 11.360000 ;
      RECT 22.400000  0.330000 22.540000 11.220000 ;
      RECT 22.680000  0.470000 22.820000 11.360000 ;
      RECT 22.960000  0.330000 23.100000 11.220000 ;
      RECT 23.240000  0.470000 23.380000 11.360000 ;
      RECT 23.520000  0.330000 23.660000 11.220000 ;
      RECT 23.800000  0.470000 23.940000 11.360000 ;
      RECT 24.080000  0.330000 24.220000 11.220000 ;
      RECT 24.360000  0.470000 24.500000 11.360000 ;
      RECT 24.640000  0.330000 24.780000 11.220000 ;
      RECT 24.920000  0.470000 25.060000 11.360000 ;
      RECT 25.200000  0.330000 25.340000 11.220000 ;
      RECT 25.480000  0.470000 25.620000 11.360000 ;
      RECT 25.760000  0.330000 25.900000 11.220000 ;
      RECT 26.040000  0.470000 26.180000 11.360000 ;
      RECT 26.320000  0.330000 26.460000 11.220000 ;
      RECT 26.600000  0.470000 26.740000 11.360000 ;
      RECT 26.880000  0.330000 27.020000 11.220000 ;
      RECT 27.160000  0.470000 27.300000 11.360000 ;
      RECT 27.440000  0.330000 27.580000 11.220000 ;
      RECT 27.720000  0.470000 27.860000 11.360000 ;
      RECT 28.000000  0.330000 28.140000 11.220000 ;
      RECT 28.280000  0.470000 28.420000 11.360000 ;
      RECT 28.560000  0.330000 28.700000 11.220000 ;
      RECT 28.840000  0.470000 28.980000 11.360000 ;
      RECT 29.120000  0.330000 29.260000 11.220000 ;
      RECT 29.400000  0.470000 29.540000 11.360000 ;
      RECT 29.680000  0.330000 29.820000 11.220000 ;
      RECT 29.960000  0.470000 30.100000 11.360000 ;
      RECT 30.240000  0.330000 30.380000 11.220000 ;
      RECT 30.520000  0.470000 30.660000 11.360000 ;
      RECT 30.800000  0.330000 30.940000 11.220000 ;
      RECT 31.080000  0.470000 31.220000 11.360000 ;
      RECT 31.360000  0.330000 31.500000 11.220000 ;
      RECT 31.640000  0.470000 31.780000 11.360000 ;
      RECT 31.920000  0.330000 32.060000 11.220000 ;
      RECT 32.200000  0.470000 32.340000 11.360000 ;
      RECT 32.480000  0.330000 32.620000 11.220000 ;
      RECT 32.760000  0.470000 32.900000 11.360000 ;
      RECT 33.040000  0.330000 33.180000 11.220000 ;
      RECT 33.320000  0.470000 33.460000 11.360000 ;
      RECT 33.600000  0.330000 33.740000 11.220000 ;
      RECT 33.880000  0.470000 34.020000 11.360000 ;
      RECT 34.160000  0.330000 34.300000 11.220000 ;
      RECT 34.440000  0.470000 34.580000 11.360000 ;
      RECT 34.720000  0.330000 34.860000 11.220000 ;
      RECT 35.000000  0.470000 35.140000 11.360000 ;
      RECT 35.280000  0.330000 35.420000 11.220000 ;
      RECT 35.560000  0.470000 35.700000 11.360000 ;
      RECT 35.840000  0.330000 35.980000 11.220000 ;
      RECT 36.120000  0.470000 36.260000 11.360000 ;
      RECT 36.400000  0.330000 36.540000 11.220000 ;
      RECT 36.680000  0.470000 36.820000 11.360000 ;
      RECT 36.960000  0.330000 37.100000 11.220000 ;
      RECT 37.240000  0.470000 37.380000 11.360000 ;
      RECT 37.520000  0.330000 37.660000 11.220000 ;
      RECT 37.800000  0.470000 37.940000 11.360000 ;
      RECT 38.080000  0.330000 38.220000 11.220000 ;
      RECT 38.360000  0.470000 38.500000 11.360000 ;
      RECT 38.640000  0.330000 38.780000 11.220000 ;
      RECT 38.920000  0.470000 39.060000 11.360000 ;
      RECT 39.200000  0.330000 39.340000 11.220000 ;
      RECT 39.480000  0.470000 39.620000 11.360000 ;
      RECT 39.760000  0.330000 39.900000 11.220000 ;
      RECT 40.040000  0.470000 40.180000 11.360000 ;
      RECT 40.320000  0.330000 40.460000 11.220000 ;
      RECT 40.600000  0.470000 40.740000 11.360000 ;
      RECT 40.880000  0.330000 41.020000 11.220000 ;
      RECT 41.160000  0.470000 41.300000 11.360000 ;
      RECT 41.440000  0.330000 41.580000 11.220000 ;
      RECT 41.720000  0.470000 41.860000 11.360000 ;
      RECT 42.000000  0.330000 42.140000 11.220000 ;
      RECT 42.280000  0.470000 42.420000 11.360000 ;
      RECT 42.560000  0.330000 42.700000 11.220000 ;
      RECT 42.840000  0.470000 42.980000 11.360000 ;
      RECT 43.120000  0.330000 43.260000 11.220000 ;
      RECT 43.400000  0.470000 43.540000 11.360000 ;
      RECT 43.680000  0.330000 43.820000 11.220000 ;
      RECT 43.960000  0.470000 44.100000 11.360000 ;
      RECT 44.240000  0.330000 44.380000 11.220000 ;
      RECT 44.520000  0.470000 44.660000 11.360000 ;
      RECT 44.800000  0.330000 44.940000 11.220000 ;
      RECT 45.080000  0.470000 45.220000 11.360000 ;
      RECT 45.360000  0.330000 45.500000 11.220000 ;
      RECT 45.640000  0.470000 45.780000 11.360000 ;
      RECT 45.920000  0.330000 46.060000 11.220000 ;
      RECT 46.200000  0.470000 46.340000 11.360000 ;
      RECT 46.480000  0.330000 46.620000 11.220000 ;
      RECT 46.760000  0.470000 46.900000 11.360000 ;
      RECT 47.040000  0.330000 47.180000 11.220000 ;
      RECT 47.320000  0.470000 47.460000 11.360000 ;
      RECT 47.600000  0.330000 47.740000 11.220000 ;
      RECT 47.880000  0.470000 48.020000 11.360000 ;
      RECT 48.160000  0.330000 48.300000 11.220000 ;
      RECT 48.440000  0.470000 48.580000 11.360000 ;
      RECT 48.720000  0.330000 48.860000 11.220000 ;
      RECT 49.000000  0.470000 49.140000 11.360000 ;
      RECT 49.280000  0.330000 49.420000 11.220000 ;
      RECT 49.560000  0.470000 49.700000 11.360000 ;
      RECT 49.840000  0.330000 49.980000 11.220000 ;
      RECT 50.120000  0.470000 50.260000 11.360000 ;
      RECT 50.400000  0.330000 50.540000 11.220000 ;
      RECT 50.680000  0.470000 50.820000 11.360000 ;
      RECT 50.960000  0.330000 51.100000 11.220000 ;
      RECT 51.240000  0.470000 51.380000 11.360000 ;
      RECT 51.520000  0.330000 51.660000 11.220000 ;
      RECT 51.800000  0.470000 51.940000 11.360000 ;
      RECT 52.080000  0.330000 52.220000 11.220000 ;
      RECT 52.360000  0.470000 52.500000 11.360000 ;
      RECT 52.640000  0.330000 52.780000 11.220000 ;
      RECT 52.920000  0.470000 53.060000 11.360000 ;
      RECT 53.200000  0.330000 53.340000 11.220000 ;
      RECT 53.480000  0.470000 53.620000 11.360000 ;
      RECT 53.760000  0.330000 53.900000 11.220000 ;
      RECT 54.040000  0.470000 54.180000 11.360000 ;
      RECT 54.320000  0.330000 54.460000 11.220000 ;
      RECT 54.600000  0.470000 54.740000 11.360000 ;
      RECT 54.880000  0.330000 55.020000 11.220000 ;
      RECT 55.160000  0.470000 55.300000 11.360000 ;
      RECT 55.440000  0.330000 55.730000 11.220000 ;
    LAYER mcon ;
      RECT  0.190000  0.080000  0.360000  0.250000 ;
      RECT  0.190000 11.440000  0.360000 11.610000 ;
      RECT  0.550000  0.080000  0.720000  0.250000 ;
      RECT  0.550000 11.440000  0.720000 11.610000 ;
      RECT  0.910000  0.080000  1.080000  0.250000 ;
      RECT  0.910000 11.440000  1.080000 11.610000 ;
      RECT  1.270000  0.080000  1.440000  0.250000 ;
      RECT  1.270000 11.440000  1.440000 11.610000 ;
      RECT  1.630000  0.080000  1.800000  0.250000 ;
      RECT  1.630000 11.440000  1.800000 11.610000 ;
      RECT  1.990000  0.080000  2.160000  0.250000 ;
      RECT  1.990000 11.440000  2.160000 11.610000 ;
      RECT  2.350000  0.080000  2.520000  0.250000 ;
      RECT  2.350000 11.440000  2.520000 11.610000 ;
      RECT  2.710000  0.080000  2.880000  0.250000 ;
      RECT  2.710000 11.440000  2.880000 11.610000 ;
      RECT  3.070000  0.080000  3.240000  0.250000 ;
      RECT  3.070000 11.440000  3.240000 11.610000 ;
      RECT  3.430000  0.080000  3.600000  0.250000 ;
      RECT  3.430000 11.440000  3.600000 11.610000 ;
      RECT  3.790000  0.080000  3.960000  0.250000 ;
      RECT  3.790000 11.440000  3.960000 11.610000 ;
      RECT  4.150000  0.080000  4.320000  0.250000 ;
      RECT  4.150000 11.440000  4.320000 11.610000 ;
      RECT  4.510000  0.080000  4.680000  0.250000 ;
      RECT  4.510000 11.440000  4.680000 11.610000 ;
      RECT  4.870000  0.080000  5.040000  0.250000 ;
      RECT  4.870000 11.440000  5.040000 11.610000 ;
      RECT  5.230000  0.080000  5.400000  0.250000 ;
      RECT  5.230000 11.440000  5.400000 11.610000 ;
      RECT  5.590000  0.080000  5.760000  0.250000 ;
      RECT  5.590000 11.440000  5.760000 11.610000 ;
      RECT  5.950000  0.080000  6.120000  0.250000 ;
      RECT  5.950000 11.440000  6.120000 11.610000 ;
      RECT  6.310000  0.080000  6.480000  0.250000 ;
      RECT  6.310000 11.440000  6.480000 11.610000 ;
      RECT  6.670000  0.080000  6.840000  0.250000 ;
      RECT  6.670000 11.440000  6.840000 11.610000 ;
      RECT  7.030000  0.080000  7.200000  0.250000 ;
      RECT  7.030000 11.440000  7.200000 11.610000 ;
      RECT  7.390000  0.080000  7.560000  0.250000 ;
      RECT  7.390000 11.440000  7.560000 11.610000 ;
      RECT  7.750000  0.080000  7.920000  0.250000 ;
      RECT  7.750000 11.440000  7.920000 11.610000 ;
      RECT  8.110000  0.080000  8.280000  0.250000 ;
      RECT  8.110000 11.440000  8.280000 11.610000 ;
      RECT  8.470000  0.080000  8.640000  0.250000 ;
      RECT  8.470000 11.440000  8.640000 11.610000 ;
      RECT  8.830000  0.080000  9.000000  0.250000 ;
      RECT  8.830000 11.440000  9.000000 11.610000 ;
      RECT  9.190000  0.080000  9.360000  0.250000 ;
      RECT  9.190000 11.440000  9.360000 11.610000 ;
      RECT  9.550000  0.080000  9.720000  0.250000 ;
      RECT  9.550000 11.440000  9.720000 11.610000 ;
      RECT  9.910000  0.080000 10.080000  0.250000 ;
      RECT  9.910000 11.440000 10.080000 11.610000 ;
      RECT 10.270000  0.080000 10.440000  0.250000 ;
      RECT 10.270000 11.440000 10.440000 11.610000 ;
      RECT 10.630000  0.080000 10.800000  0.250000 ;
      RECT 10.630000 11.440000 10.800000 11.610000 ;
      RECT 10.990000  0.080000 11.160000  0.250000 ;
      RECT 10.990000 11.440000 11.160000 11.610000 ;
      RECT 11.350000  0.080000 11.520000  0.250000 ;
      RECT 11.350000 11.440000 11.520000 11.610000 ;
      RECT 11.710000  0.080000 11.880000  0.250000 ;
      RECT 11.710000 11.440000 11.880000 11.610000 ;
      RECT 12.070000  0.080000 12.240000  0.250000 ;
      RECT 12.070000 11.440000 12.240000 11.610000 ;
      RECT 12.430000  0.080000 12.600000  0.250000 ;
      RECT 12.430000 11.440000 12.600000 11.610000 ;
      RECT 12.790000  0.080000 12.960000  0.250000 ;
      RECT 12.790000 11.440000 12.960000 11.610000 ;
      RECT 13.150000  0.080000 13.320000  0.250000 ;
      RECT 13.150000 11.440000 13.320000 11.610000 ;
      RECT 13.510000  0.080000 13.680000  0.250000 ;
      RECT 13.510000 11.440000 13.680000 11.610000 ;
      RECT 13.870000  0.080000 14.040000  0.250000 ;
      RECT 13.870000 11.440000 14.040000 11.610000 ;
      RECT 14.230000  0.080000 14.400000  0.250000 ;
      RECT 14.230000 11.440000 14.400000 11.610000 ;
      RECT 14.590000  0.080000 14.760000  0.250000 ;
      RECT 14.590000 11.440000 14.760000 11.610000 ;
      RECT 14.950000  0.080000 15.120000  0.250000 ;
      RECT 14.950000 11.440000 15.120000 11.610000 ;
      RECT 15.310000  0.080000 15.480000  0.250000 ;
      RECT 15.310000 11.440000 15.480000 11.610000 ;
      RECT 15.670000  0.080000 15.840000  0.250000 ;
      RECT 15.670000 11.440000 15.840000 11.610000 ;
      RECT 16.030000  0.080000 16.200000  0.250000 ;
      RECT 16.030000 11.440000 16.200000 11.610000 ;
      RECT 16.390000  0.080000 16.560000  0.250000 ;
      RECT 16.390000 11.440000 16.560000 11.610000 ;
      RECT 16.750000  0.080000 16.920000  0.250000 ;
      RECT 16.750000 11.440000 16.920000 11.610000 ;
      RECT 17.110000  0.080000 17.280000  0.250000 ;
      RECT 17.110000 11.440000 17.280000 11.610000 ;
      RECT 17.470000  0.080000 17.640000  0.250000 ;
      RECT 17.470000 11.440000 17.640000 11.610000 ;
      RECT 17.830000  0.080000 18.000000  0.250000 ;
      RECT 17.830000 11.440000 18.000000 11.610000 ;
      RECT 18.190000  0.080000 18.360000  0.250000 ;
      RECT 18.190000 11.440000 18.360000 11.610000 ;
      RECT 18.550000  0.080000 18.720000  0.250000 ;
      RECT 18.550000 11.440000 18.720000 11.610000 ;
      RECT 18.910000  0.080000 19.080000  0.250000 ;
      RECT 18.910000 11.440000 19.080000 11.610000 ;
      RECT 19.270000  0.080000 19.440000  0.250000 ;
      RECT 19.270000 11.440000 19.440000 11.610000 ;
      RECT 19.630000  0.080000 19.800000  0.250000 ;
      RECT 19.630000 11.440000 19.800000 11.610000 ;
      RECT 19.990000  0.080000 20.160000  0.250000 ;
      RECT 19.990000 11.440000 20.160000 11.610000 ;
      RECT 20.350000  0.080000 20.520000  0.250000 ;
      RECT 20.350000 11.440000 20.520000 11.610000 ;
      RECT 20.710000  0.080000 20.880000  0.250000 ;
      RECT 20.710000 11.440000 20.880000 11.610000 ;
      RECT 21.070000  0.080000 21.240000  0.250000 ;
      RECT 21.070000 11.440000 21.240000 11.610000 ;
      RECT 21.430000  0.080000 21.600000  0.250000 ;
      RECT 21.430000 11.440000 21.600000 11.610000 ;
      RECT 21.790000  0.080000 21.960000  0.250000 ;
      RECT 21.790000 11.440000 21.960000 11.610000 ;
      RECT 22.150000  0.080000 22.320000  0.250000 ;
      RECT 22.150000 11.440000 22.320000 11.610000 ;
      RECT 22.510000  0.080000 22.680000  0.250000 ;
      RECT 22.510000 11.440000 22.680000 11.610000 ;
      RECT 22.870000  0.080000 23.040000  0.250000 ;
      RECT 22.870000 11.440000 23.040000 11.610000 ;
      RECT 23.230000  0.080000 23.400000  0.250000 ;
      RECT 23.230000 11.440000 23.400000 11.610000 ;
      RECT 23.590000  0.080000 23.760000  0.250000 ;
      RECT 23.590000 11.440000 23.760000 11.610000 ;
      RECT 23.950000  0.080000 24.120000  0.250000 ;
      RECT 23.950000 11.440000 24.120000 11.610000 ;
      RECT 24.310000  0.080000 24.480000  0.250000 ;
      RECT 24.310000 11.440000 24.480000 11.610000 ;
      RECT 24.670000  0.080000 24.840000  0.250000 ;
      RECT 24.670000 11.440000 24.840000 11.610000 ;
      RECT 25.030000  0.080000 25.200000  0.250000 ;
      RECT 25.030000 11.440000 25.200000 11.610000 ;
      RECT 25.390000  0.080000 25.560000  0.250000 ;
      RECT 25.390000 11.440000 25.560000 11.610000 ;
      RECT 25.750000  0.080000 25.920000  0.250000 ;
      RECT 25.750000 11.440000 25.920000 11.610000 ;
      RECT 26.110000  0.080000 26.280000  0.250000 ;
      RECT 26.110000 11.440000 26.280000 11.610000 ;
      RECT 26.470000  0.080000 26.640000  0.250000 ;
      RECT 26.470000 11.440000 26.640000 11.610000 ;
      RECT 26.830000  0.080000 27.000000  0.250000 ;
      RECT 26.830000 11.440000 27.000000 11.610000 ;
      RECT 27.190000  0.080000 27.360000  0.250000 ;
      RECT 27.190000 11.440000 27.360000 11.610000 ;
      RECT 27.550000  0.080000 27.720000  0.250000 ;
      RECT 27.550000 11.440000 27.720000 11.610000 ;
      RECT 27.910000  0.080000 28.080000  0.250000 ;
      RECT 27.910000 11.440000 28.080000 11.610000 ;
      RECT 28.270000  0.080000 28.440000  0.250000 ;
      RECT 28.270000 11.440000 28.440000 11.610000 ;
      RECT 28.630000  0.080000 28.800000  0.250000 ;
      RECT 28.630000 11.440000 28.800000 11.610000 ;
      RECT 28.990000  0.080000 29.160000  0.250000 ;
      RECT 28.990000 11.440000 29.160000 11.610000 ;
      RECT 29.350000  0.080000 29.520000  0.250000 ;
      RECT 29.350000 11.440000 29.520000 11.610000 ;
      RECT 29.710000  0.080000 29.880000  0.250000 ;
      RECT 29.710000 11.440000 29.880000 11.610000 ;
      RECT 30.070000  0.080000 30.240000  0.250000 ;
      RECT 30.070000 11.440000 30.240000 11.610000 ;
      RECT 30.430000  0.080000 30.600000  0.250000 ;
      RECT 30.430000 11.440000 30.600000 11.610000 ;
      RECT 30.790000  0.080000 30.960000  0.250000 ;
      RECT 30.790000 11.440000 30.960000 11.610000 ;
      RECT 31.150000  0.080000 31.320000  0.250000 ;
      RECT 31.150000 11.440000 31.320000 11.610000 ;
      RECT 31.510000  0.080000 31.680000  0.250000 ;
      RECT 31.510000 11.440000 31.680000 11.610000 ;
      RECT 31.870000  0.080000 32.040000  0.250000 ;
      RECT 31.870000 11.440000 32.040000 11.610000 ;
      RECT 32.230000  0.080000 32.400000  0.250000 ;
      RECT 32.230000 11.440000 32.400000 11.610000 ;
      RECT 32.590000  0.080000 32.760000  0.250000 ;
      RECT 32.590000 11.440000 32.760000 11.610000 ;
      RECT 32.950000  0.080000 33.120000  0.250000 ;
      RECT 32.950000 11.440000 33.120000 11.610000 ;
      RECT 33.310000  0.080000 33.480000  0.250000 ;
      RECT 33.310000 11.440000 33.480000 11.610000 ;
      RECT 33.670000  0.080000 33.840000  0.250000 ;
      RECT 33.670000 11.440000 33.840000 11.610000 ;
      RECT 34.030000  0.080000 34.200000  0.250000 ;
      RECT 34.030000 11.440000 34.200000 11.610000 ;
      RECT 34.390000  0.080000 34.560000  0.250000 ;
      RECT 34.390000 11.440000 34.560000 11.610000 ;
      RECT 34.750000  0.080000 34.920000  0.250000 ;
      RECT 34.750000 11.440000 34.920000 11.610000 ;
      RECT 35.110000  0.080000 35.280000  0.250000 ;
      RECT 35.110000 11.440000 35.280000 11.610000 ;
      RECT 35.470000  0.080000 35.640000  0.250000 ;
      RECT 35.470000 11.440000 35.640000 11.610000 ;
      RECT 35.830000  0.080000 36.000000  0.250000 ;
      RECT 35.830000 11.440000 36.000000 11.610000 ;
      RECT 36.190000  0.080000 36.360000  0.250000 ;
      RECT 36.190000 11.440000 36.360000 11.610000 ;
      RECT 36.550000  0.080000 36.720000  0.250000 ;
      RECT 36.550000 11.440000 36.720000 11.610000 ;
      RECT 36.910000  0.080000 37.080000  0.250000 ;
      RECT 36.910000 11.440000 37.080000 11.610000 ;
      RECT 37.270000  0.080000 37.440000  0.250000 ;
      RECT 37.270000 11.440000 37.440000 11.610000 ;
      RECT 37.630000  0.080000 37.800000  0.250000 ;
      RECT 37.630000 11.440000 37.800000 11.610000 ;
      RECT 37.990000  0.080000 38.160000  0.250000 ;
      RECT 37.990000 11.440000 38.160000 11.610000 ;
      RECT 38.350000  0.080000 38.520000  0.250000 ;
      RECT 38.350000 11.440000 38.520000 11.610000 ;
      RECT 38.710000  0.080000 38.880000  0.250000 ;
      RECT 38.710000 11.440000 38.880000 11.610000 ;
      RECT 39.070000  0.080000 39.240000  0.250000 ;
      RECT 39.070000 11.440000 39.240000 11.610000 ;
      RECT 39.430000  0.080000 39.600000  0.250000 ;
      RECT 39.430000 11.440000 39.600000 11.610000 ;
      RECT 39.790000  0.080000 39.960000  0.250000 ;
      RECT 39.790000 11.440000 39.960000 11.610000 ;
      RECT 40.150000  0.080000 40.320000  0.250000 ;
      RECT 40.150000 11.440000 40.320000 11.610000 ;
      RECT 40.510000  0.080000 40.680000  0.250000 ;
      RECT 40.510000 11.440000 40.680000 11.610000 ;
      RECT 40.870000  0.080000 41.040000  0.250000 ;
      RECT 40.870000 11.440000 41.040000 11.610000 ;
      RECT 41.230000  0.080000 41.400000  0.250000 ;
      RECT 41.230000 11.440000 41.400000 11.610000 ;
      RECT 41.590000  0.080000 41.760000  0.250000 ;
      RECT 41.590000 11.440000 41.760000 11.610000 ;
      RECT 41.950000  0.080000 42.120000  0.250000 ;
      RECT 41.950000 11.440000 42.120000 11.610000 ;
      RECT 42.310000  0.080000 42.480000  0.250000 ;
      RECT 42.310000 11.440000 42.480000 11.610000 ;
      RECT 42.670000  0.080000 42.840000  0.250000 ;
      RECT 42.670000 11.440000 42.840000 11.610000 ;
      RECT 43.030000  0.080000 43.200000  0.250000 ;
      RECT 43.030000 11.440000 43.200000 11.610000 ;
      RECT 43.390000  0.080000 43.560000  0.250000 ;
      RECT 43.390000 11.440000 43.560000 11.610000 ;
      RECT 43.750000  0.080000 43.920000  0.250000 ;
      RECT 43.750000 11.440000 43.920000 11.610000 ;
      RECT 44.110000  0.080000 44.280000  0.250000 ;
      RECT 44.110000 11.440000 44.280000 11.610000 ;
      RECT 44.470000  0.080000 44.640000  0.250000 ;
      RECT 44.470000 11.440000 44.640000 11.610000 ;
      RECT 44.830000  0.080000 45.000000  0.250000 ;
      RECT 44.830000 11.440000 45.000000 11.610000 ;
      RECT 45.190000  0.080000 45.360000  0.250000 ;
      RECT 45.190000 11.440000 45.360000 11.610000 ;
      RECT 45.550000  0.080000 45.720000  0.250000 ;
      RECT 45.550000 11.440000 45.720000 11.610000 ;
      RECT 45.910000  0.080000 46.080000  0.250000 ;
      RECT 45.910000 11.440000 46.080000 11.610000 ;
      RECT 46.270000  0.080000 46.440000  0.250000 ;
      RECT 46.270000 11.440000 46.440000 11.610000 ;
      RECT 46.630000  0.080000 46.800000  0.250000 ;
      RECT 46.630000 11.440000 46.800000 11.610000 ;
      RECT 46.990000  0.080000 47.160000  0.250000 ;
      RECT 46.990000 11.440000 47.160000 11.610000 ;
      RECT 47.350000  0.080000 47.520000  0.250000 ;
      RECT 47.350000 11.440000 47.520000 11.610000 ;
      RECT 47.710000  0.080000 47.880000  0.250000 ;
      RECT 47.710000 11.440000 47.880000 11.610000 ;
      RECT 48.070000  0.080000 48.240000  0.250000 ;
      RECT 48.070000 11.440000 48.240000 11.610000 ;
      RECT 48.430000  0.080000 48.600000  0.250000 ;
      RECT 48.430000 11.440000 48.600000 11.610000 ;
      RECT 48.790000  0.080000 48.960000  0.250000 ;
      RECT 48.790000 11.440000 48.960000 11.610000 ;
      RECT 49.150000  0.080000 49.320000  0.250000 ;
      RECT 49.150000 11.440000 49.320000 11.610000 ;
      RECT 49.510000  0.080000 49.680000  0.250000 ;
      RECT 49.510000 11.440000 49.680000 11.610000 ;
      RECT 49.870000  0.080000 50.040000  0.250000 ;
      RECT 49.870000 11.440000 50.040000 11.610000 ;
      RECT 50.230000  0.080000 50.400000  0.250000 ;
      RECT 50.230000 11.440000 50.400000 11.610000 ;
      RECT 50.590000  0.080000 50.760000  0.250000 ;
      RECT 50.590000 11.440000 50.760000 11.610000 ;
      RECT 50.950000  0.080000 51.120000  0.250000 ;
      RECT 50.950000 11.440000 51.120000 11.610000 ;
      RECT 51.310000  0.080000 51.480000  0.250000 ;
      RECT 51.310000 11.440000 51.480000 11.610000 ;
      RECT 51.670000  0.080000 51.840000  0.250000 ;
      RECT 51.670000 11.440000 51.840000 11.610000 ;
      RECT 52.030000  0.080000 52.200000  0.250000 ;
      RECT 52.030000 11.440000 52.200000 11.610000 ;
      RECT 52.390000  0.080000 52.560000  0.250000 ;
      RECT 52.390000 11.440000 52.560000 11.610000 ;
      RECT 52.750000  0.080000 52.920000  0.250000 ;
      RECT 52.750000 11.440000 52.920000 11.610000 ;
      RECT 53.110000  0.080000 53.280000  0.250000 ;
      RECT 53.110000 11.440000 53.280000 11.610000 ;
      RECT 53.470000  0.080000 53.640000  0.250000 ;
      RECT 53.470000 11.440000 53.640000 11.610000 ;
      RECT 53.830000  0.080000 54.000000  0.250000 ;
      RECT 53.830000 11.440000 54.000000 11.610000 ;
      RECT 54.190000  0.080000 54.360000  0.250000 ;
      RECT 54.190000 11.440000 54.360000 11.610000 ;
      RECT 54.550000  0.080000 54.720000  0.250000 ;
      RECT 54.550000 11.440000 54.720000 11.610000 ;
      RECT 54.910000  0.080000 55.080000  0.250000 ;
      RECT 54.910000 11.440000 55.080000 11.610000 ;
      RECT 55.270000  0.080000 55.440000  0.250000 ;
      RECT 55.270000 11.440000 55.440000 11.610000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 55.730000  0.330000 ;
      RECT  0.000000  0.470000  0.140000 11.360000 ;
      RECT  0.000000 11.360000 55.730000 11.690000 ;
      RECT  0.280000  0.330000  0.420000 11.220000 ;
      RECT  0.560000  0.470000  0.700000 11.360000 ;
      RECT  0.840000  0.330000  0.980000 11.220000 ;
      RECT  1.120000  0.470000  1.260000 11.360000 ;
      RECT  1.400000  0.330000  1.540000 11.220000 ;
      RECT  1.680000  0.470000  1.820000 11.360000 ;
      RECT  1.960000  0.330000  2.100000 11.220000 ;
      RECT  2.240000  0.470000  2.380000 11.360000 ;
      RECT  2.520000  0.330000  2.660000 11.220000 ;
      RECT  2.800000  0.470000  2.940000 11.360000 ;
      RECT  3.080000  0.330000  3.220000 11.220000 ;
      RECT  3.360000  0.470000  3.500000 11.360000 ;
      RECT  3.640000  0.330000  3.780000 11.220000 ;
      RECT  3.920000  0.470000  4.060000 11.360000 ;
      RECT  4.200000  0.330000  4.340000 11.220000 ;
      RECT  4.480000  0.470000  4.620000 11.360000 ;
      RECT  4.760000  0.330000  4.900000 11.220000 ;
      RECT  5.040000  0.470000  5.180000 11.360000 ;
      RECT  5.320000  0.330000  5.460000 11.220000 ;
      RECT  5.600000  0.470000  5.740000 11.360000 ;
      RECT  5.880000  0.330000  6.020000 11.220000 ;
      RECT  6.160000  0.470000  6.300000 11.360000 ;
      RECT  6.440000  0.330000  6.580000 11.220000 ;
      RECT  6.720000  0.470000  6.860000 11.360000 ;
      RECT  7.000000  0.330000  7.140000 11.220000 ;
      RECT  7.280000  0.470000  7.420000 11.360000 ;
      RECT  7.560000  0.330000  7.700000 11.220000 ;
      RECT  7.840000  0.470000  7.980000 11.360000 ;
      RECT  8.120000  0.330000  8.260000 11.220000 ;
      RECT  8.400000  0.470000  8.540000 11.360000 ;
      RECT  8.680000  0.330000  8.820000 11.220000 ;
      RECT  8.960000  0.470000  9.100000 11.360000 ;
      RECT  9.240000  0.330000  9.380000 11.220000 ;
      RECT  9.520000  0.470000  9.660000 11.360000 ;
      RECT  9.800000  0.330000  9.940000 11.220000 ;
      RECT 10.080000  0.470000 10.220000 11.360000 ;
      RECT 10.360000  0.330000 10.500000 11.220000 ;
      RECT 10.640000  0.470000 10.780000 11.360000 ;
      RECT 10.920000  0.330000 11.060000 11.220000 ;
      RECT 11.200000  0.470000 11.340000 11.360000 ;
      RECT 11.480000  0.330000 11.620000 11.220000 ;
      RECT 11.760000  0.470000 11.900000 11.360000 ;
      RECT 12.040000  0.330000 12.180000 11.220000 ;
      RECT 12.320000  0.470000 12.460000 11.360000 ;
      RECT 12.600000  0.330000 12.740000 11.220000 ;
      RECT 12.880000  0.470000 13.020000 11.360000 ;
      RECT 13.160000  0.330000 13.300000 11.220000 ;
      RECT 13.440000  0.470000 13.580000 11.360000 ;
      RECT 13.720000  0.330000 13.860000 11.220000 ;
      RECT 14.000000  0.470000 14.140000 11.360000 ;
      RECT 14.280000  0.330000 14.420000 11.220000 ;
      RECT 14.560000  0.470000 14.700000 11.360000 ;
      RECT 14.840000  0.330000 14.980000 11.220000 ;
      RECT 15.120000  0.470000 15.260000 11.360000 ;
      RECT 15.400000  0.330000 15.540000 11.220000 ;
      RECT 15.680000  0.470000 15.820000 11.360000 ;
      RECT 15.960000  0.330000 16.100000 11.220000 ;
      RECT 16.240000  0.470000 16.380000 11.360000 ;
      RECT 16.520000  0.330000 16.660000 11.220000 ;
      RECT 16.800000  0.470000 16.940000 11.360000 ;
      RECT 17.080000  0.330000 17.220000 11.220000 ;
      RECT 17.360000  0.470000 17.500000 11.360000 ;
      RECT 17.640000  0.330000 17.780000 11.220000 ;
      RECT 17.920000  0.470000 18.060000 11.360000 ;
      RECT 18.200000  0.330000 18.340000 11.220000 ;
      RECT 18.480000  0.470000 18.620000 11.360000 ;
      RECT 18.760000  0.330000 18.900000 11.220000 ;
      RECT 19.040000  0.470000 19.180000 11.360000 ;
      RECT 19.320000  0.330000 19.460000 11.220000 ;
      RECT 19.600000  0.470000 19.740000 11.360000 ;
      RECT 19.880000  0.330000 20.020000 11.220000 ;
      RECT 20.160000  0.470000 20.300000 11.360000 ;
      RECT 20.440000  0.330000 20.580000 11.220000 ;
      RECT 20.720000  0.470000 20.860000 11.360000 ;
      RECT 21.000000  0.330000 21.140000 11.220000 ;
      RECT 21.280000  0.470000 21.420000 11.360000 ;
      RECT 21.560000  0.330000 21.700000 11.220000 ;
      RECT 21.840000  0.470000 21.980000 11.360000 ;
      RECT 22.120000  0.330000 22.260000 11.220000 ;
      RECT 22.400000  0.470000 22.540000 11.360000 ;
      RECT 22.680000  0.330000 22.820000 11.220000 ;
      RECT 22.960000  0.470000 23.100000 11.360000 ;
      RECT 23.240000  0.330000 23.380000 11.220000 ;
      RECT 23.520000  0.470000 23.660000 11.360000 ;
      RECT 23.800000  0.330000 23.940000 11.220000 ;
      RECT 24.080000  0.470000 24.220000 11.360000 ;
      RECT 24.360000  0.330000 24.500000 11.220000 ;
      RECT 24.640000  0.470000 24.780000 11.360000 ;
      RECT 24.920000  0.330000 25.060000 11.220000 ;
      RECT 25.200000  0.470000 25.340000 11.360000 ;
      RECT 25.480000  0.330000 25.620000 11.220000 ;
      RECT 25.760000  0.470000 25.900000 11.360000 ;
      RECT 26.040000  0.330000 26.180000 11.220000 ;
      RECT 26.320000  0.470000 26.460000 11.360000 ;
      RECT 26.600000  0.330000 26.740000 11.220000 ;
      RECT 26.880000  0.470000 27.020000 11.360000 ;
      RECT 27.160000  0.330000 27.300000 11.220000 ;
      RECT 27.440000  0.470000 27.580000 11.360000 ;
      RECT 27.720000  0.330000 27.860000 11.220000 ;
      RECT 28.000000  0.470000 28.140000 11.360000 ;
      RECT 28.280000  0.330000 28.420000 11.220000 ;
      RECT 28.560000  0.470000 28.700000 11.360000 ;
      RECT 28.840000  0.330000 28.980000 11.220000 ;
      RECT 29.120000  0.470000 29.260000 11.360000 ;
      RECT 29.400000  0.330000 29.540000 11.220000 ;
      RECT 29.680000  0.470000 29.820000 11.360000 ;
      RECT 29.960000  0.330000 30.100000 11.220000 ;
      RECT 30.240000  0.470000 30.380000 11.360000 ;
      RECT 30.520000  0.330000 30.660000 11.220000 ;
      RECT 30.800000  0.470000 30.940000 11.360000 ;
      RECT 31.080000  0.330000 31.220000 11.220000 ;
      RECT 31.360000  0.470000 31.500000 11.360000 ;
      RECT 31.640000  0.330000 31.780000 11.220000 ;
      RECT 31.920000  0.470000 32.060000 11.360000 ;
      RECT 32.200000  0.330000 32.340000 11.220000 ;
      RECT 32.480000  0.470000 32.620000 11.360000 ;
      RECT 32.760000  0.330000 32.900000 11.220000 ;
      RECT 33.040000  0.470000 33.180000 11.360000 ;
      RECT 33.320000  0.330000 33.460000 11.220000 ;
      RECT 33.600000  0.470000 33.740000 11.360000 ;
      RECT 33.880000  0.330000 34.020000 11.220000 ;
      RECT 34.160000  0.470000 34.300000 11.360000 ;
      RECT 34.440000  0.330000 34.580000 11.220000 ;
      RECT 34.720000  0.470000 34.860000 11.360000 ;
      RECT 35.000000  0.330000 35.140000 11.220000 ;
      RECT 35.280000  0.470000 35.420000 11.360000 ;
      RECT 35.560000  0.330000 35.700000 11.220000 ;
      RECT 35.840000  0.470000 35.980000 11.360000 ;
      RECT 36.120000  0.330000 36.260000 11.220000 ;
      RECT 36.400000  0.470000 36.540000 11.360000 ;
      RECT 36.680000  0.330000 36.820000 11.220000 ;
      RECT 36.960000  0.470000 37.100000 11.360000 ;
      RECT 37.240000  0.330000 37.380000 11.220000 ;
      RECT 37.520000  0.470000 37.660000 11.360000 ;
      RECT 37.800000  0.330000 37.940000 11.220000 ;
      RECT 38.080000  0.470000 38.220000 11.360000 ;
      RECT 38.360000  0.330000 38.500000 11.220000 ;
      RECT 38.640000  0.470000 38.780000 11.360000 ;
      RECT 38.920000  0.330000 39.060000 11.220000 ;
      RECT 39.200000  0.470000 39.340000 11.360000 ;
      RECT 39.480000  0.330000 39.620000 11.220000 ;
      RECT 39.760000  0.470000 39.900000 11.360000 ;
      RECT 40.040000  0.330000 40.180000 11.220000 ;
      RECT 40.320000  0.470000 40.460000 11.360000 ;
      RECT 40.600000  0.330000 40.740000 11.220000 ;
      RECT 40.880000  0.470000 41.020000 11.360000 ;
      RECT 41.160000  0.330000 41.300000 11.220000 ;
      RECT 41.440000  0.470000 41.580000 11.360000 ;
      RECT 41.720000  0.330000 41.860000 11.220000 ;
      RECT 42.000000  0.470000 42.140000 11.360000 ;
      RECT 42.280000  0.330000 42.420000 11.220000 ;
      RECT 42.560000  0.470000 42.700000 11.360000 ;
      RECT 42.840000  0.330000 42.980000 11.220000 ;
      RECT 43.120000  0.470000 43.260000 11.360000 ;
      RECT 43.400000  0.330000 43.540000 11.220000 ;
      RECT 43.680000  0.470000 43.820000 11.360000 ;
      RECT 43.960000  0.330000 44.100000 11.220000 ;
      RECT 44.240000  0.470000 44.380000 11.360000 ;
      RECT 44.520000  0.330000 44.660000 11.220000 ;
      RECT 44.800000  0.470000 44.940000 11.360000 ;
      RECT 45.080000  0.330000 45.220000 11.220000 ;
      RECT 45.360000  0.470000 45.500000 11.360000 ;
      RECT 45.640000  0.330000 45.780000 11.220000 ;
      RECT 45.920000  0.470000 46.060000 11.360000 ;
      RECT 46.200000  0.330000 46.340000 11.220000 ;
      RECT 46.480000  0.470000 46.620000 11.360000 ;
      RECT 46.760000  0.330000 46.900000 11.220000 ;
      RECT 47.040000  0.470000 47.180000 11.360000 ;
      RECT 47.320000  0.330000 47.460000 11.220000 ;
      RECT 47.600000  0.470000 47.740000 11.360000 ;
      RECT 47.880000  0.330000 48.020000 11.220000 ;
      RECT 48.160000  0.470000 48.300000 11.360000 ;
      RECT 48.440000  0.330000 48.580000 11.220000 ;
      RECT 48.720000  0.470000 48.860000 11.360000 ;
      RECT 49.000000  0.330000 49.140000 11.220000 ;
      RECT 49.280000  0.470000 49.420000 11.360000 ;
      RECT 49.560000  0.330000 49.700000 11.220000 ;
      RECT 49.840000  0.470000 49.980000 11.360000 ;
      RECT 50.120000  0.330000 50.260000 11.220000 ;
      RECT 50.400000  0.470000 50.540000 11.360000 ;
      RECT 50.680000  0.330000 50.820000 11.220000 ;
      RECT 50.960000  0.470000 51.100000 11.360000 ;
      RECT 51.240000  0.330000 51.380000 11.220000 ;
      RECT 51.520000  0.470000 51.660000 11.360000 ;
      RECT 51.800000  0.330000 51.940000 11.220000 ;
      RECT 52.080000  0.470000 52.220000 11.360000 ;
      RECT 52.360000  0.330000 52.500000 11.220000 ;
      RECT 52.640000  0.470000 52.780000 11.360000 ;
      RECT 52.920000  0.330000 53.060000 11.220000 ;
      RECT 53.200000  0.470000 53.340000 11.360000 ;
      RECT 53.480000  0.330000 53.620000 11.220000 ;
      RECT 53.760000  0.470000 53.900000 11.360000 ;
      RECT 54.040000  0.330000 54.180000 11.220000 ;
      RECT 54.320000  0.470000 54.460000 11.360000 ;
      RECT 54.600000  0.330000 54.740000 11.220000 ;
      RECT 54.880000  0.470000 55.020000 11.360000 ;
      RECT 55.160000  0.330000 55.300000 11.220000 ;
      RECT 55.440000  0.470000 55.730000 11.360000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  0.700000  0.330000 ;
      RECT  0.000000  0.330000  0.140000 11.690000 ;
      RECT  0.280000  0.470000  0.420000 11.360000 ;
      RECT  0.280000 11.360000  0.980000 11.690000 ;
      RECT  0.560000  0.330000  0.700000 11.220000 ;
      RECT  0.840000  0.000000  0.980000 11.360000 ;
      RECT  1.120000  0.000000  1.820000  0.330000 ;
      RECT  1.120000  0.330000  1.260000 11.690000 ;
      RECT  1.400000  0.470000  1.540000 11.360000 ;
      RECT  1.400000 11.360000  2.100000 11.690000 ;
      RECT  1.680000  0.330000  1.820000 11.220000 ;
      RECT  1.960000  0.000000  2.100000 11.360000 ;
      RECT  2.240000  0.000000  2.940000  0.330000 ;
      RECT  2.240000  0.330000  2.380000 11.690000 ;
      RECT  2.520000  0.470000  2.660000 11.360000 ;
      RECT  2.520000 11.360000  3.220000 11.690000 ;
      RECT  2.800000  0.330000  2.940000 11.220000 ;
      RECT  3.080000  0.000000  3.220000 11.360000 ;
      RECT  3.360000  0.000000  4.060000  0.330000 ;
      RECT  3.360000  0.330000  3.500000 11.690000 ;
      RECT  3.640000  0.470000  3.780000 11.360000 ;
      RECT  3.640000 11.360000  4.340000 11.690000 ;
      RECT  3.920000  0.330000  4.060000 11.220000 ;
      RECT  4.200000  0.000000  4.340000 11.360000 ;
      RECT  4.480000  0.000000  5.180000  0.330000 ;
      RECT  4.480000  0.330000  4.620000 11.690000 ;
      RECT  4.760000  0.470000  4.900000 11.360000 ;
      RECT  4.760000 11.360000  5.460000 11.690000 ;
      RECT  5.040000  0.330000  5.180000 11.220000 ;
      RECT  5.320000  0.000000  5.460000 11.360000 ;
      RECT  5.600000  0.000000  6.300000  0.330000 ;
      RECT  5.600000  0.330000  5.740000 11.690000 ;
      RECT  5.880000  0.470000  6.020000 11.360000 ;
      RECT  5.880000 11.360000  6.580000 11.690000 ;
      RECT  6.160000  0.330000  6.300000 11.220000 ;
      RECT  6.440000  0.000000  6.580000 11.360000 ;
      RECT  6.720000  0.000000  7.420000  0.330000 ;
      RECT  6.720000  0.330000  6.860000 11.690000 ;
      RECT  7.000000  0.470000  7.140000 11.360000 ;
      RECT  7.000000 11.360000  7.700000 11.690000 ;
      RECT  7.280000  0.330000  7.420000 11.220000 ;
      RECT  7.560000  0.000000  7.700000 11.360000 ;
      RECT  7.840000  0.000000  8.540000  0.330000 ;
      RECT  7.840000  0.330000  7.980000 11.690000 ;
      RECT  8.120000  0.470000  8.260000 11.360000 ;
      RECT  8.120000 11.360000  8.820000 11.690000 ;
      RECT  8.400000  0.330000  8.540000 11.220000 ;
      RECT  8.680000  0.000000  8.820000 11.360000 ;
      RECT  8.960000  0.000000  9.660000  0.330000 ;
      RECT  8.960000  0.330000  9.100000 11.690000 ;
      RECT  9.240000  0.470000  9.380000 11.360000 ;
      RECT  9.240000 11.360000  9.940000 11.690000 ;
      RECT  9.520000  0.330000  9.660000 11.220000 ;
      RECT  9.800000  0.000000  9.940000 11.360000 ;
      RECT 10.080000  0.000000 10.780000  0.330000 ;
      RECT 10.080000  0.330000 10.220000 11.690000 ;
      RECT 10.360000  0.470000 10.500000 11.360000 ;
      RECT 10.360000 11.360000 11.060000 11.690000 ;
      RECT 10.640000  0.330000 10.780000 11.220000 ;
      RECT 10.920000  0.000000 11.060000 11.360000 ;
      RECT 11.200000  0.000000 11.900000  0.330000 ;
      RECT 11.200000  0.330000 11.340000 11.690000 ;
      RECT 11.480000  0.470000 11.620000 11.360000 ;
      RECT 11.480000 11.360000 12.180000 11.690000 ;
      RECT 11.760000  0.330000 11.900000 11.220000 ;
      RECT 12.040000  0.000000 12.180000 11.360000 ;
      RECT 12.320000  0.000000 13.020000  0.330000 ;
      RECT 12.320000  0.330000 12.460000 11.690000 ;
      RECT 12.600000  0.470000 12.740000 11.360000 ;
      RECT 12.600000 11.360000 13.300000 11.690000 ;
      RECT 12.880000  0.330000 13.020000 11.220000 ;
      RECT 13.160000  0.000000 13.300000 11.360000 ;
      RECT 13.440000  0.000000 14.140000  0.330000 ;
      RECT 13.440000  0.330000 13.580000 11.690000 ;
      RECT 13.720000  0.470000 13.860000 11.360000 ;
      RECT 13.720000 11.360000 14.420000 11.690000 ;
      RECT 14.000000  0.330000 14.140000 11.220000 ;
      RECT 14.280000  0.000000 14.420000 11.360000 ;
      RECT 14.560000  0.000000 15.260000  0.330000 ;
      RECT 14.560000  0.330000 14.700000 11.690000 ;
      RECT 14.840000  0.470000 14.980000 11.360000 ;
      RECT 14.840000 11.360000 15.540000 11.690000 ;
      RECT 15.120000  0.330000 15.260000 11.220000 ;
      RECT 15.400000  0.000000 15.540000 11.360000 ;
      RECT 15.680000  0.000000 16.380000  0.330000 ;
      RECT 15.680000  0.330000 15.820000 11.690000 ;
      RECT 15.960000  0.470000 16.100000 11.360000 ;
      RECT 15.960000 11.360000 16.660000 11.690000 ;
      RECT 16.240000  0.330000 16.380000 11.220000 ;
      RECT 16.520000  0.000000 16.660000 11.360000 ;
      RECT 16.800000  0.000000 17.500000  0.330000 ;
      RECT 16.800000  0.330000 16.940000 11.690000 ;
      RECT 17.080000  0.470000 17.220000 11.360000 ;
      RECT 17.080000 11.360000 17.780000 11.690000 ;
      RECT 17.360000  0.330000 17.500000 11.220000 ;
      RECT 17.640000  0.000000 17.780000 11.360000 ;
      RECT 17.920000  0.000000 18.620000  0.330000 ;
      RECT 17.920000  0.330000 18.060000 11.690000 ;
      RECT 18.200000  0.470000 18.340000 11.360000 ;
      RECT 18.200000 11.360000 18.900000 11.690000 ;
      RECT 18.480000  0.330000 18.620000 11.220000 ;
      RECT 18.760000  0.000000 18.900000 11.360000 ;
      RECT 19.040000  0.000000 19.740000  0.330000 ;
      RECT 19.040000  0.330000 19.180000 11.690000 ;
      RECT 19.320000  0.470000 19.460000 11.360000 ;
      RECT 19.320000 11.360000 20.020000 11.690000 ;
      RECT 19.600000  0.330000 19.740000 11.220000 ;
      RECT 19.880000  0.000000 20.020000 11.360000 ;
      RECT 20.160000  0.000000 20.860000  0.330000 ;
      RECT 20.160000  0.330000 20.300000 11.690000 ;
      RECT 20.440000  0.470000 20.580000 11.360000 ;
      RECT 20.440000 11.360000 21.140000 11.690000 ;
      RECT 20.720000  0.330000 20.860000 11.220000 ;
      RECT 21.000000  0.000000 21.140000 11.360000 ;
      RECT 21.280000  0.000000 21.980000  0.330000 ;
      RECT 21.280000  0.330000 21.420000 11.690000 ;
      RECT 21.560000  0.470000 21.700000 11.360000 ;
      RECT 21.560000 11.360000 22.260000 11.690000 ;
      RECT 21.840000  0.330000 21.980000 11.220000 ;
      RECT 22.120000  0.000000 22.260000 11.360000 ;
      RECT 22.400000  0.000000 23.100000  0.330000 ;
      RECT 22.400000  0.330000 22.540000 11.690000 ;
      RECT 22.680000  0.470000 22.820000 11.360000 ;
      RECT 22.680000 11.360000 23.380000 11.690000 ;
      RECT 22.960000  0.330000 23.100000 11.220000 ;
      RECT 23.240000  0.000000 23.380000 11.360000 ;
      RECT 23.520000  0.000000 24.220000  0.330000 ;
      RECT 23.520000  0.330000 23.660000 11.690000 ;
      RECT 23.800000  0.470000 23.940000 11.360000 ;
      RECT 23.800000 11.360000 24.500000 11.690000 ;
      RECT 24.080000  0.330000 24.220000 11.220000 ;
      RECT 24.360000  0.000000 24.500000 11.360000 ;
      RECT 24.640000  0.000000 25.340000  0.330000 ;
      RECT 24.640000  0.330000 24.780000 11.690000 ;
      RECT 24.920000  0.470000 25.060000 11.360000 ;
      RECT 24.920000 11.360000 25.620000 11.690000 ;
      RECT 25.200000  0.330000 25.340000 11.220000 ;
      RECT 25.480000  0.000000 25.620000 11.360000 ;
      RECT 25.760000  0.000000 26.460000  0.330000 ;
      RECT 25.760000  0.330000 25.900000 11.690000 ;
      RECT 26.040000  0.470000 26.180000 11.360000 ;
      RECT 26.040000 11.360000 26.740000 11.690000 ;
      RECT 26.320000  0.330000 26.460000 11.220000 ;
      RECT 26.600000  0.000000 26.740000 11.360000 ;
      RECT 26.880000  0.000000 27.580000  0.330000 ;
      RECT 26.880000  0.330000 27.020000 11.690000 ;
      RECT 27.160000  0.470000 27.300000 11.360000 ;
      RECT 27.160000 11.360000 27.860000 11.690000 ;
      RECT 27.440000  0.330000 27.580000 11.220000 ;
      RECT 27.720000  0.000000 27.860000 11.360000 ;
      RECT 28.000000  0.000000 28.700000  0.330000 ;
      RECT 28.000000  0.330000 28.140000 11.690000 ;
      RECT 28.280000  0.470000 28.420000 11.360000 ;
      RECT 28.280000 11.360000 28.980000 11.690000 ;
      RECT 28.560000  0.330000 28.700000 11.220000 ;
      RECT 28.840000  0.000000 28.980000 11.360000 ;
      RECT 29.120000  0.000000 29.820000  0.330000 ;
      RECT 29.120000  0.330000 29.260000 11.690000 ;
      RECT 29.400000  0.470000 29.540000 11.360000 ;
      RECT 29.400000 11.360000 30.100000 11.690000 ;
      RECT 29.680000  0.330000 29.820000 11.220000 ;
      RECT 29.960000  0.000000 30.100000 11.360000 ;
      RECT 30.240000  0.000000 30.940000  0.330000 ;
      RECT 30.240000  0.330000 30.380000 11.690000 ;
      RECT 30.520000  0.470000 30.660000 11.360000 ;
      RECT 30.520000 11.360000 31.220000 11.690000 ;
      RECT 30.800000  0.330000 30.940000 11.220000 ;
      RECT 31.080000  0.000000 31.220000 11.360000 ;
      RECT 31.360000  0.000000 32.060000  0.330000 ;
      RECT 31.360000  0.330000 31.500000 11.690000 ;
      RECT 31.640000  0.470000 31.780000 11.360000 ;
      RECT 31.640000 11.360000 32.340000 11.690000 ;
      RECT 31.920000  0.330000 32.060000 11.220000 ;
      RECT 32.200000  0.000000 32.340000 11.360000 ;
      RECT 32.480000  0.000000 33.180000  0.330000 ;
      RECT 32.480000  0.330000 32.620000 11.690000 ;
      RECT 32.760000  0.470000 32.900000 11.360000 ;
      RECT 32.760000 11.360000 33.460000 11.690000 ;
      RECT 33.040000  0.330000 33.180000 11.220000 ;
      RECT 33.320000  0.000000 33.460000 11.360000 ;
      RECT 33.600000  0.000000 34.300000  0.330000 ;
      RECT 33.600000  0.330000 33.740000 11.690000 ;
      RECT 33.880000  0.470000 34.020000 11.360000 ;
      RECT 33.880000 11.360000 34.580000 11.690000 ;
      RECT 34.160000  0.330000 34.300000 11.220000 ;
      RECT 34.440000  0.000000 34.580000 11.360000 ;
      RECT 34.720000  0.000000 35.420000  0.330000 ;
      RECT 34.720000  0.330000 34.860000 11.690000 ;
      RECT 35.000000  0.470000 35.140000 11.360000 ;
      RECT 35.000000 11.360000 35.700000 11.690000 ;
      RECT 35.280000  0.330000 35.420000 11.220000 ;
      RECT 35.560000  0.000000 35.700000 11.360000 ;
      RECT 35.840000  0.000000 36.540000  0.330000 ;
      RECT 35.840000  0.330000 35.980000 11.690000 ;
      RECT 36.120000  0.470000 36.260000 11.360000 ;
      RECT 36.120000 11.360000 36.820000 11.690000 ;
      RECT 36.400000  0.330000 36.540000 11.220000 ;
      RECT 36.680000  0.000000 36.820000 11.360000 ;
      RECT 36.960000  0.000000 37.660000  0.330000 ;
      RECT 36.960000  0.330000 37.100000 11.690000 ;
      RECT 37.240000  0.470000 37.380000 11.360000 ;
      RECT 37.240000 11.360000 37.940000 11.690000 ;
      RECT 37.520000  0.330000 37.660000 11.220000 ;
      RECT 37.800000  0.000000 37.940000 11.360000 ;
      RECT 38.080000  0.000000 38.780000  0.330000 ;
      RECT 38.080000  0.330000 38.220000 11.690000 ;
      RECT 38.360000  0.470000 38.500000 11.360000 ;
      RECT 38.360000 11.360000 39.060000 11.690000 ;
      RECT 38.640000  0.330000 38.780000 11.220000 ;
      RECT 38.920000  0.000000 39.060000 11.360000 ;
      RECT 39.200000  0.000000 39.900000  0.330000 ;
      RECT 39.200000  0.330000 39.340000 11.690000 ;
      RECT 39.480000  0.470000 39.620000 11.360000 ;
      RECT 39.480000 11.360000 40.180000 11.690000 ;
      RECT 39.760000  0.330000 39.900000 11.220000 ;
      RECT 40.040000  0.000000 40.180000 11.360000 ;
      RECT 40.320000  0.000000 41.020000  0.330000 ;
      RECT 40.320000  0.330000 40.460000 11.690000 ;
      RECT 40.600000  0.470000 40.740000 11.360000 ;
      RECT 40.600000 11.360000 41.300000 11.690000 ;
      RECT 40.880000  0.330000 41.020000 11.220000 ;
      RECT 41.160000  0.000000 41.300000 11.360000 ;
      RECT 41.440000  0.000000 42.140000  0.330000 ;
      RECT 41.440000  0.330000 41.580000 11.690000 ;
      RECT 41.720000  0.470000 41.860000 11.360000 ;
      RECT 41.720000 11.360000 42.420000 11.690000 ;
      RECT 42.000000  0.330000 42.140000 11.220000 ;
      RECT 42.280000  0.000000 42.420000 11.360000 ;
      RECT 42.560000  0.000000 43.260000  0.330000 ;
      RECT 42.560000  0.330000 42.700000 11.690000 ;
      RECT 42.840000  0.470000 42.980000 11.360000 ;
      RECT 42.840000 11.360000 43.540000 11.690000 ;
      RECT 43.120000  0.330000 43.260000 11.220000 ;
      RECT 43.400000  0.000000 43.540000 11.360000 ;
      RECT 43.680000  0.000000 44.380000  0.330000 ;
      RECT 43.680000  0.330000 43.820000 11.690000 ;
      RECT 43.960000  0.470000 44.100000 11.360000 ;
      RECT 43.960000 11.360000 44.660000 11.690000 ;
      RECT 44.240000  0.330000 44.380000 11.220000 ;
      RECT 44.520000  0.000000 44.660000 11.360000 ;
      RECT 44.800000  0.000000 45.500000  0.330000 ;
      RECT 44.800000  0.330000 44.940000 11.690000 ;
      RECT 45.080000  0.470000 45.220000 11.360000 ;
      RECT 45.080000 11.360000 45.780000 11.690000 ;
      RECT 45.360000  0.330000 45.500000 11.220000 ;
      RECT 45.640000  0.000000 45.780000 11.360000 ;
      RECT 45.920000  0.000000 46.620000  0.330000 ;
      RECT 45.920000  0.330000 46.060000 11.690000 ;
      RECT 46.200000  0.470000 46.340000 11.360000 ;
      RECT 46.200000 11.360000 46.900000 11.690000 ;
      RECT 46.480000  0.330000 46.620000 11.220000 ;
      RECT 46.760000  0.000000 46.900000 11.360000 ;
      RECT 47.040000  0.000000 47.740000  0.330000 ;
      RECT 47.040000  0.330000 47.180000 11.690000 ;
      RECT 47.320000  0.470000 47.460000 11.360000 ;
      RECT 47.320000 11.360000 48.020000 11.690000 ;
      RECT 47.600000  0.330000 47.740000 11.220000 ;
      RECT 47.880000  0.000000 48.020000 11.360000 ;
      RECT 48.160000  0.000000 48.860000  0.330000 ;
      RECT 48.160000  0.330000 48.300000 11.690000 ;
      RECT 48.440000  0.470000 48.580000 11.360000 ;
      RECT 48.440000 11.360000 49.140000 11.690000 ;
      RECT 48.720000  0.330000 48.860000 11.220000 ;
      RECT 49.000000  0.000000 49.140000 11.360000 ;
      RECT 49.280000  0.000000 49.980000  0.330000 ;
      RECT 49.280000  0.330000 49.420000 11.690000 ;
      RECT 49.560000  0.470000 49.700000 11.360000 ;
      RECT 49.560000 11.360000 50.260000 11.690000 ;
      RECT 49.840000  0.330000 49.980000 11.220000 ;
      RECT 50.120000  0.000000 50.260000 11.360000 ;
      RECT 50.400000  0.000000 51.100000  0.330000 ;
      RECT 50.400000  0.330000 50.540000 11.690000 ;
      RECT 50.680000  0.470000 50.820000 11.360000 ;
      RECT 50.680000 11.360000 51.380000 11.690000 ;
      RECT 50.960000  0.330000 51.100000 11.220000 ;
      RECT 51.240000  0.000000 51.380000 11.360000 ;
      RECT 51.520000  0.000000 52.220000  0.330000 ;
      RECT 51.520000  0.330000 51.660000 11.690000 ;
      RECT 51.800000  0.470000 51.940000 11.360000 ;
      RECT 51.800000 11.360000 52.500000 11.690000 ;
      RECT 52.080000  0.330000 52.220000 11.220000 ;
      RECT 52.360000  0.000000 52.500000 11.360000 ;
      RECT 52.640000  0.000000 53.340000  0.330000 ;
      RECT 52.640000  0.330000 52.780000 11.690000 ;
      RECT 52.920000  0.470000 53.060000 11.360000 ;
      RECT 52.920000 11.360000 53.620000 11.690000 ;
      RECT 53.200000  0.330000 53.340000 11.220000 ;
      RECT 53.480000  0.000000 53.620000 11.360000 ;
      RECT 53.760000  0.000000 54.460000  0.330000 ;
      RECT 53.760000  0.330000 53.900000 11.690000 ;
      RECT 54.040000  0.470000 54.180000 11.360000 ;
      RECT 54.040000 11.360000 55.730000 11.690000 ;
      RECT 54.320000  0.330000 54.460000 11.220000 ;
      RECT 54.600000  0.000000 54.740000 11.360000 ;
      RECT 54.880000  0.000000 55.730000  0.330000 ;
      RECT 54.880000  0.330000 55.020000 11.220000 ;
      RECT 55.160000  0.470000 55.300000 11.360000 ;
      RECT 55.440000  0.330000 55.730000 11.220000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 55.730000  0.330000 ;
      RECT  0.000000  0.630000  0.300000 11.360000 ;
      RECT  0.000000 11.360000 55.730000 11.690000 ;
      RECT  0.600000  0.330000  0.900000 11.060000 ;
      RECT  1.200000  0.630000  1.500000 11.360000 ;
      RECT  1.800000  0.330000  2.100000 11.060000 ;
      RECT  2.400000  0.630000  2.700000 11.360000 ;
      RECT  3.000000  0.330000  3.300000 11.060000 ;
      RECT  3.600000  0.630000  3.900000 11.360000 ;
      RECT  4.200000  0.330000  4.500000 11.060000 ;
      RECT  4.800000  0.630000  5.100000 11.360000 ;
      RECT  5.400000  0.330000  5.700000 11.060000 ;
      RECT  6.000000  0.630000  6.300000 11.360000 ;
      RECT  6.600000  0.330000  6.900000 11.060000 ;
      RECT  7.200000  0.630000  7.500000 11.360000 ;
      RECT  7.800000  0.330000  8.100000 11.060000 ;
      RECT  8.400000  0.630000  8.700000 11.360000 ;
      RECT  9.000000  0.330000  9.300000 11.060000 ;
      RECT  9.600000  0.630000  9.900000 11.360000 ;
      RECT 10.200000  0.330000 10.500000 11.060000 ;
      RECT 10.800000  0.630000 11.100000 11.360000 ;
      RECT 11.400000  0.330000 11.700000 11.060000 ;
      RECT 12.000000  0.630000 12.300000 11.360000 ;
      RECT 12.600000  0.330000 12.900000 11.060000 ;
      RECT 13.200000  0.630000 13.500000 11.360000 ;
      RECT 13.800000  0.330000 14.100000 11.060000 ;
      RECT 14.400000  0.630000 14.700000 11.360000 ;
      RECT 15.000000  0.330000 15.300000 11.060000 ;
      RECT 15.600000  0.630000 15.900000 11.360000 ;
      RECT 16.200000  0.330000 16.500000 11.060000 ;
      RECT 16.800000  0.630000 17.100000 11.360000 ;
      RECT 17.400000  0.330000 17.700000 11.060000 ;
      RECT 18.000000  0.630000 18.300000 11.360000 ;
      RECT 18.600000  0.330000 18.900000 11.060000 ;
      RECT 19.200000  0.630000 19.500000 11.360000 ;
      RECT 19.800000  0.330000 20.100000 11.060000 ;
      RECT 20.400000  0.630000 20.700000 11.360000 ;
      RECT 21.000000  0.330000 21.300000 11.060000 ;
      RECT 21.600000  0.630000 21.900000 11.360000 ;
      RECT 22.200000  0.330000 22.500000 11.060000 ;
      RECT 22.800000  0.630000 23.100000 11.360000 ;
      RECT 23.400000  0.330000 23.700000 11.060000 ;
      RECT 24.000000  0.630000 24.300000 11.360000 ;
      RECT 24.600000  0.330000 24.900000 11.060000 ;
      RECT 25.200000  0.630000 25.500000 11.360000 ;
      RECT 25.800000  0.330000 26.100000 11.060000 ;
      RECT 26.400000  0.630000 26.700000 11.360000 ;
      RECT 27.000000  0.330000 27.300000 11.060000 ;
      RECT 27.600000  0.630000 27.900000 11.360000 ;
      RECT 28.200000  0.330000 28.500000 11.060000 ;
      RECT 28.800000  0.630000 29.100000 11.360000 ;
      RECT 29.400000  0.330000 29.700000 11.060000 ;
      RECT 30.000000  0.630000 30.300000 11.360000 ;
      RECT 30.600000  0.330000 30.900000 11.060000 ;
      RECT 31.200000  0.630000 31.500000 11.360000 ;
      RECT 31.800000  0.330000 32.100000 11.060000 ;
      RECT 32.400000  0.630000 32.700000 11.360000 ;
      RECT 33.000000  0.330000 33.300000 11.060000 ;
      RECT 33.600000  0.630000 33.900000 11.360000 ;
      RECT 34.200000  0.330000 34.500000 11.060000 ;
      RECT 34.800000  0.630000 35.100000 11.360000 ;
      RECT 35.400000  0.330000 35.700000 11.060000 ;
      RECT 36.000000  0.630000 36.300000 11.360000 ;
      RECT 36.600000  0.330000 36.900000 11.060000 ;
      RECT 37.200000  0.630000 37.500000 11.360000 ;
      RECT 37.800000  0.330000 38.100000 11.060000 ;
      RECT 38.400000  0.630000 38.700000 11.360000 ;
      RECT 39.000000  0.330000 39.300000 11.060000 ;
      RECT 39.600000  0.630000 39.900000 11.360000 ;
      RECT 40.200000  0.330000 40.500000 11.060000 ;
      RECT 40.800000  0.630000 41.100000 11.360000 ;
      RECT 41.400000  0.330000 41.700000 11.060000 ;
      RECT 42.000000  0.630000 42.300000 11.360000 ;
      RECT 42.600000  0.330000 42.900000 11.060000 ;
      RECT 43.200000  0.630000 43.500000 11.360000 ;
      RECT 43.800000  0.330000 44.100000 11.060000 ;
      RECT 44.400000  0.630000 44.700000 11.360000 ;
      RECT 45.000000  0.330000 45.300000 11.060000 ;
      RECT 45.600000  0.630000 45.900000 11.360000 ;
      RECT 46.200000  0.330000 46.500000 11.060000 ;
      RECT 46.800000  0.630000 47.100000 11.360000 ;
      RECT 47.400000  0.330000 47.700000 11.060000 ;
      RECT 48.000000  0.630000 48.300000 11.360000 ;
      RECT 48.600000  0.330000 48.900000 11.060000 ;
      RECT 49.200000  0.630000 49.500000 11.360000 ;
      RECT 49.800000  0.330000 50.100000 11.060000 ;
      RECT 50.400000  0.630000 50.700000 11.360000 ;
      RECT 51.000000  0.330000 51.300000 11.060000 ;
      RECT 51.600000  0.630000 51.900000 11.360000 ;
      RECT 52.200000  0.330000 52.500000 11.060000 ;
      RECT 52.800000  0.630000 53.100000 11.360000 ;
      RECT 53.400000  0.330000 53.700000 11.060000 ;
      RECT 54.000000  0.630000 54.300000 11.360000 ;
      RECT 54.600000  0.330000 54.900000 11.060000 ;
      RECT 55.200000  0.630000 55.730000 11.360000 ;
    LAYER met4 ;
      RECT  0.000000  0.000000 55.730000  0.330000 ;
      RECT  0.000000  0.330000  0.300000 11.060000 ;
      RECT  0.000000 11.360000 55.730000 11.690000 ;
      RECT  0.600000  0.630000  0.900000  9.990000 ;
      RECT  0.600000  9.990000  2.100000 11.360000 ;
      RECT  1.200000  0.330000  2.700000  1.700000 ;
      RECT  1.200000  1.700000  1.500000  9.690000 ;
      RECT  1.800000  2.000000  2.100000  9.990000 ;
      RECT  2.400000  1.700000  2.700000 11.060000 ;
      RECT  3.000000  0.630000  3.300000 11.360000 ;
      RECT  3.600000  0.330000  3.900000 11.060000 ;
      RECT  4.200000  0.630000  4.500000 11.360000 ;
      RECT  4.800000  0.330000  5.100000 11.060000 ;
      RECT  5.400000  0.630000  5.700000 11.360000 ;
      RECT  6.000000  0.330000  6.300000 11.060000 ;
      RECT  6.600000  0.630000  6.900000 11.360000 ;
      RECT  7.200000  0.330000  7.500000 11.060000 ;
      RECT  7.800000  0.630000  8.100000  9.990000 ;
      RECT  7.800000  9.990000  9.300000 11.360000 ;
      RECT  8.400000  0.330000  9.900000  1.700000 ;
      RECT  8.400000  1.700000  8.700000  9.690000 ;
      RECT  9.000000  2.000000  9.300000  9.990000 ;
      RECT  9.600000  1.700000  9.900000 11.060000 ;
      RECT 10.200000  0.630000 10.500000 11.360000 ;
      RECT 10.800000  0.330000 11.100000 11.060000 ;
      RECT 11.400000  0.630000 11.700000 11.360000 ;
      RECT 12.000000  0.330000 12.300000 11.060000 ;
      RECT 12.600000  0.630000 12.900000 11.360000 ;
      RECT 13.200000  0.330000 13.500000 11.060000 ;
      RECT 13.800000  0.630000 14.100000 11.360000 ;
      RECT 14.400000  0.330000 14.700000 11.060000 ;
      RECT 15.000000  0.630000 15.300000  9.990000 ;
      RECT 15.000000  9.990000 16.500000 11.360000 ;
      RECT 15.600000  0.330000 17.100000  1.700000 ;
      RECT 15.600000  1.700000 15.900000  9.690000 ;
      RECT 16.200000  2.000000 16.500000  9.990000 ;
      RECT 16.800000  1.700000 17.100000 11.060000 ;
      RECT 17.400000  0.630000 17.700000 11.360000 ;
      RECT 18.000000  0.330000 18.300000 11.060000 ;
      RECT 18.600000  0.630000 18.900000 11.360000 ;
      RECT 19.200000  0.330000 19.500000 11.060000 ;
      RECT 19.800000  0.630000 20.100000 11.360000 ;
      RECT 20.400000  0.330000 20.700000 11.060000 ;
      RECT 21.000000  0.630000 21.300000 11.360000 ;
      RECT 21.600000  0.330000 21.900000 11.060000 ;
      RECT 22.200000  0.630000 22.500000  9.990000 ;
      RECT 22.200000  9.990000 23.700000 11.360000 ;
      RECT 22.800000  0.330000 24.300000  1.700000 ;
      RECT 22.800000  1.700000 23.100000  9.690000 ;
      RECT 23.400000  2.000000 23.700000  9.990000 ;
      RECT 24.000000  1.700000 24.300000 11.060000 ;
      RECT 24.600000  0.630000 24.900000 11.360000 ;
      RECT 25.200000  0.330000 25.500000 11.060000 ;
      RECT 25.800000  0.630000 26.100000 11.360000 ;
      RECT 26.400000  0.330000 26.700000 11.060000 ;
      RECT 27.000000  0.630000 27.300000 11.360000 ;
      RECT 27.600000  0.330000 27.900000 11.060000 ;
      RECT 28.200000  0.630000 28.500000 11.360000 ;
      RECT 28.800000  0.330000 29.100000 11.060000 ;
      RECT 29.400000  0.630000 29.700000  9.990000 ;
      RECT 29.400000  9.990000 30.900000 11.360000 ;
      RECT 30.000000  0.330000 31.500000  1.700000 ;
      RECT 30.000000  1.700000 30.300000  9.690000 ;
      RECT 30.600000  2.000000 30.900000  9.990000 ;
      RECT 31.200000  1.700000 31.500000 11.060000 ;
      RECT 31.800000  0.630000 32.100000 11.360000 ;
      RECT 32.400000  0.330000 32.700000 11.060000 ;
      RECT 33.000000  0.630000 33.300000 11.360000 ;
      RECT 33.600000  0.330000 33.900000 11.060000 ;
      RECT 34.200000  0.630000 34.500000 11.360000 ;
      RECT 34.800000  0.330000 35.100000 11.060000 ;
      RECT 35.400000  0.630000 35.700000 11.360000 ;
      RECT 36.000000  0.330000 36.300000 11.060000 ;
      RECT 36.600000  0.630000 36.900000  9.990000 ;
      RECT 36.600000  9.990000 38.100000 11.360000 ;
      RECT 37.200000  0.330000 38.700000  1.700000 ;
      RECT 37.200000  1.700000 37.500000  9.690000 ;
      RECT 37.800000  2.000000 38.100000  9.990000 ;
      RECT 38.400000  1.700000 38.700000 11.060000 ;
      RECT 39.000000  0.630000 39.300000 11.360000 ;
      RECT 39.600000  0.330000 39.900000 11.060000 ;
      RECT 40.200000  0.630000 40.500000 11.360000 ;
      RECT 40.800000  0.330000 41.100000 11.060000 ;
      RECT 41.400000  0.630000 41.700000 11.360000 ;
      RECT 42.000000  0.330000 42.300000 11.060000 ;
      RECT 42.600000  0.630000 42.900000 11.360000 ;
      RECT 43.200000  0.330000 43.500000 11.060000 ;
      RECT 43.800000  0.630000 44.100000  9.990000 ;
      RECT 43.800000  9.990000 45.300000 11.360000 ;
      RECT 44.400000  0.330000 45.900000  1.700000 ;
      RECT 44.400000  1.700000 44.700000  9.690000 ;
      RECT 45.000000  2.000000 45.300000  9.990000 ;
      RECT 45.600000  1.700000 45.900000 11.060000 ;
      RECT 46.200000  0.630000 46.500000 11.360000 ;
      RECT 46.800000  0.330000 47.100000 11.060000 ;
      RECT 47.400000  0.630000 47.700000 11.360000 ;
      RECT 48.000000  0.330000 48.300000 11.060000 ;
      RECT 48.600000  0.630000 48.900000 11.360000 ;
      RECT 49.200000  0.330000 49.500000 11.060000 ;
      RECT 49.800000  0.630000 50.100000 11.360000 ;
      RECT 50.400000  0.330000 50.700000 11.060000 ;
      RECT 51.000000  0.630000 51.300000  9.990000 ;
      RECT 51.000000  9.990000 52.500000 11.360000 ;
      RECT 51.600000  0.330000 53.100000  1.700000 ;
      RECT 51.600000  1.700000 51.900000  9.690000 ;
      RECT 52.200000  2.000000 52.500000  9.990000 ;
      RECT 52.800000  1.700000 53.100000 11.060000 ;
      RECT 53.400000  0.630000 53.700000 11.360000 ;
      RECT 54.000000  0.330000 54.300000 11.060000 ;
      RECT 54.600000  0.630000 54.900000 11.360000 ;
      RECT 55.200000  0.330000 55.730000 11.060000 ;
    LAYER met5 ;
      RECT  0.000000 0.400000 54.930000  2.000000 ;
      RECT  0.000000 3.600000  1.600000  9.690000 ;
      RECT  0.000000 9.690000 54.930000 11.290000 ;
      RECT  3.200000 2.000000  4.800000  8.090000 ;
      RECT  6.400000 3.600000  8.000000  9.690000 ;
      RECT  9.600000 2.000000 11.200000  8.090000 ;
      RECT 12.800000 3.600000 14.400000  9.690000 ;
      RECT 16.000000 2.000000 17.600000  8.090000 ;
      RECT 19.200000 3.600000 20.800000  9.690000 ;
      RECT 22.400000 2.000000 24.000000  8.090000 ;
      RECT 25.600000 3.600000 27.200000  9.690000 ;
      RECT 28.800000 2.000000 30.400000  8.090000 ;
      RECT 32.000000 3.600000 33.600000  9.690000 ;
      RECT 35.200000 2.000000 36.800000  8.090000 ;
      RECT 38.400000 3.600000 40.000000  9.690000 ;
      RECT 41.600000 2.000000 43.200000  8.090000 ;
      RECT 44.800000 3.600000 46.400000  9.690000 ;
      RECT 48.000000 2.000000 49.600000  8.090000 ;
      RECT 51.200000 3.600000 54.930000  9.690000 ;
    LAYER via ;
      RECT  0.120000  0.035000  0.380000  0.295000 ;
      RECT  0.340000 11.395000  0.600000 11.655000 ;
      RECT  0.440000  0.035000  0.700000  0.295000 ;
      RECT  0.660000 11.395000  0.920000 11.655000 ;
      RECT  1.180000  0.035000  1.440000  0.295000 ;
      RECT  1.460000 11.395000  1.720000 11.655000 ;
      RECT  1.500000  0.035000  1.760000  0.295000 ;
      RECT  1.780000 11.395000  2.040000 11.655000 ;
      RECT  2.300000  0.035000  2.560000  0.295000 ;
      RECT  2.580000 11.395000  2.840000 11.655000 ;
      RECT  2.620000  0.035000  2.880000  0.295000 ;
      RECT  2.900000 11.395000  3.160000 11.655000 ;
      RECT  3.420000  0.035000  3.680000  0.295000 ;
      RECT  3.700000 11.395000  3.960000 11.655000 ;
      RECT  3.740000  0.035000  4.000000  0.295000 ;
      RECT  4.020000 11.395000  4.280000 11.655000 ;
      RECT  4.540000  0.035000  4.800000  0.295000 ;
      RECT  4.820000 11.395000  5.080000 11.655000 ;
      RECT  4.860000  0.035000  5.120000  0.295000 ;
      RECT  5.140000 11.395000  5.400000 11.655000 ;
      RECT  5.660000  0.035000  5.920000  0.295000 ;
      RECT  5.940000 11.395000  6.200000 11.655000 ;
      RECT  5.980000  0.035000  6.240000  0.295000 ;
      RECT  6.260000 11.395000  6.520000 11.655000 ;
      RECT  6.780000  0.035000  7.040000  0.295000 ;
      RECT  7.060000 11.395000  7.320000 11.655000 ;
      RECT  7.100000  0.035000  7.360000  0.295000 ;
      RECT  7.380000 11.395000  7.640000 11.655000 ;
      RECT  7.900000  0.035000  8.160000  0.295000 ;
      RECT  8.180000 11.395000  8.440000 11.655000 ;
      RECT  8.220000  0.035000  8.480000  0.295000 ;
      RECT  8.500000 11.395000  8.760000 11.655000 ;
      RECT  9.020000  0.035000  9.280000  0.295000 ;
      RECT  9.300000 11.395000  9.560000 11.655000 ;
      RECT  9.340000  0.035000  9.600000  0.295000 ;
      RECT  9.620000 11.395000  9.880000 11.655000 ;
      RECT 10.140000  0.035000 10.400000  0.295000 ;
      RECT 10.420000 11.395000 10.680000 11.655000 ;
      RECT 10.460000  0.035000 10.720000  0.295000 ;
      RECT 10.740000 11.395000 11.000000 11.655000 ;
      RECT 11.260000  0.035000 11.520000  0.295000 ;
      RECT 11.540000 11.395000 11.800000 11.655000 ;
      RECT 11.580000  0.035000 11.840000  0.295000 ;
      RECT 11.860000 11.395000 12.120000 11.655000 ;
      RECT 12.380000  0.035000 12.640000  0.295000 ;
      RECT 12.660000 11.395000 12.920000 11.655000 ;
      RECT 12.700000  0.035000 12.960000  0.295000 ;
      RECT 12.980000 11.395000 13.240000 11.655000 ;
      RECT 13.500000  0.035000 13.760000  0.295000 ;
      RECT 13.780000 11.395000 14.040000 11.655000 ;
      RECT 13.820000  0.035000 14.080000  0.295000 ;
      RECT 14.100000 11.395000 14.360000 11.655000 ;
      RECT 14.620000  0.035000 14.880000  0.295000 ;
      RECT 14.900000 11.395000 15.160000 11.655000 ;
      RECT 14.940000  0.035000 15.200000  0.295000 ;
      RECT 15.220000 11.395000 15.480000 11.655000 ;
      RECT 15.740000  0.035000 16.000000  0.295000 ;
      RECT 16.020000 11.395000 16.280000 11.655000 ;
      RECT 16.060000  0.035000 16.320000  0.295000 ;
      RECT 16.340000 11.395000 16.600000 11.655000 ;
      RECT 16.860000  0.035000 17.120000  0.295000 ;
      RECT 17.140000 11.395000 17.400000 11.655000 ;
      RECT 17.180000  0.035000 17.440000  0.295000 ;
      RECT 17.460000 11.395000 17.720000 11.655000 ;
      RECT 17.980000  0.035000 18.240000  0.295000 ;
      RECT 18.260000 11.395000 18.520000 11.655000 ;
      RECT 18.300000  0.035000 18.560000  0.295000 ;
      RECT 18.580000 11.395000 18.840000 11.655000 ;
      RECT 19.100000  0.035000 19.360000  0.295000 ;
      RECT 19.380000 11.395000 19.640000 11.655000 ;
      RECT 19.420000  0.035000 19.680000  0.295000 ;
      RECT 19.700000 11.395000 19.960000 11.655000 ;
      RECT 20.220000  0.035000 20.480000  0.295000 ;
      RECT 20.500000 11.395000 20.760000 11.655000 ;
      RECT 20.540000  0.035000 20.800000  0.295000 ;
      RECT 20.820000 11.395000 21.080000 11.655000 ;
      RECT 21.340000  0.035000 21.600000  0.295000 ;
      RECT 21.620000 11.395000 21.880000 11.655000 ;
      RECT 21.660000  0.035000 21.920000  0.295000 ;
      RECT 21.940000 11.395000 22.200000 11.655000 ;
      RECT 22.460000  0.035000 22.720000  0.295000 ;
      RECT 22.740000 11.395000 23.000000 11.655000 ;
      RECT 22.780000  0.035000 23.040000  0.295000 ;
      RECT 23.060000 11.395000 23.320000 11.655000 ;
      RECT 23.580000  0.035000 23.840000  0.295000 ;
      RECT 23.860000 11.395000 24.120000 11.655000 ;
      RECT 23.900000  0.035000 24.160000  0.295000 ;
      RECT 24.180000 11.395000 24.440000 11.655000 ;
      RECT 24.700000  0.035000 24.960000  0.295000 ;
      RECT 24.980000 11.395000 25.240000 11.655000 ;
      RECT 25.020000  0.035000 25.280000  0.295000 ;
      RECT 25.300000 11.395000 25.560000 11.655000 ;
      RECT 25.820000  0.035000 26.080000  0.295000 ;
      RECT 26.100000 11.395000 26.360000 11.655000 ;
      RECT 26.140000  0.035000 26.400000  0.295000 ;
      RECT 26.420000 11.395000 26.680000 11.655000 ;
      RECT 26.940000  0.035000 27.200000  0.295000 ;
      RECT 27.220000 11.395000 27.480000 11.655000 ;
      RECT 27.260000  0.035000 27.520000  0.295000 ;
      RECT 27.540000 11.395000 27.800000 11.655000 ;
      RECT 28.060000  0.035000 28.320000  0.295000 ;
      RECT 28.340000 11.395000 28.600000 11.655000 ;
      RECT 28.380000  0.035000 28.640000  0.295000 ;
      RECT 28.660000 11.395000 28.920000 11.655000 ;
      RECT 29.180000  0.035000 29.440000  0.295000 ;
      RECT 29.460000 11.395000 29.720000 11.655000 ;
      RECT 29.500000  0.035000 29.760000  0.295000 ;
      RECT 29.780000 11.395000 30.040000 11.655000 ;
      RECT 30.300000  0.035000 30.560000  0.295000 ;
      RECT 30.580000 11.395000 30.840000 11.655000 ;
      RECT 30.620000  0.035000 30.880000  0.295000 ;
      RECT 30.900000 11.395000 31.160000 11.655000 ;
      RECT 31.420000  0.035000 31.680000  0.295000 ;
      RECT 31.700000 11.395000 31.960000 11.655000 ;
      RECT 31.740000  0.035000 32.000000  0.295000 ;
      RECT 32.020000 11.395000 32.280000 11.655000 ;
      RECT 32.540000  0.035000 32.800000  0.295000 ;
      RECT 32.820000 11.395000 33.080000 11.655000 ;
      RECT 32.860000  0.035000 33.120000  0.295000 ;
      RECT 33.140000 11.395000 33.400000 11.655000 ;
      RECT 33.660000  0.035000 33.920000  0.295000 ;
      RECT 33.940000 11.395000 34.200000 11.655000 ;
      RECT 33.980000  0.035000 34.240000  0.295000 ;
      RECT 34.260000 11.395000 34.520000 11.655000 ;
      RECT 34.780000  0.035000 35.040000  0.295000 ;
      RECT 35.060000 11.395000 35.320000 11.655000 ;
      RECT 35.100000  0.035000 35.360000  0.295000 ;
      RECT 35.380000 11.395000 35.640000 11.655000 ;
      RECT 35.900000  0.035000 36.160000  0.295000 ;
      RECT 36.180000 11.395000 36.440000 11.655000 ;
      RECT 36.220000  0.035000 36.480000  0.295000 ;
      RECT 36.500000 11.395000 36.760000 11.655000 ;
      RECT 37.020000  0.035000 37.280000  0.295000 ;
      RECT 37.300000 11.395000 37.560000 11.655000 ;
      RECT 37.340000  0.035000 37.600000  0.295000 ;
      RECT 37.620000 11.395000 37.880000 11.655000 ;
      RECT 38.140000  0.035000 38.400000  0.295000 ;
      RECT 38.420000 11.395000 38.680000 11.655000 ;
      RECT 38.460000  0.035000 38.720000  0.295000 ;
      RECT 38.740000 11.395000 39.000000 11.655000 ;
      RECT 39.260000  0.035000 39.520000  0.295000 ;
      RECT 39.540000 11.395000 39.800000 11.655000 ;
      RECT 39.580000  0.035000 39.840000  0.295000 ;
      RECT 39.860000 11.395000 40.120000 11.655000 ;
      RECT 40.380000  0.035000 40.640000  0.295000 ;
      RECT 40.660000 11.395000 40.920000 11.655000 ;
      RECT 40.700000  0.035000 40.960000  0.295000 ;
      RECT 40.980000 11.395000 41.240000 11.655000 ;
      RECT 41.500000  0.035000 41.760000  0.295000 ;
      RECT 41.780000 11.395000 42.040000 11.655000 ;
      RECT 41.820000  0.035000 42.080000  0.295000 ;
      RECT 42.100000 11.395000 42.360000 11.655000 ;
      RECT 42.620000  0.035000 42.880000  0.295000 ;
      RECT 42.900000 11.395000 43.160000 11.655000 ;
      RECT 42.940000  0.035000 43.200000  0.295000 ;
      RECT 43.220000 11.395000 43.480000 11.655000 ;
      RECT 43.740000  0.035000 44.000000  0.295000 ;
      RECT 44.020000 11.395000 44.280000 11.655000 ;
      RECT 44.060000  0.035000 44.320000  0.295000 ;
      RECT 44.340000 11.395000 44.600000 11.655000 ;
      RECT 44.860000  0.035000 45.120000  0.295000 ;
      RECT 45.140000 11.395000 45.400000 11.655000 ;
      RECT 45.180000  0.035000 45.440000  0.295000 ;
      RECT 45.460000 11.395000 45.720000 11.655000 ;
      RECT 45.980000  0.035000 46.240000  0.295000 ;
      RECT 46.260000 11.395000 46.520000 11.655000 ;
      RECT 46.300000  0.035000 46.560000  0.295000 ;
      RECT 46.580000 11.395000 46.840000 11.655000 ;
      RECT 47.100000  0.035000 47.360000  0.295000 ;
      RECT 47.380000 11.395000 47.640000 11.655000 ;
      RECT 47.420000  0.035000 47.680000  0.295000 ;
      RECT 47.700000 11.395000 47.960000 11.655000 ;
      RECT 48.220000  0.035000 48.480000  0.295000 ;
      RECT 48.500000 11.395000 48.760000 11.655000 ;
      RECT 48.540000  0.035000 48.800000  0.295000 ;
      RECT 48.820000 11.395000 49.080000 11.655000 ;
      RECT 49.340000  0.035000 49.600000  0.295000 ;
      RECT 49.620000 11.395000 49.880000 11.655000 ;
      RECT 49.660000  0.035000 49.920000  0.295000 ;
      RECT 49.940000 11.395000 50.200000 11.655000 ;
      RECT 50.460000  0.035000 50.720000  0.295000 ;
      RECT 50.740000 11.395000 51.000000 11.655000 ;
      RECT 50.780000  0.035000 51.040000  0.295000 ;
      RECT 51.060000 11.395000 51.320000 11.655000 ;
      RECT 51.580000  0.035000 51.840000  0.295000 ;
      RECT 51.860000 11.395000 52.120000 11.655000 ;
      RECT 51.900000  0.035000 52.160000  0.295000 ;
      RECT 52.180000 11.395000 52.440000 11.655000 ;
      RECT 52.700000  0.035000 52.960000  0.295000 ;
      RECT 52.980000 11.395000 53.240000 11.655000 ;
      RECT 53.020000  0.035000 53.280000  0.295000 ;
      RECT 53.300000 11.395000 53.560000 11.655000 ;
      RECT 53.820000  0.035000 54.080000  0.295000 ;
      RECT 54.100000 11.395000 54.360000 11.655000 ;
      RECT 54.140000  0.035000 54.400000  0.295000 ;
      RECT 54.420000 11.395000 54.680000 11.655000 ;
      RECT 54.940000  0.035000 55.200000  0.295000 ;
      RECT 55.260000  0.035000 55.520000  0.295000 ;
    LAYER via2 ;
      RECT  0.210000  0.025000  0.490000  0.305000 ;
      RECT  0.490000 11.385000  0.770000 11.665000 ;
      RECT  1.330000  0.025000  1.610000  0.305000 ;
      RECT  1.610000 11.385000  1.890000 11.665000 ;
      RECT  2.450000  0.025000  2.730000  0.305000 ;
      RECT  2.730000 11.385000  3.010000 11.665000 ;
      RECT  3.570000  0.025000  3.850000  0.305000 ;
      RECT  3.850000 11.385000  4.130000 11.665000 ;
      RECT  4.690000  0.025000  4.970000  0.305000 ;
      RECT  4.970000 11.385000  5.250000 11.665000 ;
      RECT  5.810000  0.025000  6.090000  0.305000 ;
      RECT  6.090000 11.385000  6.370000 11.665000 ;
      RECT  6.930000  0.025000  7.210000  0.305000 ;
      RECT  7.210000 11.385000  7.490000 11.665000 ;
      RECT  8.050000  0.025000  8.330000  0.305000 ;
      RECT  8.330000 11.385000  8.610000 11.665000 ;
      RECT  9.170000  0.025000  9.450000  0.305000 ;
      RECT  9.450000 11.385000  9.730000 11.665000 ;
      RECT 10.290000  0.025000 10.570000  0.305000 ;
      RECT 10.570000 11.385000 10.850000 11.665000 ;
      RECT 11.410000  0.025000 11.690000  0.305000 ;
      RECT 11.690000 11.385000 11.970000 11.665000 ;
      RECT 12.530000  0.025000 12.810000  0.305000 ;
      RECT 12.810000 11.385000 13.090000 11.665000 ;
      RECT 13.650000  0.025000 13.930000  0.305000 ;
      RECT 13.930000 11.385000 14.210000 11.665000 ;
      RECT 14.770000  0.025000 15.050000  0.305000 ;
      RECT 15.050000 11.385000 15.330000 11.665000 ;
      RECT 15.890000  0.025000 16.170000  0.305000 ;
      RECT 16.170000 11.385000 16.450000 11.665000 ;
      RECT 17.010000  0.025000 17.290000  0.305000 ;
      RECT 17.290000 11.385000 17.570000 11.665000 ;
      RECT 18.130000  0.025000 18.410000  0.305000 ;
      RECT 18.410000 11.385000 18.690000 11.665000 ;
      RECT 19.250000  0.025000 19.530000  0.305000 ;
      RECT 19.530000 11.385000 19.810000 11.665000 ;
      RECT 20.370000  0.025000 20.650000  0.305000 ;
      RECT 20.650000 11.385000 20.930000 11.665000 ;
      RECT 21.490000  0.025000 21.770000  0.305000 ;
      RECT 21.770000 11.385000 22.050000 11.665000 ;
      RECT 22.610000  0.025000 22.890000  0.305000 ;
      RECT 22.890000 11.385000 23.170000 11.665000 ;
      RECT 23.730000  0.025000 24.010000  0.305000 ;
      RECT 24.010000 11.385000 24.290000 11.665000 ;
      RECT 24.850000  0.025000 25.130000  0.305000 ;
      RECT 25.130000 11.385000 25.410000 11.665000 ;
      RECT 25.970000  0.025000 26.250000  0.305000 ;
      RECT 26.250000 11.385000 26.530000 11.665000 ;
      RECT 27.090000  0.025000 27.370000  0.305000 ;
      RECT 27.370000 11.385000 27.650000 11.665000 ;
      RECT 28.210000  0.025000 28.490000  0.305000 ;
      RECT 28.490000 11.385000 28.770000 11.665000 ;
      RECT 29.330000  0.025000 29.610000  0.305000 ;
      RECT 29.610000 11.385000 29.890000 11.665000 ;
      RECT 30.450000  0.025000 30.730000  0.305000 ;
      RECT 30.730000 11.385000 31.010000 11.665000 ;
      RECT 31.570000  0.025000 31.850000  0.305000 ;
      RECT 31.850000 11.385000 32.130000 11.665000 ;
      RECT 32.690000  0.025000 32.970000  0.305000 ;
      RECT 32.970000 11.385000 33.250000 11.665000 ;
      RECT 33.810000  0.025000 34.090000  0.305000 ;
      RECT 34.090000 11.385000 34.370000 11.665000 ;
      RECT 34.930000  0.025000 35.210000  0.305000 ;
      RECT 35.210000 11.385000 35.490000 11.665000 ;
      RECT 36.050000  0.025000 36.330000  0.305000 ;
      RECT 36.330000 11.385000 36.610000 11.665000 ;
      RECT 37.170000  0.025000 37.450000  0.305000 ;
      RECT 37.450000 11.385000 37.730000 11.665000 ;
      RECT 38.290000  0.025000 38.570000  0.305000 ;
      RECT 38.570000 11.385000 38.850000 11.665000 ;
      RECT 39.410000  0.025000 39.690000  0.305000 ;
      RECT 39.690000 11.385000 39.970000 11.665000 ;
      RECT 40.530000  0.025000 40.810000  0.305000 ;
      RECT 40.810000 11.385000 41.090000 11.665000 ;
      RECT 41.650000  0.025000 41.930000  0.305000 ;
      RECT 41.930000 11.385000 42.210000 11.665000 ;
      RECT 42.770000  0.025000 43.050000  0.305000 ;
      RECT 43.050000 11.385000 43.330000 11.665000 ;
      RECT 43.890000  0.025000 44.170000  0.305000 ;
      RECT 44.170000 11.385000 44.450000 11.665000 ;
      RECT 45.010000  0.025000 45.290000  0.305000 ;
      RECT 45.290000 11.385000 45.570000 11.665000 ;
      RECT 46.130000  0.025000 46.410000  0.305000 ;
      RECT 46.410000 11.385000 46.690000 11.665000 ;
      RECT 47.250000  0.025000 47.530000  0.305000 ;
      RECT 47.530000 11.385000 47.810000 11.665000 ;
      RECT 48.370000  0.025000 48.650000  0.305000 ;
      RECT 48.650000 11.385000 48.930000 11.665000 ;
      RECT 49.490000  0.025000 49.770000  0.305000 ;
      RECT 49.770000 11.385000 50.050000 11.665000 ;
      RECT 50.610000  0.025000 50.890000  0.305000 ;
      RECT 50.890000 11.385000 51.170000 11.665000 ;
      RECT 51.730000  0.025000 52.010000  0.305000 ;
      RECT 52.010000 11.385000 52.290000 11.665000 ;
      RECT 52.850000  0.025000 53.130000  0.305000 ;
      RECT 53.130000 11.385000 53.410000 11.665000 ;
      RECT 53.970000  0.025000 54.250000  0.305000 ;
      RECT 54.250000 11.385000 54.530000 11.665000 ;
      RECT 55.090000  0.025000 55.370000  0.305000 ;
    LAYER via3 ;
      RECT  0.140000  0.005000  0.460000  0.325000 ;
      RECT  0.140000 11.365000  0.460000 11.685000 ;
      RECT  0.540000  0.005000  0.860000  0.325000 ;
      RECT  0.540000 11.365000  0.860000 11.685000 ;
      RECT  0.940000  0.005000  1.260000  0.325000 ;
      RECT  0.940000 11.365000  1.260000 11.685000 ;
      RECT  1.340000  0.005000  1.660000  0.325000 ;
      RECT  1.340000 11.365000  1.660000 11.685000 ;
      RECT  1.740000  0.005000  2.060000  0.325000 ;
      RECT  1.740000 11.365000  2.060000 11.685000 ;
      RECT  2.140000  0.005000  2.460000  0.325000 ;
      RECT  2.140000 11.365000  2.460000 11.685000 ;
      RECT  2.540000  0.005000  2.860000  0.325000 ;
      RECT  2.540000 11.365000  2.860000 11.685000 ;
      RECT  2.940000  0.005000  3.260000  0.325000 ;
      RECT  2.940000 11.365000  3.260000 11.685000 ;
      RECT  3.340000  0.005000  3.660000  0.325000 ;
      RECT  3.340000 11.365000  3.660000 11.685000 ;
      RECT  3.740000  0.005000  4.060000  0.325000 ;
      RECT  3.740000 11.365000  4.060000 11.685000 ;
      RECT  4.140000  0.005000  4.460000  0.325000 ;
      RECT  4.140000 11.365000  4.460000 11.685000 ;
      RECT  4.540000  0.005000  4.860000  0.325000 ;
      RECT  4.540000 11.365000  4.860000 11.685000 ;
      RECT  4.940000  0.005000  5.260000  0.325000 ;
      RECT  4.940000 11.365000  5.260000 11.685000 ;
      RECT  5.340000  0.005000  5.660000  0.325000 ;
      RECT  5.340000 11.365000  5.660000 11.685000 ;
      RECT  5.740000  0.005000  6.060000  0.325000 ;
      RECT  5.740000 11.365000  6.060000 11.685000 ;
      RECT  6.140000  0.005000  6.460000  0.325000 ;
      RECT  6.140000 11.365000  6.460000 11.685000 ;
      RECT  6.540000  0.005000  6.860000  0.325000 ;
      RECT  6.540000 11.365000  6.860000 11.685000 ;
      RECT  6.940000  0.005000  7.260000  0.325000 ;
      RECT  6.940000 11.365000  7.260000 11.685000 ;
      RECT  7.340000  0.005000  7.660000  0.325000 ;
      RECT  7.340000 11.365000  7.660000 11.685000 ;
      RECT  7.740000  0.005000  8.060000  0.325000 ;
      RECT  7.740000 11.365000  8.060000 11.685000 ;
      RECT  8.140000  0.005000  8.460000  0.325000 ;
      RECT  8.140000 11.365000  8.460000 11.685000 ;
      RECT  8.540000  0.005000  8.860000  0.325000 ;
      RECT  8.540000 11.365000  8.860000 11.685000 ;
      RECT  8.940000  0.005000  9.260000  0.325000 ;
      RECT  8.940000 11.365000  9.260000 11.685000 ;
      RECT  9.340000  0.005000  9.660000  0.325000 ;
      RECT  9.340000 11.365000  9.660000 11.685000 ;
      RECT  9.740000  0.005000 10.060000  0.325000 ;
      RECT  9.740000 11.365000 10.060000 11.685000 ;
      RECT 10.140000  0.005000 10.460000  0.325000 ;
      RECT 10.140000 11.365000 10.460000 11.685000 ;
      RECT 10.540000  0.005000 10.860000  0.325000 ;
      RECT 10.540000 11.365000 10.860000 11.685000 ;
      RECT 10.940000  0.005000 11.260000  0.325000 ;
      RECT 10.940000 11.365000 11.260000 11.685000 ;
      RECT 11.340000  0.005000 11.660000  0.325000 ;
      RECT 11.340000 11.365000 11.660000 11.685000 ;
      RECT 11.740000  0.005000 12.060000  0.325000 ;
      RECT 11.740000 11.365000 12.060000 11.685000 ;
      RECT 12.140000  0.005000 12.460000  0.325000 ;
      RECT 12.140000 11.365000 12.460000 11.685000 ;
      RECT 12.540000  0.005000 12.860000  0.325000 ;
      RECT 12.540000 11.365000 12.860000 11.685000 ;
      RECT 12.940000  0.005000 13.260000  0.325000 ;
      RECT 12.940000 11.365000 13.260000 11.685000 ;
      RECT 13.340000  0.005000 13.660000  0.325000 ;
      RECT 13.340000 11.365000 13.660000 11.685000 ;
      RECT 13.740000  0.005000 14.060000  0.325000 ;
      RECT 13.740000 11.365000 14.060000 11.685000 ;
      RECT 14.140000  0.005000 14.460000  0.325000 ;
      RECT 14.140000 11.365000 14.460000 11.685000 ;
      RECT 14.540000  0.005000 14.860000  0.325000 ;
      RECT 14.540000 11.365000 14.860000 11.685000 ;
      RECT 14.940000  0.005000 15.260000  0.325000 ;
      RECT 14.940000 11.365000 15.260000 11.685000 ;
      RECT 15.340000  0.005000 15.660000  0.325000 ;
      RECT 15.340000 11.365000 15.660000 11.685000 ;
      RECT 15.740000  0.005000 16.060000  0.325000 ;
      RECT 15.740000 11.365000 16.060000 11.685000 ;
      RECT 16.140000  0.005000 16.460000  0.325000 ;
      RECT 16.140000 11.365000 16.460000 11.685000 ;
      RECT 16.540000  0.005000 16.860000  0.325000 ;
      RECT 16.540000 11.365000 16.860000 11.685000 ;
      RECT 16.940000  0.005000 17.260000  0.325000 ;
      RECT 16.940000 11.365000 17.260000 11.685000 ;
      RECT 17.340000  0.005000 17.660000  0.325000 ;
      RECT 17.340000 11.365000 17.660000 11.685000 ;
      RECT 17.740000  0.005000 18.060000  0.325000 ;
      RECT 17.740000 11.365000 18.060000 11.685000 ;
      RECT 18.140000  0.005000 18.460000  0.325000 ;
      RECT 18.140000 11.365000 18.460000 11.685000 ;
      RECT 18.540000  0.005000 18.860000  0.325000 ;
      RECT 18.540000 11.365000 18.860000 11.685000 ;
      RECT 18.940000  0.005000 19.260000  0.325000 ;
      RECT 18.940000 11.365000 19.260000 11.685000 ;
      RECT 19.340000  0.005000 19.660000  0.325000 ;
      RECT 19.340000 11.365000 19.660000 11.685000 ;
      RECT 19.740000  0.005000 20.060000  0.325000 ;
      RECT 19.740000 11.365000 20.060000 11.685000 ;
      RECT 20.140000  0.005000 20.460000  0.325000 ;
      RECT 20.140000 11.365000 20.460000 11.685000 ;
      RECT 20.540000  0.005000 20.860000  0.325000 ;
      RECT 20.540000 11.365000 20.860000 11.685000 ;
      RECT 20.940000  0.005000 21.260000  0.325000 ;
      RECT 20.940000 11.365000 21.260000 11.685000 ;
      RECT 21.340000  0.005000 21.660000  0.325000 ;
      RECT 21.340000 11.365000 21.660000 11.685000 ;
      RECT 21.740000  0.005000 22.060000  0.325000 ;
      RECT 21.740000 11.365000 22.060000 11.685000 ;
      RECT 22.140000  0.005000 22.460000  0.325000 ;
      RECT 22.140000 11.365000 22.460000 11.685000 ;
      RECT 22.540000  0.005000 22.860000  0.325000 ;
      RECT 22.540000 11.365000 22.860000 11.685000 ;
      RECT 22.940000  0.005000 23.260000  0.325000 ;
      RECT 22.940000 11.365000 23.260000 11.685000 ;
      RECT 23.340000  0.005000 23.660000  0.325000 ;
      RECT 23.340000 11.365000 23.660000 11.685000 ;
      RECT 23.740000  0.005000 24.060000  0.325000 ;
      RECT 23.740000 11.365000 24.060000 11.685000 ;
      RECT 24.140000  0.005000 24.460000  0.325000 ;
      RECT 24.140000 11.365000 24.460000 11.685000 ;
      RECT 24.540000  0.005000 24.860000  0.325000 ;
      RECT 24.540000 11.365000 24.860000 11.685000 ;
      RECT 24.940000  0.005000 25.260000  0.325000 ;
      RECT 24.940000 11.365000 25.260000 11.685000 ;
      RECT 25.340000  0.005000 25.660000  0.325000 ;
      RECT 25.340000 11.365000 25.660000 11.685000 ;
      RECT 25.740000  0.005000 26.060000  0.325000 ;
      RECT 25.740000 11.365000 26.060000 11.685000 ;
      RECT 26.140000  0.005000 26.460000  0.325000 ;
      RECT 26.140000 11.365000 26.460000 11.685000 ;
      RECT 26.540000  0.005000 26.860000  0.325000 ;
      RECT 26.540000 11.365000 26.860000 11.685000 ;
      RECT 26.940000  0.005000 27.260000  0.325000 ;
      RECT 26.940000 11.365000 27.260000 11.685000 ;
      RECT 27.340000  0.005000 27.660000  0.325000 ;
      RECT 27.340000 11.365000 27.660000 11.685000 ;
      RECT 27.740000  0.005000 28.060000  0.325000 ;
      RECT 27.740000 11.365000 28.060000 11.685000 ;
      RECT 28.140000  0.005000 28.460000  0.325000 ;
      RECT 28.140000 11.365000 28.460000 11.685000 ;
      RECT 28.540000  0.005000 28.860000  0.325000 ;
      RECT 28.540000 11.365000 28.860000 11.685000 ;
      RECT 28.940000  0.005000 29.260000  0.325000 ;
      RECT 28.940000 11.365000 29.260000 11.685000 ;
      RECT 29.340000  0.005000 29.660000  0.325000 ;
      RECT 29.340000 11.365000 29.660000 11.685000 ;
      RECT 29.740000  0.005000 30.060000  0.325000 ;
      RECT 29.740000 11.365000 30.060000 11.685000 ;
      RECT 30.140000  0.005000 30.460000  0.325000 ;
      RECT 30.140000 11.365000 30.460000 11.685000 ;
      RECT 30.540000  0.005000 30.860000  0.325000 ;
      RECT 30.540000 11.365000 30.860000 11.685000 ;
      RECT 30.940000  0.005000 31.260000  0.325000 ;
      RECT 30.940000 11.365000 31.260000 11.685000 ;
      RECT 31.340000  0.005000 31.660000  0.325000 ;
      RECT 31.340000 11.365000 31.660000 11.685000 ;
      RECT 31.740000  0.005000 32.060000  0.325000 ;
      RECT 31.740000 11.365000 32.060000 11.685000 ;
      RECT 32.140000  0.005000 32.460000  0.325000 ;
      RECT 32.140000 11.365000 32.460000 11.685000 ;
      RECT 32.540000  0.005000 32.860000  0.325000 ;
      RECT 32.540000 11.365000 32.860000 11.685000 ;
      RECT 32.940000  0.005000 33.260000  0.325000 ;
      RECT 32.940000 11.365000 33.260000 11.685000 ;
      RECT 33.340000  0.005000 33.660000  0.325000 ;
      RECT 33.340000 11.365000 33.660000 11.685000 ;
      RECT 33.740000  0.005000 34.060000  0.325000 ;
      RECT 33.740000 11.365000 34.060000 11.685000 ;
      RECT 34.140000  0.005000 34.460000  0.325000 ;
      RECT 34.140000 11.365000 34.460000 11.685000 ;
      RECT 34.540000  0.005000 34.860000  0.325000 ;
      RECT 34.540000 11.365000 34.860000 11.685000 ;
      RECT 34.940000  0.005000 35.260000  0.325000 ;
      RECT 34.940000 11.365000 35.260000 11.685000 ;
      RECT 35.340000  0.005000 35.660000  0.325000 ;
      RECT 35.340000 11.365000 35.660000 11.685000 ;
      RECT 35.740000  0.005000 36.060000  0.325000 ;
      RECT 35.740000 11.365000 36.060000 11.685000 ;
      RECT 36.140000  0.005000 36.460000  0.325000 ;
      RECT 36.140000 11.365000 36.460000 11.685000 ;
      RECT 36.540000  0.005000 36.860000  0.325000 ;
      RECT 36.540000 11.365000 36.860000 11.685000 ;
      RECT 36.940000  0.005000 37.260000  0.325000 ;
      RECT 36.940000 11.365000 37.260000 11.685000 ;
      RECT 37.340000  0.005000 37.660000  0.325000 ;
      RECT 37.340000 11.365000 37.660000 11.685000 ;
      RECT 37.740000  0.005000 38.060000  0.325000 ;
      RECT 37.740000 11.365000 38.060000 11.685000 ;
      RECT 38.140000  0.005000 38.460000  0.325000 ;
      RECT 38.140000 11.365000 38.460000 11.685000 ;
      RECT 38.540000  0.005000 38.860000  0.325000 ;
      RECT 38.540000 11.365000 38.860000 11.685000 ;
      RECT 38.940000  0.005000 39.260000  0.325000 ;
      RECT 38.940000 11.365000 39.260000 11.685000 ;
      RECT 39.340000  0.005000 39.660000  0.325000 ;
      RECT 39.340000 11.365000 39.660000 11.685000 ;
      RECT 39.740000  0.005000 40.060000  0.325000 ;
      RECT 39.740000 11.365000 40.060000 11.685000 ;
      RECT 40.140000  0.005000 40.460000  0.325000 ;
      RECT 40.140000 11.365000 40.460000 11.685000 ;
      RECT 40.540000  0.005000 40.860000  0.325000 ;
      RECT 40.540000 11.365000 40.860000 11.685000 ;
      RECT 40.940000  0.005000 41.260000  0.325000 ;
      RECT 40.940000 11.365000 41.260000 11.685000 ;
      RECT 41.340000  0.005000 41.660000  0.325000 ;
      RECT 41.340000 11.365000 41.660000 11.685000 ;
      RECT 41.740000  0.005000 42.060000  0.325000 ;
      RECT 41.740000 11.365000 42.060000 11.685000 ;
      RECT 42.140000  0.005000 42.460000  0.325000 ;
      RECT 42.140000 11.365000 42.460000 11.685000 ;
      RECT 42.540000  0.005000 42.860000  0.325000 ;
      RECT 42.540000 11.365000 42.860000 11.685000 ;
      RECT 42.940000  0.005000 43.260000  0.325000 ;
      RECT 42.940000 11.365000 43.260000 11.685000 ;
      RECT 43.340000  0.005000 43.660000  0.325000 ;
      RECT 43.340000 11.365000 43.660000 11.685000 ;
      RECT 43.740000  0.005000 44.060000  0.325000 ;
      RECT 43.740000 11.365000 44.060000 11.685000 ;
      RECT 44.140000  0.005000 44.460000  0.325000 ;
      RECT 44.140000 11.365000 44.460000 11.685000 ;
      RECT 44.540000  0.005000 44.860000  0.325000 ;
      RECT 44.540000 11.365000 44.860000 11.685000 ;
      RECT 44.940000  0.005000 45.260000  0.325000 ;
      RECT 44.940000 11.365000 45.260000 11.685000 ;
      RECT 45.340000  0.005000 45.660000  0.325000 ;
      RECT 45.340000 11.365000 45.660000 11.685000 ;
      RECT 45.740000  0.005000 46.060000  0.325000 ;
      RECT 45.740000 11.365000 46.060000 11.685000 ;
      RECT 46.140000  0.005000 46.460000  0.325000 ;
      RECT 46.140000 11.365000 46.460000 11.685000 ;
      RECT 46.540000  0.005000 46.860000  0.325000 ;
      RECT 46.540000 11.365000 46.860000 11.685000 ;
      RECT 46.940000  0.005000 47.260000  0.325000 ;
      RECT 46.940000 11.365000 47.260000 11.685000 ;
      RECT 47.340000  0.005000 47.660000  0.325000 ;
      RECT 47.340000 11.365000 47.660000 11.685000 ;
      RECT 47.740000  0.005000 48.060000  0.325000 ;
      RECT 47.740000 11.365000 48.060000 11.685000 ;
      RECT 48.140000  0.005000 48.460000  0.325000 ;
      RECT 48.140000 11.365000 48.460000 11.685000 ;
      RECT 48.540000  0.005000 48.860000  0.325000 ;
      RECT 48.540000 11.365000 48.860000 11.685000 ;
      RECT 48.940000  0.005000 49.260000  0.325000 ;
      RECT 48.940000 11.365000 49.260000 11.685000 ;
      RECT 49.340000  0.005000 49.660000  0.325000 ;
      RECT 49.340000 11.365000 49.660000 11.685000 ;
      RECT 49.740000  0.005000 50.060000  0.325000 ;
      RECT 49.740000 11.365000 50.060000 11.685000 ;
      RECT 50.140000  0.005000 50.460000  0.325000 ;
      RECT 50.140000 11.365000 50.460000 11.685000 ;
      RECT 50.540000  0.005000 50.860000  0.325000 ;
      RECT 50.540000 11.365000 50.860000 11.685000 ;
      RECT 50.940000  0.005000 51.260000  0.325000 ;
      RECT 50.940000 11.365000 51.260000 11.685000 ;
      RECT 51.340000  0.005000 51.660000  0.325000 ;
      RECT 51.340000 11.365000 51.660000 11.685000 ;
      RECT 51.740000  0.005000 52.060000  0.325000 ;
      RECT 51.740000 11.365000 52.060000 11.685000 ;
      RECT 52.140000  0.005000 52.460000  0.325000 ;
      RECT 52.140000 11.365000 52.460000 11.685000 ;
      RECT 52.540000  0.005000 52.860000  0.325000 ;
      RECT 52.540000 11.365000 52.860000 11.685000 ;
      RECT 52.940000  0.005000 53.260000  0.325000 ;
      RECT 52.940000 11.365000 53.260000 11.685000 ;
      RECT 53.340000  0.005000 53.660000  0.325000 ;
      RECT 53.340000 11.365000 53.660000 11.685000 ;
      RECT 53.740000  0.005000 54.060000  0.325000 ;
      RECT 53.740000 11.365000 54.060000 11.685000 ;
      RECT 54.140000  0.005000 54.460000  0.325000 ;
      RECT 54.140000 11.365000 54.460000 11.685000 ;
      RECT 54.540000  0.005000 54.860000  0.325000 ;
      RECT 54.540000 11.365000 54.860000 11.685000 ;
      RECT 54.940000  0.005000 55.260000  0.325000 ;
      RECT 54.940000 11.365000 55.260000 11.685000 ;
    LAYER via4 ;
      RECT  0.760000 9.990000  1.940000 11.170000 ;
      RECT  1.360000 0.520000  2.540000  1.700000 ;
      RECT  7.960000 9.990000  9.140000 11.170000 ;
      RECT  8.560000 0.520000  9.740000  1.700000 ;
      RECT 15.160000 9.990000 16.340000 11.170000 ;
      RECT 15.760000 0.520000 16.940000  1.700000 ;
      RECT 22.360000 9.990000 23.540000 11.170000 ;
      RECT 22.960000 0.520000 24.140000  1.700000 ;
      RECT 29.560000 9.990000 30.740000 11.170000 ;
      RECT 30.160000 0.520000 31.340000  1.700000 ;
      RECT 36.760000 9.990000 37.940000 11.170000 ;
      RECT 37.360000 0.520000 38.540000  1.700000 ;
      RECT 43.960000 9.990000 45.140000 11.170000 ;
      RECT 44.560000 0.520000 45.740000  1.700000 ;
      RECT 51.160000 9.990000 52.340000 11.170000 ;
      RECT 51.760000 0.520000 52.940000  1.700000 ;
  END
END sky130_fd_pr__cap_vpp_55p8x11p7_pol1m1m2m3m4m5_noshield_m5pullin
END LIBRARY
