* SKY130 Spice File.
.include "../../sonos_e/begin_of_life.pm3.spice"
.include "../../sonos_p/begin_of_life.pm3.spice"
.include "../../sonos_e/begin_of_life/typical.spice"
.include "../../sonos_p/begin_of_life/typical.spice"
