# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.880000 BY  4.030000 ;
  PIN BULK
    ANTENNADIFFAREA  1.745800 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.610000 0.470000 3.420000 ;
        RECT 3.410000 0.610000 3.700000 3.420000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.140000 3.830000 3.420000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.010000 ;
    PORT
      LAYER li1 ;
        RECT 0.925000 0.100000 2.955000 0.270000 ;
        RECT 0.925000 3.760000 2.955000 3.930000 ;
      LAYER mcon ;
        RECT 0.960000 0.100000 1.130000 0.270000 ;
        RECT 0.960000 3.760000 1.130000 3.930000 ;
        RECT 1.320000 0.100000 1.490000 0.270000 ;
        RECT 1.320000 3.760000 1.490000 3.930000 ;
        RECT 1.680000 0.100000 1.850000 0.270000 ;
        RECT 1.680000 3.760000 1.850000 3.930000 ;
        RECT 2.040000 0.100000 2.210000 0.270000 ;
        RECT 2.040000 3.760000 2.210000 3.930000 ;
        RECT 2.400000 0.100000 2.570000 0.270000 ;
        RECT 2.400000 3.760000 2.570000 3.930000 ;
        RECT 2.760000 0.100000 2.930000 0.270000 ;
        RECT 2.760000 3.760000 2.930000 3.930000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.900000 0.000000 2.990000 0.330000 ;
        RECT 0.900000 3.700000 2.990000 4.030000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.528400 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.610000 3.830000 1.890000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.660000 0.410000 3.370000 ;
      RECT 0.795000 0.490000 0.965000 3.540000 ;
      RECT 1.325000 0.490000 1.495000 3.540000 ;
      RECT 1.855000 0.490000 2.025000 3.540000 ;
      RECT 2.385000 0.490000 2.555000 3.540000 ;
      RECT 2.915000 0.490000 3.085000 3.540000 ;
      RECT 3.470000 0.660000 3.640000 3.370000 ;
    LAYER mcon ;
      RECT 0.240000 0.670000 0.410000 0.840000 ;
      RECT 0.240000 1.030000 0.410000 1.200000 ;
      RECT 0.240000 1.390000 0.410000 1.560000 ;
      RECT 0.240000 1.750000 0.410000 1.920000 ;
      RECT 0.240000 2.110000 0.410000 2.280000 ;
      RECT 0.240000 2.470000 0.410000 2.640000 ;
      RECT 0.240000 2.830000 0.410000 3.000000 ;
      RECT 0.240000 3.190000 0.410000 3.360000 ;
      RECT 0.795000 0.670000 0.965000 0.840000 ;
      RECT 0.795000 1.030000 0.965000 1.200000 ;
      RECT 0.795000 1.390000 0.965000 1.560000 ;
      RECT 0.795000 1.750000 0.965000 1.920000 ;
      RECT 0.795000 2.110000 0.965000 2.280000 ;
      RECT 0.795000 2.470000 0.965000 2.640000 ;
      RECT 0.795000 2.830000 0.965000 3.000000 ;
      RECT 0.795000 3.190000 0.965000 3.360000 ;
      RECT 1.325000 0.670000 1.495000 0.840000 ;
      RECT 1.325000 1.030000 1.495000 1.200000 ;
      RECT 1.325000 1.390000 1.495000 1.560000 ;
      RECT 1.325000 1.750000 1.495000 1.920000 ;
      RECT 1.325000 2.110000 1.495000 2.280000 ;
      RECT 1.325000 2.470000 1.495000 2.640000 ;
      RECT 1.325000 2.830000 1.495000 3.000000 ;
      RECT 1.325000 3.190000 1.495000 3.360000 ;
      RECT 1.855000 0.670000 2.025000 0.840000 ;
      RECT 1.855000 1.030000 2.025000 1.200000 ;
      RECT 1.855000 1.390000 2.025000 1.560000 ;
      RECT 1.855000 1.750000 2.025000 1.920000 ;
      RECT 1.855000 2.110000 2.025000 2.280000 ;
      RECT 1.855000 2.470000 2.025000 2.640000 ;
      RECT 1.855000 2.830000 2.025000 3.000000 ;
      RECT 1.855000 3.190000 2.025000 3.360000 ;
      RECT 2.385000 0.670000 2.555000 0.840000 ;
      RECT 2.385000 1.030000 2.555000 1.200000 ;
      RECT 2.385000 1.390000 2.555000 1.560000 ;
      RECT 2.385000 1.750000 2.555000 1.920000 ;
      RECT 2.385000 2.110000 2.555000 2.280000 ;
      RECT 2.385000 2.470000 2.555000 2.640000 ;
      RECT 2.385000 2.830000 2.555000 3.000000 ;
      RECT 2.385000 3.190000 2.555000 3.360000 ;
      RECT 2.915000 0.670000 3.085000 0.840000 ;
      RECT 2.915000 1.030000 3.085000 1.200000 ;
      RECT 2.915000 1.390000 3.085000 1.560000 ;
      RECT 2.915000 1.750000 3.085000 1.920000 ;
      RECT 2.915000 2.110000 3.085000 2.280000 ;
      RECT 2.915000 2.470000 3.085000 2.640000 ;
      RECT 2.915000 2.830000 3.085000 3.000000 ;
      RECT 2.915000 3.190000 3.085000 3.360000 ;
      RECT 3.470000 0.670000 3.640000 0.840000 ;
      RECT 3.470000 1.030000 3.640000 1.200000 ;
      RECT 3.470000 1.390000 3.640000 1.560000 ;
      RECT 3.470000 1.750000 3.640000 1.920000 ;
      RECT 3.470000 2.110000 3.640000 2.280000 ;
      RECT 3.470000 2.470000 3.640000 2.640000 ;
      RECT 3.470000 2.830000 3.640000 3.000000 ;
      RECT 3.470000 3.190000 3.640000 3.360000 ;
    LAYER met1 ;
      RECT 0.750000 0.610000 1.010000 3.420000 ;
      RECT 1.280000 0.610000 1.540000 3.420000 ;
      RECT 1.810000 0.610000 2.070000 3.420000 ;
      RECT 2.340000 0.610000 2.600000 3.420000 ;
      RECT 2.870000 0.610000 3.130000 3.420000 ;
    LAYER via ;
      RECT 0.750000 0.640000 1.010000 0.900000 ;
      RECT 0.750000 0.960000 1.010000 1.220000 ;
      RECT 0.750000 1.280000 1.010000 1.540000 ;
      RECT 0.750000 1.600000 1.010000 1.860000 ;
      RECT 1.280000 2.170000 1.540000 2.430000 ;
      RECT 1.280000 2.490000 1.540000 2.750000 ;
      RECT 1.280000 2.810000 1.540000 3.070000 ;
      RECT 1.280000 3.130000 1.540000 3.390000 ;
      RECT 1.810000 0.640000 2.070000 0.900000 ;
      RECT 1.810000 0.960000 2.070000 1.220000 ;
      RECT 1.810000 1.280000 2.070000 1.540000 ;
      RECT 1.810000 1.600000 2.070000 1.860000 ;
      RECT 2.340000 2.170000 2.600000 2.430000 ;
      RECT 2.340000 2.490000 2.600000 2.750000 ;
      RECT 2.340000 2.810000 2.600000 3.070000 ;
      RECT 2.340000 3.130000 2.600000 3.390000 ;
      RECT 2.870000 0.640000 3.130000 0.900000 ;
      RECT 2.870000 0.960000 3.130000 1.220000 ;
      RECT 2.870000 1.280000 3.130000 1.540000 ;
      RECT 2.870000 1.600000 3.130000 1.860000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25
END LIBRARY
