magic
tech sky130A
magscale 1 2
timestamp 1762019803
<< pwell >>
rect -276 -813 276 813
<< nmos >>
rect -80 403 80 603
rect -80 47 80 247
rect -80 -309 80 -109
rect -80 -665 80 -465
<< ndiff >>
rect -138 591 -80 603
rect -138 415 -126 591
rect -92 415 -80 591
rect -138 403 -80 415
rect 80 591 138 603
rect 80 415 92 591
rect 126 415 138 591
rect 80 403 138 415
rect -138 235 -80 247
rect -138 59 -126 235
rect -92 59 -80 235
rect -138 47 -80 59
rect 80 235 138 247
rect 80 59 92 235
rect 126 59 138 235
rect 80 47 138 59
rect -138 -121 -80 -109
rect -138 -297 -126 -121
rect -92 -297 -80 -121
rect -138 -309 -80 -297
rect 80 -121 138 -109
rect 80 -297 92 -121
rect 126 -297 138 -121
rect 80 -309 138 -297
rect -138 -477 -80 -465
rect -138 -653 -126 -477
rect -92 -653 -80 -477
rect -138 -665 -80 -653
rect 80 -477 138 -465
rect 80 -653 92 -477
rect 126 -653 138 -477
rect 80 -665 138 -653
<< ndiffc >>
rect -126 415 -92 591
rect 92 415 126 591
rect -126 59 -92 235
rect 92 59 126 235
rect -126 -297 -92 -121
rect 92 -297 126 -121
rect -126 -653 -92 -477
rect 92 -653 126 -477
<< psubdiff >>
rect -240 743 -144 777
rect 144 743 240 777
rect -240 681 -206 743
rect 206 681 240 743
rect -240 -743 -206 -681
rect 206 -743 240 -681
rect -240 -777 -144 -743
rect 144 -777 240 -743
<< psubdiffcont >>
rect -144 743 144 777
rect -240 -681 -206 681
rect 206 -681 240 681
rect -144 -777 144 -743
<< poly >>
rect -80 675 80 691
rect -80 641 -64 675
rect 64 641 80 675
rect -80 603 80 641
rect -80 377 80 403
rect -80 319 80 335
rect -80 285 -64 319
rect 64 285 80 319
rect -80 247 80 285
rect -80 21 80 47
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -109 80 -71
rect -80 -335 80 -309
rect -80 -393 80 -377
rect -80 -427 -64 -393
rect 64 -427 80 -393
rect -80 -465 80 -427
rect -80 -691 80 -665
<< polycont >>
rect -64 641 64 675
rect -64 285 64 319
rect -64 -71 64 -37
rect -64 -427 64 -393
<< locali >>
rect -240 743 -144 777
rect 144 743 240 777
rect -240 681 -206 743
rect 206 681 240 743
rect -80 641 -64 675
rect 64 641 80 675
rect -126 591 -92 607
rect -126 399 -92 415
rect 92 591 126 607
rect 92 399 126 415
rect -80 285 -64 319
rect 64 285 80 319
rect -126 235 -92 251
rect -126 43 -92 59
rect 92 235 126 251
rect 92 43 126 59
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -121 -92 -105
rect -126 -313 -92 -297
rect 92 -121 126 -105
rect 92 -313 126 -297
rect -80 -427 -64 -393
rect 64 -427 80 -393
rect -126 -477 -92 -461
rect -126 -669 -92 -653
rect 92 -477 126 -461
rect 92 -669 126 -653
rect -240 -743 -206 -681
rect 206 -743 240 -681
rect -240 -777 -144 -743
rect 144 -777 240 -743
<< viali >>
rect -64 641 64 675
rect -126 415 -92 591
rect 92 415 126 591
rect -64 285 64 319
rect -126 59 -92 235
rect 92 59 126 235
rect -64 -71 64 -37
rect -126 -297 -92 -121
rect 92 -297 126 -121
rect -64 -427 64 -393
rect -126 -653 -92 -477
rect 92 -653 126 -477
<< metal1 >>
rect -76 675 76 681
rect -76 641 -64 675
rect 64 641 76 675
rect -76 635 76 641
rect -132 591 -86 603
rect -132 415 -126 591
rect -92 415 -86 591
rect -132 403 -86 415
rect 86 591 132 603
rect 86 415 92 591
rect 126 415 132 591
rect 86 403 132 415
rect -76 319 76 325
rect -76 285 -64 319
rect 64 285 76 319
rect -76 279 76 285
rect -132 235 -86 247
rect -132 59 -126 235
rect -92 59 -86 235
rect -132 47 -86 59
rect 86 235 132 247
rect 86 59 92 235
rect 126 59 132 235
rect 86 47 132 59
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -121 -86 -109
rect -132 -297 -126 -121
rect -92 -297 -86 -121
rect -132 -309 -86 -297
rect 86 -121 132 -109
rect 86 -297 92 -121
rect 126 -297 132 -121
rect 86 -309 132 -297
rect -76 -393 76 -387
rect -76 -427 -64 -393
rect 64 -427 76 -393
rect -76 -433 76 -427
rect -132 -477 -86 -465
rect -132 -653 -126 -477
rect -92 -653 -86 -477
rect -132 -665 -86 -653
rect 86 -477 132 -465
rect 86 -653 92 -477
rect 126 -653 132 -477
rect 86 -665 132 -653
<< labels >>
rlabel psubdiffcont 0 -760 0 -760 0 B
port 1 nsew
rlabel ndiffc -109 -565 -109 -565 0 D0
port 2 nsew
rlabel ndiffc 109 -565 109 -565 0 S0
port 3 nsew
rlabel polycont 0 -410 0 -410 0 G0
port 4 nsew
rlabel ndiffc -109 -209 -109 -209 0 D1
port 5 nsew
rlabel ndiffc 109 -209 109 -209 0 S1
port 6 nsew
rlabel polycont 0 -54 0 -54 0 G1
port 7 nsew
rlabel ndiffc -109 147 -109 147 0 D2
port 8 nsew
rlabel ndiffc 109 147 109 147 0 S2
port 9 nsew
rlabel polycont 0 302 0 302 0 G2
port 10 nsew
rlabel ndiffc -109 503 -109 503 0 D3
port 11 nsew
rlabel ndiffc 109 503 109 503 0 S3
port 12 nsew
rlabel polycont 0 658 0 658 0 G3
port 13 nsew
<< properties >>
string FIXED_BBOX -223 -760 223 760
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.8 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
