# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.280000 BY  4.030000 ;
  PIN BULK
    ANTENNADIFFAREA  1.745800 ;
    PORT
      LAYER li1 ;
        RECT 0.240000 0.660000 0.410000 3.370000 ;
        RECT 3.870000 0.660000 4.040000 3.370000 ;
      LAYER mcon ;
        RECT 0.240000 0.670000 0.410000 0.840000 ;
        RECT 0.240000 1.030000 0.410000 1.200000 ;
        RECT 0.240000 1.390000 0.410000 1.560000 ;
        RECT 0.240000 1.750000 0.410000 1.920000 ;
        RECT 0.240000 2.110000 0.410000 2.280000 ;
        RECT 0.240000 2.470000 0.410000 2.640000 ;
        RECT 0.240000 2.830000 0.410000 3.000000 ;
        RECT 0.240000 3.190000 0.410000 3.360000 ;
        RECT 3.870000 0.670000 4.040000 0.840000 ;
        RECT 3.870000 1.030000 4.040000 1.200000 ;
        RECT 3.870000 1.390000 4.040000 1.560000 ;
        RECT 3.870000 1.750000 4.040000 1.920000 ;
        RECT 3.870000 2.110000 4.040000 2.280000 ;
        RECT 3.870000 2.470000 4.040000 2.640000 ;
        RECT 3.870000 2.830000 4.040000 3.000000 ;
        RECT 3.870000 3.190000 4.040000 3.360000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.180000 0.610000 0.470000 3.420000 ;
        RECT 3.810000 0.610000 4.100000 3.420000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.140000 4.230000 3.420000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  4.214000 ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.100000 3.325000 0.270000 ;
        RECT 0.955000 3.760000 3.325000 3.930000 ;
      LAYER mcon ;
        RECT 0.975000 0.100000 1.145000 0.270000 ;
        RECT 0.975000 3.760000 1.145000 3.930000 ;
        RECT 1.335000 0.100000 1.505000 0.270000 ;
        RECT 1.335000 3.760000 1.505000 3.930000 ;
        RECT 1.695000 0.100000 1.865000 0.270000 ;
        RECT 1.695000 3.760000 1.865000 3.930000 ;
        RECT 2.055000 0.100000 2.225000 0.270000 ;
        RECT 2.055000 3.760000 2.225000 3.930000 ;
        RECT 2.415000 0.100000 2.585000 0.270000 ;
        RECT 2.415000 3.760000 2.585000 3.930000 ;
        RECT 2.775000 0.100000 2.945000 0.270000 ;
        RECT 2.775000 3.760000 2.945000 3.930000 ;
        RECT 3.135000 0.100000 3.305000 0.270000 ;
        RECT 3.135000 3.760000 3.305000 3.930000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.915000 0.000000 3.365000 0.330000 ;
        RECT 0.915000 3.700000 3.365000 4.030000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.528400 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.610000 4.230000 1.890000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.795000 0.490000 0.965000 3.540000 ;
      RECT 1.425000 0.490000 1.595000 3.540000 ;
      RECT 2.055000 0.490000 2.225000 3.540000 ;
      RECT 2.685000 0.490000 2.855000 3.540000 ;
      RECT 3.315000 0.490000 3.485000 3.540000 ;
    LAYER mcon ;
      RECT 0.795000 0.670000 0.965000 0.840000 ;
      RECT 0.795000 1.030000 0.965000 1.200000 ;
      RECT 0.795000 1.390000 0.965000 1.560000 ;
      RECT 0.795000 1.750000 0.965000 1.920000 ;
      RECT 0.795000 2.110000 0.965000 2.280000 ;
      RECT 0.795000 2.470000 0.965000 2.640000 ;
      RECT 0.795000 2.830000 0.965000 3.000000 ;
      RECT 0.795000 3.190000 0.965000 3.360000 ;
      RECT 1.425000 0.670000 1.595000 0.840000 ;
      RECT 1.425000 1.030000 1.595000 1.200000 ;
      RECT 1.425000 1.390000 1.595000 1.560000 ;
      RECT 1.425000 1.750000 1.595000 1.920000 ;
      RECT 1.425000 2.110000 1.595000 2.280000 ;
      RECT 1.425000 2.470000 1.595000 2.640000 ;
      RECT 1.425000 2.830000 1.595000 3.000000 ;
      RECT 1.425000 3.190000 1.595000 3.360000 ;
      RECT 2.055000 0.670000 2.225000 0.840000 ;
      RECT 2.055000 1.030000 2.225000 1.200000 ;
      RECT 2.055000 1.390000 2.225000 1.560000 ;
      RECT 2.055000 1.750000 2.225000 1.920000 ;
      RECT 2.055000 2.110000 2.225000 2.280000 ;
      RECT 2.055000 2.470000 2.225000 2.640000 ;
      RECT 2.055000 2.830000 2.225000 3.000000 ;
      RECT 2.055000 3.190000 2.225000 3.360000 ;
      RECT 2.685000 0.670000 2.855000 0.840000 ;
      RECT 2.685000 1.030000 2.855000 1.200000 ;
      RECT 2.685000 1.390000 2.855000 1.560000 ;
      RECT 2.685000 1.750000 2.855000 1.920000 ;
      RECT 2.685000 2.110000 2.855000 2.280000 ;
      RECT 2.685000 2.470000 2.855000 2.640000 ;
      RECT 2.685000 2.830000 2.855000 3.000000 ;
      RECT 2.685000 3.190000 2.855000 3.360000 ;
      RECT 3.315000 0.670000 3.485000 0.840000 ;
      RECT 3.315000 1.030000 3.485000 1.200000 ;
      RECT 3.315000 1.390000 3.485000 1.560000 ;
      RECT 3.315000 1.750000 3.485000 1.920000 ;
      RECT 3.315000 2.110000 3.485000 2.280000 ;
      RECT 3.315000 2.470000 3.485000 2.640000 ;
      RECT 3.315000 2.830000 3.485000 3.000000 ;
      RECT 3.315000 3.190000 3.485000 3.360000 ;
    LAYER met1 ;
      RECT 0.750000 0.610000 1.010000 3.420000 ;
      RECT 1.380000 0.610000 1.640000 3.420000 ;
      RECT 2.010000 0.610000 2.270000 3.420000 ;
      RECT 2.640000 0.610000 2.900000 3.420000 ;
      RECT 3.270000 0.610000 3.530000 3.420000 ;
    LAYER via ;
      RECT 0.750000 0.640000 1.010000 0.900000 ;
      RECT 0.750000 0.960000 1.010000 1.220000 ;
      RECT 0.750000 1.280000 1.010000 1.540000 ;
      RECT 0.750000 1.600000 1.010000 1.860000 ;
      RECT 1.380000 2.170000 1.640000 2.430000 ;
      RECT 1.380000 2.490000 1.640000 2.750000 ;
      RECT 1.380000 2.810000 1.640000 3.070000 ;
      RECT 1.380000 3.130000 1.640000 3.390000 ;
      RECT 2.010000 0.640000 2.270000 0.900000 ;
      RECT 2.010000 0.960000 2.270000 1.220000 ;
      RECT 2.010000 1.280000 2.270000 1.540000 ;
      RECT 2.010000 1.600000 2.270000 1.860000 ;
      RECT 2.640000 2.170000 2.900000 2.430000 ;
      RECT 2.640000 2.490000 2.900000 2.750000 ;
      RECT 2.640000 2.810000 2.900000 3.070000 ;
      RECT 2.640000 3.130000 2.900000 3.390000 ;
      RECT 3.270000 0.640000 3.530000 0.900000 ;
      RECT 3.270000 0.960000 3.530000 1.220000 ;
      RECT 3.270000 1.280000 3.530000 1.540000 ;
      RECT 3.270000 1.600000 3.530000 1.860000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35
END LIBRARY
