# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_20v0_withptap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_20v0_withptap ;
  ORIGIN  7.900000  9.020000 ;
  SIZE  16.55000 BY  48.04000 ;
  OBS
    LAYER li1 ;
      RECT -7.900000 -9.020000  8.650000 -8.610000 ;
      RECT -7.900000 -8.610000 -7.490000 38.610000 ;
      RECT -7.900000 38.610000  8.650000 39.020000 ;
      RECT -3.990000 -5.110000  4.740000 -3.785000 ;
      RECT -3.990000 -3.785000 -3.580000 33.785000 ;
      RECT -3.990000 33.785000  4.740000 35.110000 ;
      RECT -3.295000 -0.820000 -2.285000 30.825000 ;
      RECT -0.730000 -3.285000  1.450000 -2.215000 ;
      RECT -0.670000 -0.820000  1.420000 30.825000 ;
      RECT  3.035000 -0.820000  4.045000 30.825000 ;
      RECT  4.330000 -3.785000  4.740000 33.785000 ;
      RECT  8.240000 -8.610000  8.650000 38.610000 ;
    LAYER mcon ;
      RECT -7.780000 -8.305000 -7.610000 -8.135000 ;
      RECT -7.780000 -7.945000 -7.610000 -7.775000 ;
      RECT -7.780000 -7.585000 -7.610000 -7.415000 ;
      RECT -7.780000 -7.225000 -7.610000 -7.055000 ;
      RECT -7.780000 -6.865000 -7.610000 -6.695000 ;
      RECT -7.780000 -6.505000 -7.610000 -6.335000 ;
      RECT -7.780000 -6.145000 -7.610000 -5.975000 ;
      RECT -7.780000 -5.785000 -7.610000 -5.615000 ;
      RECT -7.780000 -5.425000 -7.610000 -5.255000 ;
      RECT -7.780000 -5.065000 -7.610000 -4.895000 ;
      RECT -7.780000 -4.705000 -7.610000 -4.535000 ;
      RECT -7.780000 -4.345000 -7.610000 -4.175000 ;
      RECT -7.780000 -3.985000 -7.610000 -3.815000 ;
      RECT -7.780000 -3.625000 -7.610000 -3.455000 ;
      RECT -7.780000 -3.265000 -7.610000 -3.095000 ;
      RECT -7.780000 -2.905000 -7.610000 -2.735000 ;
      RECT -7.780000 -2.545000 -7.610000 -2.375000 ;
      RECT -7.780000 -2.185000 -7.610000 -2.015000 ;
      RECT -7.780000 -1.825000 -7.610000 -1.655000 ;
      RECT -7.780000 -1.465000 -7.610000 -1.295000 ;
      RECT -7.780000 -1.105000 -7.610000 -0.935000 ;
      RECT -7.780000 -0.745000 -7.610000 -0.575000 ;
      RECT -7.780000 -0.385000 -7.610000 -0.215000 ;
      RECT -7.780000 -0.025000 -7.610000  0.145000 ;
      RECT -7.780000  0.335000 -7.610000  0.505000 ;
      RECT -7.780000  0.695000 -7.610000  0.865000 ;
      RECT -7.780000  1.055000 -7.610000  1.225000 ;
      RECT -7.780000  1.415000 -7.610000  1.585000 ;
      RECT -7.780000  1.775000 -7.610000  1.945000 ;
      RECT -7.780000  2.135000 -7.610000  2.305000 ;
      RECT -7.780000  2.495000 -7.610000  2.665000 ;
      RECT -7.780000  2.855000 -7.610000  3.025000 ;
      RECT -7.780000  3.215000 -7.610000  3.385000 ;
      RECT -7.780000  3.575000 -7.610000  3.745000 ;
      RECT -7.780000  3.935000 -7.610000  4.105000 ;
      RECT -7.780000  4.295000 -7.610000  4.465000 ;
      RECT -7.780000  4.655000 -7.610000  4.825000 ;
      RECT -7.780000  5.015000 -7.610000  5.185000 ;
      RECT -7.780000  5.375000 -7.610000  5.545000 ;
      RECT -7.780000  5.735000 -7.610000  5.905000 ;
      RECT -7.780000  6.095000 -7.610000  6.265000 ;
      RECT -7.780000  6.455000 -7.610000  6.625000 ;
      RECT -7.780000  6.815000 -7.610000  6.985000 ;
      RECT -7.780000  7.175000 -7.610000  7.345000 ;
      RECT -7.780000  7.535000 -7.610000  7.705000 ;
      RECT -7.780000  7.895000 -7.610000  8.065000 ;
      RECT -7.780000  8.255000 -7.610000  8.425000 ;
      RECT -7.780000  8.615000 -7.610000  8.785000 ;
      RECT -7.780000  8.975000 -7.610000  9.145000 ;
      RECT -7.780000  9.335000 -7.610000  9.505000 ;
      RECT -7.780000  9.695000 -7.610000  9.865000 ;
      RECT -7.780000 10.055000 -7.610000 10.225000 ;
      RECT -7.780000 10.415000 -7.610000 10.585000 ;
      RECT -7.780000 10.775000 -7.610000 10.945000 ;
      RECT -7.780000 11.135000 -7.610000 11.305000 ;
      RECT -7.780000 11.495000 -7.610000 11.665000 ;
      RECT -7.780000 11.855000 -7.610000 12.025000 ;
      RECT -7.780000 12.215000 -7.610000 12.385000 ;
      RECT -7.780000 12.575000 -7.610000 12.745000 ;
      RECT -7.780000 12.935000 -7.610000 13.105000 ;
      RECT -7.780000 13.295000 -7.610000 13.465000 ;
      RECT -7.780000 13.655000 -7.610000 13.825000 ;
      RECT -7.780000 14.015000 -7.610000 14.185000 ;
      RECT -7.780000 14.375000 -7.610000 14.545000 ;
      RECT -7.780000 14.735000 -7.610000 14.905000 ;
      RECT -7.780000 15.095000 -7.610000 15.265000 ;
      RECT -7.780000 15.455000 -7.610000 15.625000 ;
      RECT -7.780000 15.815000 -7.610000 15.985000 ;
      RECT -7.780000 16.175000 -7.610000 16.345000 ;
      RECT -7.780000 16.535000 -7.610000 16.705000 ;
      RECT -7.780000 16.895000 -7.610000 17.065000 ;
      RECT -7.780000 17.255000 -7.610000 17.425000 ;
      RECT -7.780000 17.615000 -7.610000 17.785000 ;
      RECT -7.780000 17.975000 -7.610000 18.145000 ;
      RECT -7.780000 18.335000 -7.610000 18.505000 ;
      RECT -7.780000 18.695000 -7.610000 18.865000 ;
      RECT -7.780000 19.055000 -7.610000 19.225000 ;
      RECT -7.780000 19.415000 -7.610000 19.585000 ;
      RECT -7.780000 19.775000 -7.610000 19.945000 ;
      RECT -7.780000 20.135000 -7.610000 20.305000 ;
      RECT -7.780000 20.495000 -7.610000 20.665000 ;
      RECT -7.780000 20.855000 -7.610000 21.025000 ;
      RECT -7.780000 21.215000 -7.610000 21.385000 ;
      RECT -7.780000 21.575000 -7.610000 21.745000 ;
      RECT -7.780000 21.935000 -7.610000 22.105000 ;
      RECT -7.780000 22.295000 -7.610000 22.465000 ;
      RECT -7.780000 22.655000 -7.610000 22.825000 ;
      RECT -7.780000 23.015000 -7.610000 23.185000 ;
      RECT -7.780000 23.375000 -7.610000 23.545000 ;
      RECT -7.780000 23.735000 -7.610000 23.905000 ;
      RECT -7.780000 24.095000 -7.610000 24.265000 ;
      RECT -7.780000 24.455000 -7.610000 24.625000 ;
      RECT -7.780000 24.815000 -7.610000 24.985000 ;
      RECT -7.780000 25.175000 -7.610000 25.345000 ;
      RECT -7.780000 25.535000 -7.610000 25.705000 ;
      RECT -7.780000 25.895000 -7.610000 26.065000 ;
      RECT -7.780000 26.255000 -7.610000 26.425000 ;
      RECT -7.780000 26.615000 -7.610000 26.785000 ;
      RECT -7.780000 26.975000 -7.610000 27.145000 ;
      RECT -7.780000 27.335000 -7.610000 27.505000 ;
      RECT -7.780000 27.695000 -7.610000 27.865000 ;
      RECT -7.780000 28.055000 -7.610000 28.225000 ;
      RECT -7.780000 28.415000 -7.610000 28.585000 ;
      RECT -7.780000 28.775000 -7.610000 28.945000 ;
      RECT -7.780000 29.135000 -7.610000 29.305000 ;
      RECT -7.780000 29.495000 -7.610000 29.665000 ;
      RECT -7.780000 29.855000 -7.610000 30.025000 ;
      RECT -7.780000 30.215000 -7.610000 30.385000 ;
      RECT -7.780000 30.575000 -7.610000 30.745000 ;
      RECT -7.780000 30.935000 -7.610000 31.105000 ;
      RECT -7.780000 31.295000 -7.610000 31.465000 ;
      RECT -7.780000 31.655000 -7.610000 31.825000 ;
      RECT -7.780000 32.015000 -7.610000 32.185000 ;
      RECT -7.780000 32.375000 -7.610000 32.545000 ;
      RECT -7.780000 32.735000 -7.610000 32.905000 ;
      RECT -7.780000 33.095000 -7.610000 33.265000 ;
      RECT -7.780000 33.455000 -7.610000 33.625000 ;
      RECT -7.780000 33.815000 -7.610000 33.985000 ;
      RECT -7.780000 34.175000 -7.610000 34.345000 ;
      RECT -7.780000 34.535000 -7.610000 34.705000 ;
      RECT -7.780000 34.895000 -7.610000 35.065000 ;
      RECT -7.780000 35.255000 -7.610000 35.425000 ;
      RECT -7.780000 35.615000 -7.610000 35.785000 ;
      RECT -7.780000 35.975000 -7.610000 36.145000 ;
      RECT -7.780000 36.335000 -7.610000 36.505000 ;
      RECT -7.780000 36.695000 -7.610000 36.865000 ;
      RECT -7.780000 37.055000 -7.610000 37.225000 ;
      RECT -7.780000 37.415000 -7.610000 37.585000 ;
      RECT -7.780000 37.775000 -7.610000 37.945000 ;
      RECT -7.780000 38.135000 -7.610000 38.305000 ;
      RECT -7.270000 -8.900000 -7.100000 -8.730000 ;
      RECT -7.270000 38.730000 -7.100000 38.900000 ;
      RECT -6.910000 -8.900000 -6.740000 -8.730000 ;
      RECT -6.910000 38.730000 -6.740000 38.900000 ;
      RECT -6.550000 -8.900000 -6.380000 -8.730000 ;
      RECT -6.550000 38.730000 -6.380000 38.900000 ;
      RECT -6.190000 -8.900000 -6.020000 -8.730000 ;
      RECT -6.190000 38.730000 -6.020000 38.900000 ;
      RECT -5.830000 -8.900000 -5.660000 -8.730000 ;
      RECT -5.830000 38.730000 -5.660000 38.900000 ;
      RECT -5.470000 -8.900000 -5.300000 -8.730000 ;
      RECT -5.470000 38.730000 -5.300000 38.900000 ;
      RECT -5.110000 -8.900000 -4.940000 -8.730000 ;
      RECT -5.110000 38.730000 -4.940000 38.900000 ;
      RECT -4.750000 -8.900000 -4.580000 -8.730000 ;
      RECT -4.750000 38.730000 -4.580000 38.900000 ;
      RECT -4.390000 -8.900000 -4.220000 -8.730000 ;
      RECT -4.390000 38.730000 -4.220000 38.900000 ;
      RECT -4.030000 -8.900000 -3.860000 -8.730000 ;
      RECT -4.030000 38.730000 -3.860000 38.900000 ;
      RECT -3.870000 -3.280000 -3.700000 -3.110000 ;
      RECT -3.870000 -2.920000 -3.700000 -2.750000 ;
      RECT -3.870000 -2.560000 -3.700000 -2.390000 ;
      RECT -3.870000 -2.200000 -3.700000 -2.030000 ;
      RECT -3.870000 -1.840000 -3.700000 -1.670000 ;
      RECT -3.870000 -1.480000 -3.700000 -1.310000 ;
      RECT -3.870000 -1.120000 -3.700000 -0.950000 ;
      RECT -3.870000 -0.760000 -3.700000 -0.590000 ;
      RECT -3.870000 -0.400000 -3.700000 -0.230000 ;
      RECT -3.870000 -0.040000 -3.700000  0.130000 ;
      RECT -3.870000  0.320000 -3.700000  0.490000 ;
      RECT -3.870000  0.680000 -3.700000  0.850000 ;
      RECT -3.870000  1.040000 -3.700000  1.210000 ;
      RECT -3.870000  1.400000 -3.700000  1.570000 ;
      RECT -3.870000  1.760000 -3.700000  1.930000 ;
      RECT -3.870000  2.120000 -3.700000  2.290000 ;
      RECT -3.870000  2.480000 -3.700000  2.650000 ;
      RECT -3.870000  2.840000 -3.700000  3.010000 ;
      RECT -3.870000  3.200000 -3.700000  3.370000 ;
      RECT -3.870000  3.560000 -3.700000  3.730000 ;
      RECT -3.870000  3.920000 -3.700000  4.090000 ;
      RECT -3.870000  4.280000 -3.700000  4.450000 ;
      RECT -3.870000  4.640000 -3.700000  4.810000 ;
      RECT -3.870000  5.000000 -3.700000  5.170000 ;
      RECT -3.870000  5.360000 -3.700000  5.530000 ;
      RECT -3.870000  5.720000 -3.700000  5.890000 ;
      RECT -3.870000  6.080000 -3.700000  6.250000 ;
      RECT -3.870000  6.440000 -3.700000  6.610000 ;
      RECT -3.870000  6.800000 -3.700000  6.970000 ;
      RECT -3.870000  7.160000 -3.700000  7.330000 ;
      RECT -3.870000  7.520000 -3.700000  7.690000 ;
      RECT -3.870000  7.880000 -3.700000  8.050000 ;
      RECT -3.870000  8.240000 -3.700000  8.410000 ;
      RECT -3.870000  8.600000 -3.700000  8.770000 ;
      RECT -3.870000  8.960000 -3.700000  9.130000 ;
      RECT -3.870000  9.320000 -3.700000  9.490000 ;
      RECT -3.870000  9.680000 -3.700000  9.850000 ;
      RECT -3.870000 10.040000 -3.700000 10.210000 ;
      RECT -3.870000 10.400000 -3.700000 10.570000 ;
      RECT -3.870000 10.760000 -3.700000 10.930000 ;
      RECT -3.870000 11.120000 -3.700000 11.290000 ;
      RECT -3.870000 11.480000 -3.700000 11.650000 ;
      RECT -3.870000 11.840000 -3.700000 12.010000 ;
      RECT -3.870000 12.200000 -3.700000 12.370000 ;
      RECT -3.870000 12.560000 -3.700000 12.730000 ;
      RECT -3.870000 12.920000 -3.700000 13.090000 ;
      RECT -3.870000 13.280000 -3.700000 13.450000 ;
      RECT -3.870000 13.640000 -3.700000 13.810000 ;
      RECT -3.870000 14.000000 -3.700000 14.170000 ;
      RECT -3.870000 14.360000 -3.700000 14.530000 ;
      RECT -3.870000 14.720000 -3.700000 14.890000 ;
      RECT -3.870000 15.080000 -3.700000 15.250000 ;
      RECT -3.870000 15.440000 -3.700000 15.610000 ;
      RECT -3.870000 15.800000 -3.700000 15.970000 ;
      RECT -3.870000 16.160000 -3.700000 16.330000 ;
      RECT -3.870000 16.520000 -3.700000 16.690000 ;
      RECT -3.870000 16.880000 -3.700000 17.050000 ;
      RECT -3.870000 17.240000 -3.700000 17.410000 ;
      RECT -3.870000 17.600000 -3.700000 17.770000 ;
      RECT -3.870000 17.960000 -3.700000 18.130000 ;
      RECT -3.870000 18.320000 -3.700000 18.490000 ;
      RECT -3.870000 18.680000 -3.700000 18.850000 ;
      RECT -3.870000 19.040000 -3.700000 19.210000 ;
      RECT -3.870000 19.400000 -3.700000 19.570000 ;
      RECT -3.870000 19.760000 -3.700000 19.930000 ;
      RECT -3.870000 20.120000 -3.700000 20.290000 ;
      RECT -3.870000 20.480000 -3.700000 20.650000 ;
      RECT -3.870000 20.840000 -3.700000 21.010000 ;
      RECT -3.870000 21.200000 -3.700000 21.370000 ;
      RECT -3.870000 21.560000 -3.700000 21.730000 ;
      RECT -3.870000 21.920000 -3.700000 22.090000 ;
      RECT -3.870000 22.280000 -3.700000 22.450000 ;
      RECT -3.870000 22.640000 -3.700000 22.810000 ;
      RECT -3.870000 23.000000 -3.700000 23.170000 ;
      RECT -3.870000 23.360000 -3.700000 23.530000 ;
      RECT -3.870000 23.720000 -3.700000 23.890000 ;
      RECT -3.870000 24.080000 -3.700000 24.250000 ;
      RECT -3.870000 24.440000 -3.700000 24.610000 ;
      RECT -3.870000 24.800000 -3.700000 24.970000 ;
      RECT -3.870000 25.160000 -3.700000 25.330000 ;
      RECT -3.870000 25.520000 -3.700000 25.690000 ;
      RECT -3.870000 25.880000 -3.700000 26.050000 ;
      RECT -3.870000 26.240000 -3.700000 26.410000 ;
      RECT -3.870000 26.600000 -3.700000 26.770000 ;
      RECT -3.870000 26.960000 -3.700000 27.130000 ;
      RECT -3.870000 27.320000 -3.700000 27.490000 ;
      RECT -3.870000 27.680000 -3.700000 27.850000 ;
      RECT -3.870000 28.040000 -3.700000 28.210000 ;
      RECT -3.870000 28.400000 -3.700000 28.570000 ;
      RECT -3.870000 28.760000 -3.700000 28.930000 ;
      RECT -3.870000 29.120000 -3.700000 29.290000 ;
      RECT -3.870000 29.480000 -3.700000 29.650000 ;
      RECT -3.870000 29.840000 -3.700000 30.010000 ;
      RECT -3.870000 30.200000 -3.700000 30.370000 ;
      RECT -3.870000 30.560000 -3.700000 30.730000 ;
      RECT -3.870000 30.920000 -3.700000 31.090000 ;
      RECT -3.870000 31.280000 -3.700000 31.450000 ;
      RECT -3.870000 31.640000 -3.700000 31.810000 ;
      RECT -3.870000 32.000000 -3.700000 32.170000 ;
      RECT -3.870000 32.360000 -3.700000 32.530000 ;
      RECT -3.870000 32.720000 -3.700000 32.890000 ;
      RECT -3.870000 33.080000 -3.700000 33.250000 ;
      RECT -3.670000 -8.900000 -3.500000 -8.730000 ;
      RECT -3.670000 38.730000 -3.500000 38.900000 ;
      RECT -3.310000 -8.900000 -3.140000 -8.730000 ;
      RECT -3.310000 38.730000 -3.140000 38.900000 ;
      RECT -3.235000 -0.760000 -2.345000 30.730000 ;
      RECT -2.950000 -8.900000 -2.780000 -8.730000 ;
      RECT -2.950000 38.730000 -2.780000 38.900000 ;
      RECT -2.770000 -4.990000  3.520000 -4.100000 ;
      RECT -2.770000 34.100000  3.520000 34.990000 ;
      RECT -2.590000 -8.900000 -2.420000 -8.730000 ;
      RECT -2.590000 38.730000 -2.420000 38.900000 ;
      RECT -2.230000 -8.900000 -2.060000 -8.730000 ;
      RECT -2.230000 38.730000 -2.060000 38.900000 ;
      RECT -1.870000 -8.900000 -1.700000 -8.730000 ;
      RECT -1.870000 38.730000 -1.700000 38.900000 ;
      RECT -1.510000 -8.900000 -1.340000 -8.730000 ;
      RECT -1.510000 38.730000 -1.340000 38.900000 ;
      RECT -1.150000 -8.900000 -0.980000 -8.730000 ;
      RECT -1.150000 38.730000 -0.980000 38.900000 ;
      RECT -0.790000 -8.900000 -0.620000 -8.730000 ;
      RECT -0.790000 38.730000 -0.620000 38.900000 ;
      RECT -0.650000 -3.205000 -0.480000 -3.035000 ;
      RECT -0.650000 -2.835000 -0.480000 -2.665000 ;
      RECT -0.650000 -2.465000 -0.480000 -2.295000 ;
      RECT -0.610000 -0.760000  1.360000 30.730000 ;
      RECT -0.430000 -8.900000 -0.260000 -8.730000 ;
      RECT -0.430000 38.730000 -0.260000 38.900000 ;
      RECT -0.280000 -3.205000 -0.110000 -3.035000 ;
      RECT -0.280000 -2.835000 -0.110000 -2.665000 ;
      RECT -0.280000 -2.465000 -0.110000 -2.295000 ;
      RECT -0.070000 -8.900000  0.100000 -8.730000 ;
      RECT -0.070000 38.730000  0.100000 38.900000 ;
      RECT  0.090000 -3.205000  0.260000 -3.035000 ;
      RECT  0.090000 -2.835000  0.260000 -2.665000 ;
      RECT  0.090000 -2.465000  0.260000 -2.295000 ;
      RECT  0.290000 -8.900000  0.460000 -8.730000 ;
      RECT  0.290000 38.730000  0.460000 38.900000 ;
      RECT  0.460000 -3.205000  0.630000 -3.035000 ;
      RECT  0.460000 -2.835000  0.630000 -2.665000 ;
      RECT  0.460000 -2.465000  0.630000 -2.295000 ;
      RECT  0.650000 -8.900000  0.820000 -8.730000 ;
      RECT  0.650000 38.730000  0.820000 38.900000 ;
      RECT  0.830000 -3.205000  1.000000 -3.035000 ;
      RECT  0.830000 -2.835000  1.000000 -2.665000 ;
      RECT  0.830000 -2.465000  1.000000 -2.295000 ;
      RECT  1.010000 -8.900000  1.180000 -8.730000 ;
      RECT  1.010000 38.730000  1.180000 38.900000 ;
      RECT  1.200000 -3.205000  1.370000 -3.035000 ;
      RECT  1.200000 -2.835000  1.370000 -2.665000 ;
      RECT  1.200000 -2.465000  1.370000 -2.295000 ;
      RECT  1.370000 -8.900000  1.540000 -8.730000 ;
      RECT  1.370000 38.730000  1.540000 38.900000 ;
      RECT  1.730000 -8.900000  1.900000 -8.730000 ;
      RECT  1.730000 38.730000  1.900000 38.900000 ;
      RECT  2.090000 -8.900000  2.260000 -8.730000 ;
      RECT  2.090000 38.730000  2.260000 38.900000 ;
      RECT  2.450000 -8.900000  2.620000 -8.730000 ;
      RECT  2.450000 38.730000  2.620000 38.900000 ;
      RECT  2.810000 -8.900000  2.980000 -8.730000 ;
      RECT  2.810000 38.730000  2.980000 38.900000 ;
      RECT  3.095000 -0.760000  3.985000 30.730000 ;
      RECT  3.170000 -8.900000  3.340000 -8.730000 ;
      RECT  3.170000 38.730000  3.340000 38.900000 ;
      RECT  3.530000 -8.900000  3.700000 -8.730000 ;
      RECT  3.530000 38.730000  3.700000 38.900000 ;
      RECT  3.890000 -8.900000  4.060000 -8.730000 ;
      RECT  3.890000 38.730000  4.060000 38.900000 ;
      RECT  4.250000 -8.900000  4.420000 -8.730000 ;
      RECT  4.250000 38.730000  4.420000 38.900000 ;
      RECT  4.450000 -3.280000  4.620000 -3.110000 ;
      RECT  4.450000 -2.920000  4.620000 -2.750000 ;
      RECT  4.450000 -2.560000  4.620000 -2.390000 ;
      RECT  4.450000 -2.200000  4.620000 -2.030000 ;
      RECT  4.450000 -1.840000  4.620000 -1.670000 ;
      RECT  4.450000 -1.480000  4.620000 -1.310000 ;
      RECT  4.450000 -1.120000  4.620000 -0.950000 ;
      RECT  4.450000 -0.760000  4.620000 -0.590000 ;
      RECT  4.450000 -0.400000  4.620000 -0.230000 ;
      RECT  4.450000 -0.040000  4.620000  0.130000 ;
      RECT  4.450000  0.320000  4.620000  0.490000 ;
      RECT  4.450000  0.680000  4.620000  0.850000 ;
      RECT  4.450000  1.040000  4.620000  1.210000 ;
      RECT  4.450000  1.400000  4.620000  1.570000 ;
      RECT  4.450000  1.760000  4.620000  1.930000 ;
      RECT  4.450000  2.120000  4.620000  2.290000 ;
      RECT  4.450000  2.480000  4.620000  2.650000 ;
      RECT  4.450000  2.840000  4.620000  3.010000 ;
      RECT  4.450000  3.200000  4.620000  3.370000 ;
      RECT  4.450000  3.560000  4.620000  3.730000 ;
      RECT  4.450000  3.920000  4.620000  4.090000 ;
      RECT  4.450000  4.280000  4.620000  4.450000 ;
      RECT  4.450000  4.640000  4.620000  4.810000 ;
      RECT  4.450000  5.000000  4.620000  5.170000 ;
      RECT  4.450000  5.360000  4.620000  5.530000 ;
      RECT  4.450000  5.720000  4.620000  5.890000 ;
      RECT  4.450000  6.080000  4.620000  6.250000 ;
      RECT  4.450000  6.440000  4.620000  6.610000 ;
      RECT  4.450000  6.800000  4.620000  6.970000 ;
      RECT  4.450000  7.160000  4.620000  7.330000 ;
      RECT  4.450000  7.520000  4.620000  7.690000 ;
      RECT  4.450000  7.880000  4.620000  8.050000 ;
      RECT  4.450000  8.240000  4.620000  8.410000 ;
      RECT  4.450000  8.600000  4.620000  8.770000 ;
      RECT  4.450000  8.960000  4.620000  9.130000 ;
      RECT  4.450000  9.320000  4.620000  9.490000 ;
      RECT  4.450000  9.680000  4.620000  9.850000 ;
      RECT  4.450000 10.040000  4.620000 10.210000 ;
      RECT  4.450000 10.400000  4.620000 10.570000 ;
      RECT  4.450000 10.760000  4.620000 10.930000 ;
      RECT  4.450000 11.120000  4.620000 11.290000 ;
      RECT  4.450000 11.480000  4.620000 11.650000 ;
      RECT  4.450000 11.840000  4.620000 12.010000 ;
      RECT  4.450000 12.200000  4.620000 12.370000 ;
      RECT  4.450000 12.560000  4.620000 12.730000 ;
      RECT  4.450000 12.920000  4.620000 13.090000 ;
      RECT  4.450000 13.280000  4.620000 13.450000 ;
      RECT  4.450000 13.640000  4.620000 13.810000 ;
      RECT  4.450000 14.000000  4.620000 14.170000 ;
      RECT  4.450000 14.360000  4.620000 14.530000 ;
      RECT  4.450000 14.720000  4.620000 14.890000 ;
      RECT  4.450000 15.080000  4.620000 15.250000 ;
      RECT  4.450000 15.440000  4.620000 15.610000 ;
      RECT  4.450000 15.800000  4.620000 15.970000 ;
      RECT  4.450000 16.160000  4.620000 16.330000 ;
      RECT  4.450000 16.520000  4.620000 16.690000 ;
      RECT  4.450000 16.880000  4.620000 17.050000 ;
      RECT  4.450000 17.240000  4.620000 17.410000 ;
      RECT  4.450000 17.600000  4.620000 17.770000 ;
      RECT  4.450000 17.960000  4.620000 18.130000 ;
      RECT  4.450000 18.320000  4.620000 18.490000 ;
      RECT  4.450000 18.680000  4.620000 18.850000 ;
      RECT  4.450000 19.040000  4.620000 19.210000 ;
      RECT  4.450000 19.400000  4.620000 19.570000 ;
      RECT  4.450000 19.760000  4.620000 19.930000 ;
      RECT  4.450000 20.120000  4.620000 20.290000 ;
      RECT  4.450000 20.480000  4.620000 20.650000 ;
      RECT  4.450000 20.840000  4.620000 21.010000 ;
      RECT  4.450000 21.200000  4.620000 21.370000 ;
      RECT  4.450000 21.560000  4.620000 21.730000 ;
      RECT  4.450000 21.920000  4.620000 22.090000 ;
      RECT  4.450000 22.280000  4.620000 22.450000 ;
      RECT  4.450000 22.640000  4.620000 22.810000 ;
      RECT  4.450000 23.000000  4.620000 23.170000 ;
      RECT  4.450000 23.360000  4.620000 23.530000 ;
      RECT  4.450000 23.720000  4.620000 23.890000 ;
      RECT  4.450000 24.080000  4.620000 24.250000 ;
      RECT  4.450000 24.440000  4.620000 24.610000 ;
      RECT  4.450000 24.800000  4.620000 24.970000 ;
      RECT  4.450000 25.160000  4.620000 25.330000 ;
      RECT  4.450000 25.520000  4.620000 25.690000 ;
      RECT  4.450000 25.880000  4.620000 26.050000 ;
      RECT  4.450000 26.240000  4.620000 26.410000 ;
      RECT  4.450000 26.600000  4.620000 26.770000 ;
      RECT  4.450000 26.960000  4.620000 27.130000 ;
      RECT  4.450000 27.320000  4.620000 27.490000 ;
      RECT  4.450000 27.680000  4.620000 27.850000 ;
      RECT  4.450000 28.040000  4.620000 28.210000 ;
      RECT  4.450000 28.400000  4.620000 28.570000 ;
      RECT  4.450000 28.760000  4.620000 28.930000 ;
      RECT  4.450000 29.120000  4.620000 29.290000 ;
      RECT  4.450000 29.480000  4.620000 29.650000 ;
      RECT  4.450000 29.840000  4.620000 30.010000 ;
      RECT  4.450000 30.200000  4.620000 30.370000 ;
      RECT  4.450000 30.560000  4.620000 30.730000 ;
      RECT  4.450000 30.920000  4.620000 31.090000 ;
      RECT  4.450000 31.280000  4.620000 31.450000 ;
      RECT  4.450000 31.640000  4.620000 31.810000 ;
      RECT  4.450000 32.000000  4.620000 32.170000 ;
      RECT  4.450000 32.360000  4.620000 32.530000 ;
      RECT  4.450000 32.720000  4.620000 32.890000 ;
      RECT  4.450000 33.080000  4.620000 33.250000 ;
      RECT  4.610000 -8.900000  4.780000 -8.730000 ;
      RECT  4.610000 38.730000  4.780000 38.900000 ;
      RECT  4.970000 -8.900000  5.140000 -8.730000 ;
      RECT  4.970000 38.730000  5.140000 38.900000 ;
      RECT  5.330000 -8.900000  5.500000 -8.730000 ;
      RECT  5.330000 38.730000  5.500000 38.900000 ;
      RECT  5.690000 -8.900000  5.860000 -8.730000 ;
      RECT  5.690000 38.730000  5.860000 38.900000 ;
      RECT  6.050000 -8.900000  6.220000 -8.730000 ;
      RECT  6.050000 38.730000  6.220000 38.900000 ;
      RECT  6.410000 -8.900000  6.580000 -8.730000 ;
      RECT  6.410000 38.730000  6.580000 38.900000 ;
      RECT  6.770000 -8.900000  6.940000 -8.730000 ;
      RECT  6.770000 38.730000  6.940000 38.900000 ;
      RECT  7.130000 -8.900000  7.300000 -8.730000 ;
      RECT  7.130000 38.730000  7.300000 38.900000 ;
      RECT  7.490000 -8.900000  7.660000 -8.730000 ;
      RECT  7.490000 38.730000  7.660000 38.900000 ;
      RECT  7.850000 -8.900000  8.020000 -8.730000 ;
      RECT  7.850000 38.730000  8.020000 38.900000 ;
      RECT  8.360000 -8.305000  8.530000 -8.135000 ;
      RECT  8.360000 -7.945000  8.530000 -7.775000 ;
      RECT  8.360000 -7.585000  8.530000 -7.415000 ;
      RECT  8.360000 -7.225000  8.530000 -7.055000 ;
      RECT  8.360000 -6.865000  8.530000 -6.695000 ;
      RECT  8.360000 -6.505000  8.530000 -6.335000 ;
      RECT  8.360000 -6.145000  8.530000 -5.975000 ;
      RECT  8.360000 -5.785000  8.530000 -5.615000 ;
      RECT  8.360000 -5.425000  8.530000 -5.255000 ;
      RECT  8.360000 -5.065000  8.530000 -4.895000 ;
      RECT  8.360000 -4.705000  8.530000 -4.535000 ;
      RECT  8.360000 -4.345000  8.530000 -4.175000 ;
      RECT  8.360000 -3.985000  8.530000 -3.815000 ;
      RECT  8.360000 -3.625000  8.530000 -3.455000 ;
      RECT  8.360000 -3.265000  8.530000 -3.095000 ;
      RECT  8.360000 -2.905000  8.530000 -2.735000 ;
      RECT  8.360000 -2.545000  8.530000 -2.375000 ;
      RECT  8.360000 -2.185000  8.530000 -2.015000 ;
      RECT  8.360000 -1.825000  8.530000 -1.655000 ;
      RECT  8.360000 -1.465000  8.530000 -1.295000 ;
      RECT  8.360000 -1.105000  8.530000 -0.935000 ;
      RECT  8.360000 -0.745000  8.530000 -0.575000 ;
      RECT  8.360000 -0.385000  8.530000 -0.215000 ;
      RECT  8.360000 -0.025000  8.530000  0.145000 ;
      RECT  8.360000  0.335000  8.530000  0.505000 ;
      RECT  8.360000  0.695000  8.530000  0.865000 ;
      RECT  8.360000  1.055000  8.530000  1.225000 ;
      RECT  8.360000  1.415000  8.530000  1.585000 ;
      RECT  8.360000  1.775000  8.530000  1.945000 ;
      RECT  8.360000  2.135000  8.530000  2.305000 ;
      RECT  8.360000  2.495000  8.530000  2.665000 ;
      RECT  8.360000  2.855000  8.530000  3.025000 ;
      RECT  8.360000  3.215000  8.530000  3.385000 ;
      RECT  8.360000  3.575000  8.530000  3.745000 ;
      RECT  8.360000  3.935000  8.530000  4.105000 ;
      RECT  8.360000  4.295000  8.530000  4.465000 ;
      RECT  8.360000  4.655000  8.530000  4.825000 ;
      RECT  8.360000  5.015000  8.530000  5.185000 ;
      RECT  8.360000  5.375000  8.530000  5.545000 ;
      RECT  8.360000  5.735000  8.530000  5.905000 ;
      RECT  8.360000  6.095000  8.530000  6.265000 ;
      RECT  8.360000  6.455000  8.530000  6.625000 ;
      RECT  8.360000  6.815000  8.530000  6.985000 ;
      RECT  8.360000  7.175000  8.530000  7.345000 ;
      RECT  8.360000  7.535000  8.530000  7.705000 ;
      RECT  8.360000  7.895000  8.530000  8.065000 ;
      RECT  8.360000  8.255000  8.530000  8.425000 ;
      RECT  8.360000  8.615000  8.530000  8.785000 ;
      RECT  8.360000  8.975000  8.530000  9.145000 ;
      RECT  8.360000  9.335000  8.530000  9.505000 ;
      RECT  8.360000  9.695000  8.530000  9.865000 ;
      RECT  8.360000 10.055000  8.530000 10.225000 ;
      RECT  8.360000 10.415000  8.530000 10.585000 ;
      RECT  8.360000 10.775000  8.530000 10.945000 ;
      RECT  8.360000 11.135000  8.530000 11.305000 ;
      RECT  8.360000 11.495000  8.530000 11.665000 ;
      RECT  8.360000 11.855000  8.530000 12.025000 ;
      RECT  8.360000 12.215000  8.530000 12.385000 ;
      RECT  8.360000 12.575000  8.530000 12.745000 ;
      RECT  8.360000 12.935000  8.530000 13.105000 ;
      RECT  8.360000 13.295000  8.530000 13.465000 ;
      RECT  8.360000 13.655000  8.530000 13.825000 ;
      RECT  8.360000 14.015000  8.530000 14.185000 ;
      RECT  8.360000 14.375000  8.530000 14.545000 ;
      RECT  8.360000 14.735000  8.530000 14.905000 ;
      RECT  8.360000 15.095000  8.530000 15.265000 ;
      RECT  8.360000 15.455000  8.530000 15.625000 ;
      RECT  8.360000 15.815000  8.530000 15.985000 ;
      RECT  8.360000 16.175000  8.530000 16.345000 ;
      RECT  8.360000 16.535000  8.530000 16.705000 ;
      RECT  8.360000 16.895000  8.530000 17.065000 ;
      RECT  8.360000 17.255000  8.530000 17.425000 ;
      RECT  8.360000 17.615000  8.530000 17.785000 ;
      RECT  8.360000 17.975000  8.530000 18.145000 ;
      RECT  8.360000 18.335000  8.530000 18.505000 ;
      RECT  8.360000 18.695000  8.530000 18.865000 ;
      RECT  8.360000 19.055000  8.530000 19.225000 ;
      RECT  8.360000 19.415000  8.530000 19.585000 ;
      RECT  8.360000 19.775000  8.530000 19.945000 ;
      RECT  8.360000 20.135000  8.530000 20.305000 ;
      RECT  8.360000 20.495000  8.530000 20.665000 ;
      RECT  8.360000 20.855000  8.530000 21.025000 ;
      RECT  8.360000 21.215000  8.530000 21.385000 ;
      RECT  8.360000 21.575000  8.530000 21.745000 ;
      RECT  8.360000 21.935000  8.530000 22.105000 ;
      RECT  8.360000 22.295000  8.530000 22.465000 ;
      RECT  8.360000 22.655000  8.530000 22.825000 ;
      RECT  8.360000 23.015000  8.530000 23.185000 ;
      RECT  8.360000 23.375000  8.530000 23.545000 ;
      RECT  8.360000 23.735000  8.530000 23.905000 ;
      RECT  8.360000 24.095000  8.530000 24.265000 ;
      RECT  8.360000 24.455000  8.530000 24.625000 ;
      RECT  8.360000 24.815000  8.530000 24.985000 ;
      RECT  8.360000 25.175000  8.530000 25.345000 ;
      RECT  8.360000 25.535000  8.530000 25.705000 ;
      RECT  8.360000 25.895000  8.530000 26.065000 ;
      RECT  8.360000 26.255000  8.530000 26.425000 ;
      RECT  8.360000 26.615000  8.530000 26.785000 ;
      RECT  8.360000 26.975000  8.530000 27.145000 ;
      RECT  8.360000 27.335000  8.530000 27.505000 ;
      RECT  8.360000 27.695000  8.530000 27.865000 ;
      RECT  8.360000 28.055000  8.530000 28.225000 ;
      RECT  8.360000 28.415000  8.530000 28.585000 ;
      RECT  8.360000 28.775000  8.530000 28.945000 ;
      RECT  8.360000 29.135000  8.530000 29.305000 ;
      RECT  8.360000 29.495000  8.530000 29.665000 ;
      RECT  8.360000 29.855000  8.530000 30.025000 ;
      RECT  8.360000 30.215000  8.530000 30.385000 ;
      RECT  8.360000 30.575000  8.530000 30.745000 ;
      RECT  8.360000 30.935000  8.530000 31.105000 ;
      RECT  8.360000 31.295000  8.530000 31.465000 ;
      RECT  8.360000 31.655000  8.530000 31.825000 ;
      RECT  8.360000 32.015000  8.530000 32.185000 ;
      RECT  8.360000 32.375000  8.530000 32.545000 ;
      RECT  8.360000 32.735000  8.530000 32.905000 ;
      RECT  8.360000 33.095000  8.530000 33.265000 ;
      RECT  8.360000 33.455000  8.530000 33.625000 ;
      RECT  8.360000 33.815000  8.530000 33.985000 ;
      RECT  8.360000 34.175000  8.530000 34.345000 ;
      RECT  8.360000 34.535000  8.530000 34.705000 ;
      RECT  8.360000 34.895000  8.530000 35.065000 ;
      RECT  8.360000 35.255000  8.530000 35.425000 ;
      RECT  8.360000 35.615000  8.530000 35.785000 ;
      RECT  8.360000 35.975000  8.530000 36.145000 ;
      RECT  8.360000 36.335000  8.530000 36.505000 ;
      RECT  8.360000 36.695000  8.530000 36.865000 ;
      RECT  8.360000 37.055000  8.530000 37.225000 ;
      RECT  8.360000 37.415000  8.530000 37.585000 ;
      RECT  8.360000 37.775000  8.530000 37.945000 ;
      RECT  8.360000 38.135000  8.530000 38.305000 ;
    LAYER met1 ;
      RECT -7.900000 -9.020000  8.650000 -8.610000 ;
      RECT -7.900000 -8.610000 -7.490000 38.610000 ;
      RECT -7.900000 38.610000  8.650000 39.020000 ;
      RECT -3.990000 -5.110000  4.740000 -3.785000 ;
      RECT -3.990000 -3.785000 -3.580000 33.785000 ;
      RECT -3.990000 33.785000  4.740000 35.110000 ;
      RECT -3.295000 -0.820000 -2.285000 30.825000 ;
      RECT -0.730000 -3.285000  1.450000 -2.215000 ;
      RECT -0.670000 -0.820000  1.420000 30.825000 ;
      RECT  3.035000 -0.820000  4.045000 30.825000 ;
      RECT  4.330000 -3.785000  4.740000 33.785000 ;
      RECT  8.240000 -8.610000  8.650000 38.610000 ;
    LAYER met2 ;
      RECT -3.295000 -5.610000 -2.285000 30.825000 ;
      RECT -0.730000 -3.285000  1.450000 -2.215000 ;
      RECT -0.670000 -0.820000  1.420000 35.610000 ;
      RECT  3.035000 -5.610000  4.045000 30.825000 ;
    LAYER met3 ;
      RECT -0.750000 -3.285000 1.450000 -2.215000 ;
    LAYER via ;
      RECT -3.240000 -0.665000 -2.340000 30.635000 ;
      RECT -0.695000 -3.250000 -0.435000 -2.990000 ;
      RECT -0.695000 -2.880000 -0.435000 -2.620000 ;
      RECT -0.695000 -2.510000 -0.435000 -2.250000 ;
      RECT -0.555000 -0.665000  1.305000 30.635000 ;
      RECT -0.325000 -3.250000 -0.065000 -2.990000 ;
      RECT -0.325000 -2.880000 -0.065000 -2.620000 ;
      RECT -0.325000 -2.510000 -0.065000 -2.250000 ;
      RECT  0.045000 -3.250000  0.305000 -2.990000 ;
      RECT  0.045000 -2.880000  0.305000 -2.620000 ;
      RECT  0.045000 -2.510000  0.305000 -2.250000 ;
      RECT  0.415000 -3.250000  0.675000 -2.990000 ;
      RECT  0.415000 -2.880000  0.675000 -2.620000 ;
      RECT  0.415000 -2.510000  0.675000 -2.250000 ;
      RECT  0.785000 -3.250000  1.045000 -2.990000 ;
      RECT  0.785000 -2.880000  1.045000 -2.620000 ;
      RECT  0.785000 -2.510000  1.045000 -2.250000 ;
      RECT  1.155000 -3.250000  1.415000 -2.990000 ;
      RECT  1.155000 -2.880000  1.415000 -2.620000 ;
      RECT  1.155000 -2.510000  1.415000 -2.250000 ;
      RECT  3.090000 -0.665000  3.990000 30.635000 ;
    LAYER via2 ;
      RECT -0.580000 -3.075000 1.300000 -2.395000 ;
  END
END sky130_fd_pr__rf_pfet_20v0_withptap
END LIBRARY
