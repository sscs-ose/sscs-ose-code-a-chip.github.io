# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2 ;
  ORIGIN  0.440000  0.000000 ;
  SIZE  4.380000 BY  4.590000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT -0.440000 0.000000  3.940000 0.320000 ;
        RECT -0.440000 0.320000 -0.170000 4.130000 ;
        RECT  0.280000 0.320000  0.420000 4.130000 ;
        RECT  0.840000 0.320000  0.980000 4.130000 ;
        RECT  1.400000 0.320000  1.540000 4.130000 ;
        RECT  1.960000 0.320000  2.100000 4.130000 ;
        RECT  2.520000 0.320000  2.660000 4.130000 ;
        RECT  3.080000 0.320000  3.220000 4.130000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT -0.440000 4.270000 3.940000 4.590000 ;
        RECT  0.000000 0.460000 0.140000 4.270000 ;
        RECT  0.560000 0.460000 0.700000 4.270000 ;
        RECT  1.120000 0.460000 1.260000 4.270000 ;
        RECT  1.680000 0.460000 1.820000 4.270000 ;
        RECT  2.240000 0.460000 2.380000 4.270000 ;
        RECT  2.800000 0.460000 2.940000 4.270000 ;
        RECT  3.360000 0.460000 3.500000 4.270000 ;
        RECT  3.670000 0.460000 3.940000 4.270000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 1.850000 2.430000 1.930000 2.515000 ;
    END
  END SUB
  OBS
    LAYER met1 ;
      RECT -0.440000 0.000000  3.940000 0.320000 ;
      RECT -0.440000 0.320000 -0.170000 4.130000 ;
      RECT -0.440000 4.270000  3.940000 4.590000 ;
      RECT  0.000000 0.320000  0.140000 4.130000 ;
      RECT  0.280000 0.460000  0.420000 4.270000 ;
      RECT  0.560000 0.320000  0.700000 4.130000 ;
      RECT  0.840000 0.460000  0.980000 4.270000 ;
      RECT  1.120000 0.320000  1.260000 4.130000 ;
      RECT  1.400000 0.460000  1.540000 4.270000 ;
      RECT  1.680000 0.320000  1.820000 4.130000 ;
      RECT  1.960000 0.460000  2.100000 4.270000 ;
      RECT  2.240000 0.320000  2.380000 4.130000 ;
      RECT  2.520000 0.460000  2.660000 4.270000 ;
      RECT  2.800000 0.320000  2.940000 4.130000 ;
      RECT  3.080000 0.460000  3.220000 4.270000 ;
      RECT  3.360000 0.320000  3.500000 4.130000 ;
      RECT  3.670000 0.460000  3.940000 4.270000 ;
    LAYER via ;
      RECT -0.435000 0.265000 -0.175000 0.525000 ;
      RECT -0.435000 0.585000 -0.175000 0.845000 ;
      RECT -0.435000 0.905000 -0.175000 1.165000 ;
      RECT -0.435000 1.225000 -0.175000 1.485000 ;
      RECT -0.435000 1.545000 -0.175000 1.805000 ;
      RECT -0.435000 1.865000 -0.175000 2.125000 ;
      RECT -0.435000 2.185000 -0.175000 2.445000 ;
      RECT -0.435000 2.505000 -0.175000 2.765000 ;
      RECT -0.435000 2.825000 -0.175000 3.085000 ;
      RECT -0.435000 3.145000 -0.175000 3.405000 ;
      RECT -0.435000 3.465000 -0.175000 3.725000 ;
      RECT -0.435000 3.785000 -0.175000 4.045000 ;
      RECT -0.060000 0.030000  0.200000 0.290000 ;
      RECT -0.060000 4.300000  0.200000 4.560000 ;
      RECT  0.260000 0.030000  0.520000 0.290000 ;
      RECT  0.260000 4.300000  0.520000 4.560000 ;
      RECT  0.580000 0.030000  0.840000 0.290000 ;
      RECT  0.580000 4.300000  0.840000 4.560000 ;
      RECT  0.900000 0.030000  1.160000 0.290000 ;
      RECT  0.900000 4.300000  1.160000 4.560000 ;
      RECT  1.220000 0.030000  1.480000 0.290000 ;
      RECT  1.220000 4.300000  1.480000 4.560000 ;
      RECT  1.540000 0.030000  1.800000 0.290000 ;
      RECT  1.540000 4.300000  1.800000 4.560000 ;
      RECT  1.860000 0.030000  2.120000 0.290000 ;
      RECT  1.860000 4.300000  2.120000 4.560000 ;
      RECT  2.180000 0.030000  2.440000 0.290000 ;
      RECT  2.180000 4.300000  2.440000 4.560000 ;
      RECT  2.500000 0.030000  2.760000 0.290000 ;
      RECT  2.500000 4.300000  2.760000 4.560000 ;
      RECT  2.820000 0.030000  3.080000 0.290000 ;
      RECT  2.820000 4.300000  3.080000 4.560000 ;
      RECT  3.140000 0.030000  3.400000 0.290000 ;
      RECT  3.140000 4.300000  3.400000 4.560000 ;
      RECT  3.675000 0.490000  3.935000 0.750000 ;
      RECT  3.675000 0.810000  3.935000 1.070000 ;
      RECT  3.675000 1.130000  3.935000 1.390000 ;
      RECT  3.675000 1.450000  3.935000 1.710000 ;
      RECT  3.675000 1.770000  3.935000 2.030000 ;
      RECT  3.675000 2.090000  3.935000 2.350000 ;
      RECT  3.675000 2.410000  3.935000 2.670000 ;
      RECT  3.675000 2.730000  3.935000 2.990000 ;
      RECT  3.675000 3.050000  3.935000 3.310000 ;
      RECT  3.675000 3.370000  3.935000 3.630000 ;
      RECT  3.675000 3.690000  3.935000 3.950000 ;
  END
END sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2
END LIBRARY
