# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF06W1p65L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF06W1p65L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  2.860000 BY  2.760000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.386000 ;
    PORT
      LAYER met3 ;
        RECT 0.585000 1.015000 0.915000 1.455000 ;
        RECT 0.585000 1.455000 2.635000 1.785000 ;
        RECT 1.445000 1.015000 1.775000 1.455000 ;
        RECT 2.305000 1.015000 2.635000 1.455000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.485000 ;
    PORT
      LAYER met1 ;
        RECT 0.565000 2.005000 2.655000 2.295000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.848000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 3.015000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  1.785000 ;
        RECT 1.065000 -0.145000 1.295000  1.785000 ;
        RECT 1.925000 -0.145000 2.155000  1.785000 ;
        RECT 2.785000 -0.145000 3.015000  1.785000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.395000 1.850000 0.445000 1.935000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.255000 0.405000 1.785000 ;
      RECT 0.595000 1.985000 2.625000 2.315000 ;
      RECT 0.665000 0.255000 0.835000 1.785000 ;
      RECT 1.095000 0.255000 1.265000 1.785000 ;
      RECT 1.525000 0.255000 1.695000 1.785000 ;
      RECT 1.955000 0.255000 2.125000 1.785000 ;
      RECT 2.385000 0.255000 2.555000 1.785000 ;
      RECT 2.815000 0.255000 2.985000 1.785000 ;
    LAYER mcon ;
      RECT 0.235000 0.395000 0.405000 0.565000 ;
      RECT 0.235000 0.755000 0.405000 0.925000 ;
      RECT 0.235000 1.115000 0.405000 1.285000 ;
      RECT 0.235000 1.475000 0.405000 1.645000 ;
      RECT 0.625000 2.065000 0.795000 2.235000 ;
      RECT 0.665000 0.395000 0.835000 0.565000 ;
      RECT 0.665000 0.755000 0.835000 0.925000 ;
      RECT 0.665000 1.115000 0.835000 1.285000 ;
      RECT 0.665000 1.475000 0.835000 1.645000 ;
      RECT 0.985000 2.065000 1.155000 2.235000 ;
      RECT 1.095000 0.395000 1.265000 0.565000 ;
      RECT 1.095000 0.755000 1.265000 0.925000 ;
      RECT 1.095000 1.115000 1.265000 1.285000 ;
      RECT 1.095000 1.475000 1.265000 1.645000 ;
      RECT 1.345000 2.065000 1.515000 2.235000 ;
      RECT 1.525000 0.395000 1.695000 0.565000 ;
      RECT 1.525000 0.755000 1.695000 0.925000 ;
      RECT 1.525000 1.115000 1.695000 1.285000 ;
      RECT 1.525000 1.475000 1.695000 1.645000 ;
      RECT 1.705000 2.065000 1.875000 2.235000 ;
      RECT 1.955000 0.395000 2.125000 0.565000 ;
      RECT 1.955000 0.755000 2.125000 0.925000 ;
      RECT 1.955000 1.115000 2.125000 1.285000 ;
      RECT 1.955000 1.475000 2.125000 1.645000 ;
      RECT 2.065000 2.065000 2.235000 2.235000 ;
      RECT 2.385000 0.395000 2.555000 0.565000 ;
      RECT 2.385000 0.755000 2.555000 0.925000 ;
      RECT 2.385000 1.115000 2.555000 1.285000 ;
      RECT 2.385000 1.475000 2.555000 1.645000 ;
      RECT 2.425000 2.065000 2.595000 2.235000 ;
      RECT 2.815000 0.395000 2.985000 0.565000 ;
      RECT 2.815000 0.755000 2.985000 0.925000 ;
      RECT 2.815000 1.115000 2.985000 1.285000 ;
      RECT 2.815000 1.475000 2.985000 1.645000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 1.785000 ;
      RECT 1.480000 0.255000 1.740000 1.785000 ;
      RECT 2.340000 0.255000 2.600000 1.785000 ;
    LAYER met2 ;
      RECT 0.585000 1.015000 0.915000 1.785000 ;
      RECT 1.445000 1.015000 1.775000 1.785000 ;
      RECT 2.305000 1.015000 2.635000 1.785000 ;
    LAYER via ;
      RECT 0.620000 1.110000 0.880000 1.370000 ;
      RECT 0.620000 1.430000 0.880000 1.690000 ;
      RECT 1.480000 1.110000 1.740000 1.370000 ;
      RECT 1.480000 1.430000 1.740000 1.690000 ;
      RECT 2.340000 1.110000 2.600000 1.370000 ;
      RECT 2.340000 1.430000 2.600000 1.690000 ;
    LAYER via2 ;
      RECT 0.610000 1.060000 0.890000 1.340000 ;
      RECT 0.610000 1.460000 0.890000 1.740000 ;
      RECT 1.470000 1.060000 1.750000 1.340000 ;
      RECT 1.470000 1.460000 1.750000 1.740000 ;
      RECT 2.330000 1.060000 2.610000 1.340000 ;
      RECT 2.330000 1.460000 2.610000 1.740000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF06W1p65L0p15
END LIBRARY
