** sch_path: /home/evadeltor/OpenSourceAMS/NAND.sch
**.subckt NAND
**.ends
.end
