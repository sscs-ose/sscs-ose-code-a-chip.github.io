# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__esd_rf_nfet_20v0_hbm_32vW60p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__esd_rf_nfet_20v0_hbm_32vW60p00 ;
  ORIGIN  6.040000  5.910000 ;
  SIZE  13.58000 BY  41.82000 ;
  OBS
    LAYER li1 ;
      RECT -6.040000 -5.910000  7.540000 -4.470000 ;
      RECT -6.040000 -4.470000 -4.480000 34.350000 ;
      RECT -6.040000 34.350000  7.540000 35.910000 ;
      RECT -0.950000 -4.470000  2.445000 -3.255000 ;
      RECT -0.945000 -3.255000  2.445000 -3.245000 ;
      RECT  0.000000  0.000000  1.500000 30.000000 ;
      RECT  5.980000 -4.470000  7.540000 34.350000 ;
    LAYER mcon ;
      RECT -5.810000 -5.785000 -4.560000 35.785000 ;
      RECT -4.195000 -5.785000  5.695000 -4.535000 ;
      RECT -4.195000 34.535000  5.695000 35.785000 ;
      RECT  0.125000  0.155000  1.375000 29.845000 ;
      RECT  6.060000 -5.785000  7.310000 35.785000 ;
    LAYER met1 ;
      POLYGON -3.545000 -1.740000 -3.035000 -2.250000 -3.545000 -2.250000 ;
      POLYGON -3.545000 32.250000 -3.035000 32.250000 -3.545000 31.740000 ;
      POLYGON -3.035000 -2.250000 -1.785000 -3.500000 -3.035000 -3.500000 ;
      POLYGON -3.035000 33.500000 -1.785000 33.500000 -3.035000 32.250000 ;
      POLYGON -2.245000 -1.870000 -2.155000 -1.870000 -2.155000 -1.960000 ;
      POLYGON -2.155000 -1.960000 -1.865000 -1.960000 -1.865000 -2.250000 ;
      POLYGON -2.155000 31.960000 -2.155000 31.870000 -2.245000 31.870000 ;
      POLYGON -1.865000 32.250000 -1.865000 31.960000 -2.155000 31.960000 ;
      POLYGON  3.290000 33.500000  4.540000 33.500000  4.540000 32.250000 ;
      POLYGON  3.370000 -1.960000  3.660000 -1.960000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.660000 31.960000  3.370000 31.960000 ;
      POLYGON  3.660000 -1.870000  3.750000 -1.870000  3.660000 -1.960000 ;
      POLYGON  3.660000 31.960000  3.750000 31.870000  3.660000 31.870000 ;
      POLYGON  4.540000 -2.250000  4.540000 -3.500000  3.290000 -3.500000 ;
      POLYGON  4.540000 32.250000  4.830000 32.250000  4.830000 31.960000 ;
      POLYGON  4.830000 -1.960000  4.830000 -2.250000  4.540000 -2.250000 ;
      POLYGON  4.830000 31.960000  5.050000 31.960000  5.050000 31.740000 ;
      POLYGON  5.050000 -1.740000  5.050000 -1.960000  4.830000 -1.960000 ;
      RECT -6.040000 -5.910000  7.540000 -3.500000 ;
      RECT -6.040000 -3.500000 -3.035000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.545000 32.250000 ;
      RECT -6.040000 32.250000 -3.035000 33.500000 ;
      RECT -6.040000 33.500000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.155000 -1.960000  3.660000 -1.870000 ;
      RECT -2.155000 31.870000  3.660000 31.960000 ;
      RECT -1.865000 -2.250000  3.370000 -1.960000 ;
      RECT -1.865000 31.960000  3.370000 32.250000 ;
      RECT  4.540000 -3.500000  7.540000 -2.250000 ;
      RECT  4.540000 32.250000  7.540000 33.500000 ;
      RECT  4.830000 -2.250000  7.540000 -1.960000 ;
      RECT  4.830000 31.960000  7.540000 32.250000 ;
      RECT  5.050000 -1.960000  7.540000 31.960000 ;
    LAYER met2 ;
      POLYGON -3.545000 -1.740000 -3.035000 -2.250000 -3.545000 -2.250000 ;
      POLYGON -3.545000 32.250000 -3.035000 32.250000 -3.545000 31.740000 ;
      POLYGON -3.035000 -2.250000 -1.785000 -3.500000 -3.035000 -3.500000 ;
      POLYGON -3.035000 33.500000 -1.785000 33.500000 -3.035000 32.250000 ;
      POLYGON -2.245000 -1.870000 -2.130000 -1.870000 -2.130000 -1.985000 ;
      POLYGON -2.130000 -1.985000 -1.865000 -1.985000 -1.865000 -2.250000 ;
      POLYGON -2.130000 31.985000 -2.130000 31.870000 -2.245000 31.870000 ;
      POLYGON -1.865000 32.250000 -1.865000 31.985000 -2.130000 31.985000 ;
      POLYGON  3.290000 33.500000  4.540000 33.500000  4.540000 32.250000 ;
      POLYGON  3.370000 -1.985000  3.635000 -1.985000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.635000 31.985000  3.370000 31.985000 ;
      POLYGON  3.635000 -1.870000  3.750000 -1.870000  3.635000 -1.985000 ;
      POLYGON  3.635000 31.985000  3.750000 31.870000  3.635000 31.870000 ;
      POLYGON  4.540000 -2.250000  4.540000 -3.500000  3.290000 -3.500000 ;
      POLYGON  4.540000 32.250000  4.805000 32.250000  4.805000 31.985000 ;
      POLYGON  4.805000 -1.985000  4.805000 -2.250000  4.540000 -2.250000 ;
      POLYGON  4.805000 31.985000  5.050000 31.985000  5.050000 31.740000 ;
      POLYGON  5.050000 -1.740000  5.050000 -1.985000  4.805000 -1.985000 ;
      RECT -6.040000 -5.910000  7.540000 -3.500000 ;
      RECT -6.040000 -3.500000 -3.035000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.545000 32.250000 ;
      RECT -6.040000 32.250000 -3.035000 33.500000 ;
      RECT -6.040000 33.500000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.130000 -1.985000  3.635000 -1.870000 ;
      RECT -2.130000 31.870000  3.635000 31.985000 ;
      RECT -1.865000 -2.250000  3.370000 -1.985000 ;
      RECT -1.865000 31.985000  3.370000 32.250000 ;
      RECT  4.540000 -3.500000  7.540000 -2.250000 ;
      RECT  4.540000 32.250000  7.540000 33.500000 ;
      RECT  4.805000 -2.250000  7.540000 -1.985000 ;
      RECT  4.805000 31.985000  7.540000 32.250000 ;
      RECT  5.050000 -1.985000  7.540000 31.985000 ;
    LAYER met3 ;
      RECT -6.040000 -5.910000 7.540000  4.090000 ;
      RECT -6.040000 25.910000 7.540000 35.910000 ;
      RECT -4.840000  4.090000 6.340000 25.910000 ;
    LAYER via ;
      RECT -5.930000 -5.760000 -3.750000 35.780000 ;
      RECT -3.540000 -5.760000  5.040000 -3.580000 ;
      RECT -3.540000 33.600000  5.040000 35.780000 ;
      RECT -1.940000 -1.930000  3.440000 31.930000 ;
      RECT  5.250000 -5.760000  7.430000 35.780000 ;
    LAYER via2 ;
      RECT -1.985000 -1.940000 3.495000 31.940000 ;
  END
END sky130_fd_pr__esd_rf_nfet_20v0_hbm_32vW60p00
END LIBRARY
