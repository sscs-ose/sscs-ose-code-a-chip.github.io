# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  3.990000 BY  6.940000 ;
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 3.595000 4.060000 5.955000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.636000 ;
    PORT
      LAYER li1 ;
        RECT 1.190000 0.000000 2.940000 0.695000 ;
        RECT 1.190000 6.245000 2.940000 6.940000 ;
      LAYER mcon ;
        RECT 1.260000 0.095000 2.870000 0.625000 ;
        RECT 1.260000 6.315000 2.870000 6.845000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.180000 0.000000 2.950000 0.685000 ;
        RECT 1.180000 6.255000 2.950000 6.940000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 0.985000 4.060000 3.345000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  3.282500 ;
    ANTENNAGATEAREA  0.757500 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 0.985000 0.500000 5.955000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.630000 0.985000 3.925000 5.955000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 0.800000 6.015000 ;
      RECT 0.580000 0.485000 0.910000 0.815000 ;
      RECT 0.580000 0.815000 0.800000 0.925000 ;
      RECT 0.580000 6.015000 0.800000 6.125000 ;
      RECT 0.580000 6.125000 0.910000 6.455000 ;
      RECT 1.060000 0.925000 1.230000 6.015000 ;
      RECT 1.520000 0.925000 1.690000 6.015000 ;
      RECT 1.980000 0.925000 2.150000 6.015000 ;
      RECT 2.440000 0.925000 2.610000 6.015000 ;
      RECT 2.900000 0.925000 3.070000 6.015000 ;
      RECT 3.220000 0.485000 3.550000 0.815000 ;
      RECT 3.220000 6.125000 3.550000 6.455000 ;
      RECT 3.330000 0.815000 3.550000 0.925000 ;
      RECT 3.330000 0.925000 3.925000 6.015000 ;
      RECT 3.330000 6.015000 3.550000 6.125000 ;
    LAYER mcon ;
      RECT 0.300000 1.045000 0.470000 1.215000 ;
      RECT 0.300000 1.405000 0.470000 1.575000 ;
      RECT 0.300000 1.765000 0.470000 1.935000 ;
      RECT 0.300000 2.125000 0.470000 2.295000 ;
      RECT 0.300000 2.485000 0.470000 2.655000 ;
      RECT 0.300000 2.845000 0.470000 3.015000 ;
      RECT 0.300000 3.205000 0.470000 3.375000 ;
      RECT 0.300000 3.565000 0.470000 3.735000 ;
      RECT 0.300000 3.925000 0.470000 4.095000 ;
      RECT 0.300000 4.285000 0.470000 4.455000 ;
      RECT 0.300000 4.645000 0.470000 4.815000 ;
      RECT 0.300000 5.005000 0.470000 5.175000 ;
      RECT 0.300000 5.365000 0.470000 5.535000 ;
      RECT 0.300000 5.725000 0.470000 5.895000 ;
      RECT 1.060000 1.045000 1.230000 1.215000 ;
      RECT 1.060000 1.405000 1.230000 1.575000 ;
      RECT 1.060000 1.765000 1.230000 1.935000 ;
      RECT 1.060000 2.125000 1.230000 2.295000 ;
      RECT 1.060000 2.485000 1.230000 2.655000 ;
      RECT 1.060000 2.845000 1.230000 3.015000 ;
      RECT 1.060000 3.205000 1.230000 3.375000 ;
      RECT 1.060000 3.565000 1.230000 3.735000 ;
      RECT 1.060000 3.925000 1.230000 4.095000 ;
      RECT 1.060000 4.285000 1.230000 4.455000 ;
      RECT 1.060000 4.645000 1.230000 4.815000 ;
      RECT 1.060000 5.005000 1.230000 5.175000 ;
      RECT 1.060000 5.365000 1.230000 5.535000 ;
      RECT 1.060000 5.725000 1.230000 5.895000 ;
      RECT 1.520000 1.045000 1.690000 1.215000 ;
      RECT 1.520000 1.405000 1.690000 1.575000 ;
      RECT 1.520000 1.765000 1.690000 1.935000 ;
      RECT 1.520000 2.125000 1.690000 2.295000 ;
      RECT 1.520000 2.485000 1.690000 2.655000 ;
      RECT 1.520000 2.845000 1.690000 3.015000 ;
      RECT 1.520000 3.205000 1.690000 3.375000 ;
      RECT 1.520000 3.565000 1.690000 3.735000 ;
      RECT 1.520000 3.925000 1.690000 4.095000 ;
      RECT 1.520000 4.285000 1.690000 4.455000 ;
      RECT 1.520000 4.645000 1.690000 4.815000 ;
      RECT 1.520000 5.005000 1.690000 5.175000 ;
      RECT 1.520000 5.365000 1.690000 5.535000 ;
      RECT 1.520000 5.725000 1.690000 5.895000 ;
      RECT 1.980000 1.045000 2.150000 1.215000 ;
      RECT 1.980000 1.405000 2.150000 1.575000 ;
      RECT 1.980000 1.765000 2.150000 1.935000 ;
      RECT 1.980000 2.125000 2.150000 2.295000 ;
      RECT 1.980000 2.485000 2.150000 2.655000 ;
      RECT 1.980000 2.845000 2.150000 3.015000 ;
      RECT 1.980000 3.205000 2.150000 3.375000 ;
      RECT 1.980000 3.565000 2.150000 3.735000 ;
      RECT 1.980000 3.925000 2.150000 4.095000 ;
      RECT 1.980000 4.285000 2.150000 4.455000 ;
      RECT 1.980000 4.645000 2.150000 4.815000 ;
      RECT 1.980000 5.005000 2.150000 5.175000 ;
      RECT 1.980000 5.365000 2.150000 5.535000 ;
      RECT 1.980000 5.725000 2.150000 5.895000 ;
      RECT 2.440000 1.045000 2.610000 1.215000 ;
      RECT 2.440000 1.405000 2.610000 1.575000 ;
      RECT 2.440000 1.765000 2.610000 1.935000 ;
      RECT 2.440000 2.125000 2.610000 2.295000 ;
      RECT 2.440000 2.485000 2.610000 2.655000 ;
      RECT 2.440000 2.845000 2.610000 3.015000 ;
      RECT 2.440000 3.205000 2.610000 3.375000 ;
      RECT 2.440000 3.565000 2.610000 3.735000 ;
      RECT 2.440000 3.925000 2.610000 4.095000 ;
      RECT 2.440000 4.285000 2.610000 4.455000 ;
      RECT 2.440000 4.645000 2.610000 4.815000 ;
      RECT 2.440000 5.005000 2.610000 5.175000 ;
      RECT 2.440000 5.365000 2.610000 5.535000 ;
      RECT 2.440000 5.725000 2.610000 5.895000 ;
      RECT 2.900000 1.045000 3.070000 1.215000 ;
      RECT 2.900000 1.405000 3.070000 1.575000 ;
      RECT 2.900000 1.765000 3.070000 1.935000 ;
      RECT 2.900000 2.125000 3.070000 2.295000 ;
      RECT 2.900000 2.485000 3.070000 2.655000 ;
      RECT 2.900000 2.845000 3.070000 3.015000 ;
      RECT 2.900000 3.205000 3.070000 3.375000 ;
      RECT 2.900000 3.565000 3.070000 3.735000 ;
      RECT 2.900000 3.925000 3.070000 4.095000 ;
      RECT 2.900000 4.285000 3.070000 4.455000 ;
      RECT 2.900000 4.645000 3.070000 4.815000 ;
      RECT 2.900000 5.005000 3.070000 5.175000 ;
      RECT 2.900000 5.365000 3.070000 5.535000 ;
      RECT 2.900000 5.725000 3.070000 5.895000 ;
      RECT 3.660000 1.045000 3.830000 1.215000 ;
      RECT 3.660000 1.405000 3.830000 1.575000 ;
      RECT 3.660000 1.765000 3.830000 1.935000 ;
      RECT 3.660000 2.125000 3.830000 2.295000 ;
      RECT 3.660000 2.485000 3.830000 2.655000 ;
      RECT 3.660000 2.845000 3.830000 3.015000 ;
      RECT 3.660000 3.205000 3.830000 3.375000 ;
      RECT 3.660000 3.565000 3.830000 3.735000 ;
      RECT 3.660000 3.925000 3.830000 4.095000 ;
      RECT 3.660000 4.285000 3.830000 4.455000 ;
      RECT 3.660000 4.645000 3.830000 4.815000 ;
      RECT 3.660000 5.005000 3.830000 5.175000 ;
      RECT 3.660000 5.365000 3.830000 5.535000 ;
      RECT 3.660000 5.725000 3.830000 5.895000 ;
    LAYER met1 ;
      RECT 1.015000 0.985000 1.275000 5.955000 ;
      RECT 1.475000 0.985000 1.735000 5.955000 ;
      RECT 1.935000 0.985000 2.195000 5.955000 ;
      RECT 2.395000 0.985000 2.655000 5.955000 ;
      RECT 2.855000 0.985000 3.115000 5.955000 ;
    LAYER via ;
      RECT 1.015000 1.015000 1.275000 1.275000 ;
      RECT 1.015000 1.335000 1.275000 1.595000 ;
      RECT 1.015000 1.655000 1.275000 1.915000 ;
      RECT 1.015000 1.975000 1.275000 2.235000 ;
      RECT 1.015000 2.295000 1.275000 2.555000 ;
      RECT 1.015000 2.615000 1.275000 2.875000 ;
      RECT 1.015000 2.935000 1.275000 3.195000 ;
      RECT 1.475000 3.745000 1.735000 4.005000 ;
      RECT 1.475000 4.065000 1.735000 4.325000 ;
      RECT 1.475000 4.385000 1.735000 4.645000 ;
      RECT 1.475000 4.705000 1.735000 4.965000 ;
      RECT 1.475000 5.025000 1.735000 5.285000 ;
      RECT 1.475000 5.345000 1.735000 5.605000 ;
      RECT 1.475000 5.665000 1.735000 5.925000 ;
      RECT 1.935000 1.015000 2.195000 1.275000 ;
      RECT 1.935000 1.335000 2.195000 1.595000 ;
      RECT 1.935000 1.655000 2.195000 1.915000 ;
      RECT 1.935000 1.975000 2.195000 2.235000 ;
      RECT 1.935000 2.295000 2.195000 2.555000 ;
      RECT 1.935000 2.615000 2.195000 2.875000 ;
      RECT 1.935000 2.935000 2.195000 3.195000 ;
      RECT 2.395000 3.745000 2.655000 4.005000 ;
      RECT 2.395000 4.065000 2.655000 4.325000 ;
      RECT 2.395000 4.385000 2.655000 4.645000 ;
      RECT 2.395000 4.705000 2.655000 4.965000 ;
      RECT 2.395000 5.025000 2.655000 5.285000 ;
      RECT 2.395000 5.345000 2.655000 5.605000 ;
      RECT 2.395000 5.665000 2.655000 5.925000 ;
      RECT 2.855000 1.015000 3.115000 1.275000 ;
      RECT 2.855000 1.335000 3.115000 1.595000 ;
      RECT 2.855000 1.655000 3.115000 1.915000 ;
      RECT 2.855000 1.975000 3.115000 2.235000 ;
      RECT 2.855000 2.295000 3.115000 2.555000 ;
      RECT 2.855000 2.615000 3.115000 2.875000 ;
      RECT 2.855000 2.935000 3.115000 3.195000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18
END LIBRARY
