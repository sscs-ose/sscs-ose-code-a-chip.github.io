* SKY130 Spice File.
* Number of bins: 1
* 9 parameters
.param
+ sky130_fd_bs_flash__special_sonosfet_star__tox_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__overlap_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__lint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__wint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__dlc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__dwc_diff = 0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 000, W = 0.45, L = 0.22
* ------------------------------------
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0 = 9.2685e-1
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0 = -3.5390e-3
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0 = -4.3689e-1
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0 = 0.0
