# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.33000 BY  11.33000 ;
  PIN C0
    PORT
      LAYER met4 ;
        RECT  0.000000  0.000000 11.330000  0.330000 ;
        RECT  0.000000  0.330000  0.330000  1.230000 ;
        RECT  0.000000  1.230000  5.130000  1.530000 ;
        RECT  0.000000  1.530000  0.330000  2.430000 ;
        RECT  0.000000  2.430000  5.130000  2.730000 ;
        RECT  0.000000  2.730000  0.330000  3.630000 ;
        RECT  0.000000  3.630000  5.130000  3.930000 ;
        RECT  0.000000  3.930000  0.330000  4.830000 ;
        RECT  0.000000  4.830000  5.130000  5.130000 ;
        RECT  0.000000  5.130000  0.330000  6.200000 ;
        RECT  0.000000  6.200000  5.130000  6.500000 ;
        RECT  0.000000  6.500000  0.330000  7.400000 ;
        RECT  0.000000  7.400000  5.130000  7.700000 ;
        RECT  0.000000  7.700000  0.330000  8.600000 ;
        RECT  0.000000  8.600000  5.130000  8.900000 ;
        RECT  0.000000  8.900000  0.330000  9.800000 ;
        RECT  0.000000  9.800000  5.130000 10.100000 ;
        RECT  0.000000 10.100000  0.330000 11.000000 ;
        RECT  0.000000 11.000000 11.330000 11.330000 ;
        RECT  6.200000  1.230000 11.330000  1.530000 ;
        RECT  6.200000  2.430000 11.330000  2.730000 ;
        RECT  6.200000  3.630000 11.330000  3.930000 ;
        RECT  6.200000  4.830000 11.330000  5.130000 ;
        RECT  6.200000  6.200000 11.330000  6.500000 ;
        RECT  6.200000  7.400000 11.330000  7.700000 ;
        RECT  6.200000  8.600000 11.330000  8.900000 ;
        RECT  6.200000  9.800000 11.330000 10.100000 ;
        RECT 11.000000  0.330000 11.330000  1.230000 ;
        RECT 11.000000  1.530000 11.330000  2.430000 ;
        RECT 11.000000  2.730000 11.330000  3.630000 ;
        RECT 11.000000  3.930000 11.330000  4.830000 ;
        RECT 11.000000  5.130000 11.330000  6.200000 ;
        RECT 11.000000  6.500000 11.330000  7.400000 ;
        RECT 11.000000  7.700000 11.330000  8.600000 ;
        RECT 11.000000  8.900000 11.330000  9.800000 ;
        RECT 11.000000 10.100000 11.330000 11.000000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met4 ;
        RECT 0.630000  0.630000 10.700000  0.930000 ;
        RECT 0.630000  1.830000 10.700000  2.130000 ;
        RECT 0.630000  3.030000 10.700000  3.330000 ;
        RECT 0.630000  4.230000 10.700000  4.530000 ;
        RECT 0.630000  5.430000 10.700000  5.900000 ;
        RECT 0.630000  6.800000 10.700000  7.100000 ;
        RECT 0.630000  8.000000 10.700000  8.300000 ;
        RECT 0.630000  9.200000 10.700000  9.500000 ;
        RECT 0.630000 10.400000 10.700000 10.700000 ;
        RECT 5.430000  0.930000  5.900000  1.830000 ;
        RECT 5.430000  2.130000  5.900000  3.030000 ;
        RECT 5.430000  3.330000  5.900000  4.230000 ;
        RECT 5.430000  4.530000  5.900000  5.430000 ;
        RECT 5.430000  5.900000  5.900000  6.800000 ;
        RECT 5.430000  7.100000  5.900000  8.000000 ;
        RECT 5.430000  8.300000  5.900000  9.200000 ;
        RECT 5.430000  9.500000  5.900000 10.400000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 7.755000 8.735000 7.860000 8.980000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT  0.080000  0.080000 11.250000  0.250000 ;
      RECT  0.080000  0.250000  0.250000 11.080000 ;
      RECT  0.080000 11.080000 11.250000 11.250000 ;
      RECT 11.080000  0.250000 11.250000 11.080000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 11.330000  0.330000 ;
      RECT  0.000000  0.330000  0.330000 11.000000 ;
      RECT  0.000000 11.000000 11.330000 11.330000 ;
      RECT  0.470000  0.470000  0.610000  5.510000 ;
      RECT  0.470000  5.510000 10.860000  5.820000 ;
      RECT  0.470000  5.820000  0.610000 10.860000 ;
      RECT  0.750000  0.330000  0.890000  5.370000 ;
      RECT  0.750000  5.960000  0.890000 11.000000 ;
      RECT  1.030000  0.470000  1.170000  5.510000 ;
      RECT  1.030000  5.820000  1.170000 10.860000 ;
      RECT  1.310000  0.330000  1.450000  5.370000 ;
      RECT  1.310000  5.960000  1.450000 11.000000 ;
      RECT  1.590000  0.470000  1.730000  5.510000 ;
      RECT  1.590000  5.820000  1.730000 10.860000 ;
      RECT  1.870000  0.330000  2.010000  5.370000 ;
      RECT  1.870000  5.960000  2.010000 11.000000 ;
      RECT  2.150000  0.470000  2.290000  5.510000 ;
      RECT  2.150000  5.820000  2.290000 10.860000 ;
      RECT  2.430000  0.330000  2.570000  5.370000 ;
      RECT  2.430000  5.960000  2.570000 11.000000 ;
      RECT  2.710000  0.470000  2.850000  5.510000 ;
      RECT  2.710000  5.820000  2.850000 10.860000 ;
      RECT  2.990000  0.330000  3.130000  5.370000 ;
      RECT  2.990000  5.960000  3.130000 11.000000 ;
      RECT  3.270000  0.470000  3.410000  5.510000 ;
      RECT  3.270000  5.820000  3.410000 10.860000 ;
      RECT  3.550000  0.330000  3.690000  5.370000 ;
      RECT  3.550000  5.960000  3.690000 11.000000 ;
      RECT  3.830000  0.470000  3.970000  5.510000 ;
      RECT  3.830000  5.820000  3.970000 10.860000 ;
      RECT  4.110000  0.330000  4.250000  5.370000 ;
      RECT  4.110000  5.960000  4.250000 11.000000 ;
      RECT  4.390000  0.470000  4.530000  5.510000 ;
      RECT  4.390000  5.820000  4.530000 10.860000 ;
      RECT  4.670000  0.330000  4.810000  5.370000 ;
      RECT  4.670000  5.960000  4.810000 11.000000 ;
      RECT  4.950000  0.470000  5.090000  5.510000 ;
      RECT  4.950000  5.820000  5.090000 10.860000 ;
      RECT  5.230000  0.330000  5.370000  5.370000 ;
      RECT  5.230000  5.960000  5.370000 11.000000 ;
      RECT  5.510000  0.470000  5.820000  5.510000 ;
      RECT  5.510000  5.820000  5.820000 10.860000 ;
      RECT  5.960000  0.330000  6.100000  5.370000 ;
      RECT  5.960000  5.960000  6.100000 11.000000 ;
      RECT  6.240000  0.470000  6.380000  5.510000 ;
      RECT  6.240000  5.820000  6.380000 10.860000 ;
      RECT  6.520000  0.330000  6.660000  5.370000 ;
      RECT  6.520000  5.960000  6.660000 11.000000 ;
      RECT  6.800000  0.470000  6.940000  5.510000 ;
      RECT  6.800000  5.820000  6.940000 10.860000 ;
      RECT  7.080000  0.330000  7.220000  5.370000 ;
      RECT  7.080000  5.960000  7.220000 11.000000 ;
      RECT  7.360000  0.470000  7.500000  5.510000 ;
      RECT  7.360000  5.820000  7.500000 10.860000 ;
      RECT  7.640000  0.330000  7.780000  5.370000 ;
      RECT  7.640000  5.960000  7.780000 11.000000 ;
      RECT  7.920000  0.470000  8.060000  5.510000 ;
      RECT  7.920000  5.820000  8.060000 10.860000 ;
      RECT  8.200000  0.330000  8.340000  5.370000 ;
      RECT  8.200000  5.960000  8.340000 11.000000 ;
      RECT  8.480000  0.470000  8.620000  5.510000 ;
      RECT  8.480000  5.820000  8.620000 10.860000 ;
      RECT  8.760000  0.330000  8.900000  5.370000 ;
      RECT  8.760000  5.960000  8.900000 11.000000 ;
      RECT  9.040000  0.470000  9.180000  5.510000 ;
      RECT  9.040000  5.820000  9.180000 10.860000 ;
      RECT  9.320000  0.330000  9.460000  5.370000 ;
      RECT  9.320000  5.960000  9.460000 11.000000 ;
      RECT  9.600000  0.470000  9.740000  5.510000 ;
      RECT  9.600000  5.820000  9.740000 10.860000 ;
      RECT  9.880000  0.330000 10.020000  5.370000 ;
      RECT  9.880000  5.960000 10.020000 11.000000 ;
      RECT 10.160000  0.470000 10.300000  5.510000 ;
      RECT 10.160000  5.820000 10.300000 10.860000 ;
      RECT 10.440000  0.330000 10.580000  5.370000 ;
      RECT 10.440000  5.960000 10.580000 11.000000 ;
      RECT 10.720000  0.470000 10.860000  5.510000 ;
      RECT 10.720000  5.820000 10.860000 10.860000 ;
      RECT 11.000000  0.330000 11.330000 11.000000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  5.370000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.750000 ;
      RECT  0.000000  0.750000  5.370000  0.890000 ;
      RECT  0.000000  0.890000  0.330000  1.310000 ;
      RECT  0.000000  1.310000  5.370000  1.450000 ;
      RECT  0.000000  1.450000  0.330000  1.870000 ;
      RECT  0.000000  1.870000  5.370000  2.010000 ;
      RECT  0.000000  2.010000  0.330000  2.430000 ;
      RECT  0.000000  2.430000  5.370000  2.570000 ;
      RECT  0.000000  2.570000  0.330000  2.990000 ;
      RECT  0.000000  2.990000  5.370000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.550000 ;
      RECT  0.000000  3.550000  5.370000  3.690000 ;
      RECT  0.000000  3.690000  0.330000  4.110000 ;
      RECT  0.000000  4.110000  5.370000  4.250000 ;
      RECT  0.000000  4.250000  0.330000  4.670000 ;
      RECT  0.000000  4.670000  5.370000  4.810000 ;
      RECT  0.000000  4.810000  0.330000  5.230000 ;
      RECT  0.000000  5.230000  5.370000  5.370000 ;
      RECT  0.000000  5.960000  5.370000  6.100000 ;
      RECT  0.000000  6.100000  0.330000  6.520000 ;
      RECT  0.000000  6.520000  5.370000  6.660000 ;
      RECT  0.000000  6.660000  0.330000  7.080000 ;
      RECT  0.000000  7.080000  5.370000  7.220000 ;
      RECT  0.000000  7.220000  0.330000  7.640000 ;
      RECT  0.000000  7.640000  5.370000  7.780000 ;
      RECT  0.000000  7.780000  0.330000  8.200000 ;
      RECT  0.000000  8.200000  5.370000  8.340000 ;
      RECT  0.000000  8.340000  0.330000  8.760000 ;
      RECT  0.000000  8.760000  5.370000  8.900000 ;
      RECT  0.000000  8.900000  0.330000  9.320000 ;
      RECT  0.000000  9.320000  5.370000  9.460000 ;
      RECT  0.000000  9.460000  0.330000  9.880000 ;
      RECT  0.000000  9.880000  5.370000 10.020000 ;
      RECT  0.000000 10.020000  0.330000 10.440000 ;
      RECT  0.000000 10.440000  5.370000 10.580000 ;
      RECT  0.000000 10.580000  0.330000 11.000000 ;
      RECT  0.000000 11.000000  5.370000 11.330000 ;
      RECT  0.330000  5.510000 11.000000  5.820000 ;
      RECT  0.470000  0.470000 10.860000  0.610000 ;
      RECT  0.470000  1.030000 10.860000  1.170000 ;
      RECT  0.470000  1.590000 10.860000  1.730000 ;
      RECT  0.470000  2.150000 10.860000  2.290000 ;
      RECT  0.470000  2.710000 10.860000  2.850000 ;
      RECT  0.470000  3.270000 10.860000  3.410000 ;
      RECT  0.470000  3.830000 10.860000  3.970000 ;
      RECT  0.470000  4.390000 10.860000  4.530000 ;
      RECT  0.470000  4.950000 10.860000  5.090000 ;
      RECT  0.470000  6.240000 10.860000  6.380000 ;
      RECT  0.470000  6.800000 10.860000  6.940000 ;
      RECT  0.470000  7.360000 10.860000  7.500000 ;
      RECT  0.470000  7.920000 10.860000  8.060000 ;
      RECT  0.470000  8.480000 10.860000  8.620000 ;
      RECT  0.470000  9.040000 10.860000  9.180000 ;
      RECT  0.470000  9.600000 10.860000  9.740000 ;
      RECT  0.470000 10.160000 10.860000 10.300000 ;
      RECT  0.470000 10.720000 10.860000 10.860000 ;
      RECT  5.510000  0.330000  5.820000  0.470000 ;
      RECT  5.510000  0.610000  5.820000  1.030000 ;
      RECT  5.510000  1.170000  5.820000  1.590000 ;
      RECT  5.510000  1.730000  5.820000  2.150000 ;
      RECT  5.510000  2.290000  5.820000  2.710000 ;
      RECT  5.510000  2.850000  5.820000  3.270000 ;
      RECT  5.510000  3.410000  5.820000  3.830000 ;
      RECT  5.510000  3.970000  5.820000  4.390000 ;
      RECT  5.510000  4.530000  5.820000  4.950000 ;
      RECT  5.510000  5.090000  5.820000  5.510000 ;
      RECT  5.510000  5.820000  5.820000  6.240000 ;
      RECT  5.510000  6.380000  5.820000  6.800000 ;
      RECT  5.510000  6.940000  5.820000  7.360000 ;
      RECT  5.510000  7.500000  5.820000  7.920000 ;
      RECT  5.510000  8.060000  5.820000  8.480000 ;
      RECT  5.510000  8.620000  5.820000  9.040000 ;
      RECT  5.510000  9.180000  5.820000  9.600000 ;
      RECT  5.510000  9.740000  5.820000 10.160000 ;
      RECT  5.510000 10.300000  5.820000 10.720000 ;
      RECT  5.510000 10.860000  5.820000 11.000000 ;
      RECT  5.960000  0.000000 11.330000  0.330000 ;
      RECT  5.960000  0.750000 11.330000  0.890000 ;
      RECT  5.960000  1.310000 11.330000  1.450000 ;
      RECT  5.960000  1.870000 11.330000  2.010000 ;
      RECT  5.960000  2.430000 11.330000  2.570000 ;
      RECT  5.960000  2.990000 11.330000  3.130000 ;
      RECT  5.960000  3.550000 11.330000  3.690000 ;
      RECT  5.960000  4.110000 11.330000  4.250000 ;
      RECT  5.960000  4.670000 11.330000  4.810000 ;
      RECT  5.960000  5.230000 11.330000  5.370000 ;
      RECT  5.960000  5.960000 11.330000  6.100000 ;
      RECT  5.960000  6.520000 11.330000  6.660000 ;
      RECT  5.960000  7.080000 11.330000  7.220000 ;
      RECT  5.960000  7.640000 11.330000  7.780000 ;
      RECT  5.960000  8.200000 11.330000  8.340000 ;
      RECT  5.960000  8.760000 11.330000  8.900000 ;
      RECT  5.960000  9.320000 11.330000  9.460000 ;
      RECT  5.960000  9.880000 11.330000 10.020000 ;
      RECT  5.960000 10.440000 11.330000 10.580000 ;
      RECT  5.960000 11.000000 11.330000 11.330000 ;
      RECT 11.000000  0.330000 11.330000  0.750000 ;
      RECT 11.000000  0.890000 11.330000  1.310000 ;
      RECT 11.000000  1.450000 11.330000  1.870000 ;
      RECT 11.000000  2.010000 11.330000  2.430000 ;
      RECT 11.000000  2.570000 11.330000  2.990000 ;
      RECT 11.000000  3.130000 11.330000  3.550000 ;
      RECT 11.000000  3.690000 11.330000  4.110000 ;
      RECT 11.000000  4.250000 11.330000  4.670000 ;
      RECT 11.000000  4.810000 11.330000  5.230000 ;
      RECT 11.000000  6.100000 11.330000  6.520000 ;
      RECT 11.000000  6.660000 11.330000  7.080000 ;
      RECT 11.000000  7.220000 11.330000  7.640000 ;
      RECT 11.000000  7.780000 11.330000  8.200000 ;
      RECT 11.000000  8.340000 11.330000  8.760000 ;
      RECT 11.000000  8.900000 11.330000  9.320000 ;
      RECT 11.000000  9.460000 11.330000  9.880000 ;
      RECT 11.000000 10.020000 11.330000 10.440000 ;
      RECT 11.000000 10.580000 11.330000 11.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000  5.130000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  5.130000 ;
      RECT  0.000000  6.200000  0.330000 11.000000 ;
      RECT  0.000000 11.000000  5.130000 11.330000 ;
      RECT  0.330000  5.430000 11.000000  5.900000 ;
      RECT  0.630000  0.630000  0.930000  5.430000 ;
      RECT  0.630000  5.900000  0.930000 10.700000 ;
      RECT  1.230000  0.330000  1.530000  5.130000 ;
      RECT  1.230000  6.200000  1.530000 11.000000 ;
      RECT  1.830000  0.630000  2.130000  5.430000 ;
      RECT  1.830000  5.900000  2.130000 10.700000 ;
      RECT  2.430000  0.330000  2.730000  5.130000 ;
      RECT  2.430000  6.200000  2.730000 11.000000 ;
      RECT  3.030000  0.630000  3.330000  5.430000 ;
      RECT  3.030000  5.900000  3.330000 10.700000 ;
      RECT  3.630000  0.330000  3.930000  5.130000 ;
      RECT  3.630000  6.200000  3.930000 11.000000 ;
      RECT  4.230000  0.630000  4.530000  5.430000 ;
      RECT  4.230000  5.900000  4.530000 10.700000 ;
      RECT  4.830000  0.330000  5.130000  5.130000 ;
      RECT  4.830000  6.200000  5.130000 11.000000 ;
      RECT  5.430000  0.330000  5.900000  5.430000 ;
      RECT  5.430000  5.900000  5.900000 11.000000 ;
      RECT  6.200000  0.000000 11.330000  0.330000 ;
      RECT  6.200000  0.330000  6.500000  5.130000 ;
      RECT  6.200000  6.200000  6.500000 11.000000 ;
      RECT  6.200000 11.000000 11.330000 11.330000 ;
      RECT  6.800000  0.630000  7.100000  5.430000 ;
      RECT  6.800000  5.900000  7.100000 10.700000 ;
      RECT  7.400000  0.330000  7.700000  5.130000 ;
      RECT  7.400000  6.200000  7.700000 11.000000 ;
      RECT  8.000000  0.630000  8.300000  5.430000 ;
      RECT  8.000000  5.900000  8.300000 10.700000 ;
      RECT  8.600000  0.330000  8.900000  5.130000 ;
      RECT  8.600000  6.200000  8.900000 11.000000 ;
      RECT  9.200000  0.630000  9.500000  5.430000 ;
      RECT  9.200000  5.900000  9.500000 10.700000 ;
      RECT  9.800000  0.330000 10.100000  5.130000 ;
      RECT  9.800000  6.200000 10.100000 11.000000 ;
      RECT 10.400000  0.630000 10.700000  5.430000 ;
      RECT 10.400000  5.900000 10.700000 10.700000 ;
      RECT 11.000000  0.330000 11.330000  5.130000 ;
      RECT 11.000000  6.200000 11.330000 11.000000 ;
    LAYER via ;
      RECT  0.035000  0.680000  0.295000  0.940000 ;
      RECT  0.035000  1.080000  0.295000  1.340000 ;
      RECT  0.035000  1.480000  0.295000  1.740000 ;
      RECT  0.035000  1.880000  0.295000  2.140000 ;
      RECT  0.035000  2.280000  0.295000  2.540000 ;
      RECT  0.035000  2.680000  0.295000  2.940000 ;
      RECT  0.035000  3.080000  0.295000  3.340000 ;
      RECT  0.035000  3.480000  0.295000  3.740000 ;
      RECT  0.035000  3.880000  0.295000  4.140000 ;
      RECT  0.035000  4.280000  0.295000  4.540000 ;
      RECT  0.035000  4.680000  0.295000  4.940000 ;
      RECT  0.035000  5.080000  0.295000  5.340000 ;
      RECT  0.035000  5.990000  0.295000  6.250000 ;
      RECT  0.035000  6.390000  0.295000  6.650000 ;
      RECT  0.035000  6.790000  0.295000  7.050000 ;
      RECT  0.035000  7.190000  0.295000  7.450000 ;
      RECT  0.035000  7.590000  0.295000  7.850000 ;
      RECT  0.035000  7.990000  0.295000  8.250000 ;
      RECT  0.035000  8.390000  0.295000  8.650000 ;
      RECT  0.035000  8.790000  0.295000  9.050000 ;
      RECT  0.035000  9.190000  0.295000  9.450000 ;
      RECT  0.035000  9.590000  0.295000  9.850000 ;
      RECT  0.035000  9.990000  0.295000 10.250000 ;
      RECT  0.035000 10.390000  0.295000 10.650000 ;
      RECT  0.280000  0.035000  0.540000  0.295000 ;
      RECT  0.280000 11.035000  0.540000 11.295000 ;
      RECT  0.680000  0.035000  0.940000  0.295000 ;
      RECT  0.680000 11.035000  0.940000 11.295000 ;
      RECT  0.735000  5.535000  0.995000  5.795000 ;
      RECT  1.080000  0.035000  1.340000  0.295000 ;
      RECT  1.080000 11.035000  1.340000 11.295000 ;
      RECT  1.135000  5.535000  1.395000  5.795000 ;
      RECT  1.480000  0.035000  1.740000  0.295000 ;
      RECT  1.480000 11.035000  1.740000 11.295000 ;
      RECT  1.535000  5.535000  1.795000  5.795000 ;
      RECT  1.880000  0.035000  2.140000  0.295000 ;
      RECT  1.880000 11.035000  2.140000 11.295000 ;
      RECT  1.935000  5.535000  2.195000  5.795000 ;
      RECT  2.280000  0.035000  2.540000  0.295000 ;
      RECT  2.280000 11.035000  2.540000 11.295000 ;
      RECT  2.335000  5.535000  2.595000  5.795000 ;
      RECT  2.680000  0.035000  2.940000  0.295000 ;
      RECT  2.680000 11.035000  2.940000 11.295000 ;
      RECT  2.735000  5.535000  2.995000  5.795000 ;
      RECT  3.080000  0.035000  3.340000  0.295000 ;
      RECT  3.080000 11.035000  3.340000 11.295000 ;
      RECT  3.135000  5.535000  3.395000  5.795000 ;
      RECT  3.480000  0.035000  3.740000  0.295000 ;
      RECT  3.480000 11.035000  3.740000 11.295000 ;
      RECT  3.535000  5.535000  3.795000  5.795000 ;
      RECT  3.880000  0.035000  4.140000  0.295000 ;
      RECT  3.880000 11.035000  4.140000 11.295000 ;
      RECT  3.935000  5.535000  4.195000  5.795000 ;
      RECT  4.280000  0.035000  4.540000  0.295000 ;
      RECT  4.280000 11.035000  4.540000 11.295000 ;
      RECT  4.335000  5.535000  4.595000  5.795000 ;
      RECT  4.680000  0.035000  4.940000  0.295000 ;
      RECT  4.680000 11.035000  4.940000 11.295000 ;
      RECT  4.735000  5.535000  4.995000  5.795000 ;
      RECT  5.080000  0.035000  5.340000  0.295000 ;
      RECT  5.080000 11.035000  5.340000 11.295000 ;
      RECT  5.135000  5.535000  5.395000  5.795000 ;
      RECT  5.535000  0.735000  5.795000  0.995000 ;
      RECT  5.535000  1.135000  5.795000  1.395000 ;
      RECT  5.535000  1.535000  5.795000  1.795000 ;
      RECT  5.535000  1.935000  5.795000  2.195000 ;
      RECT  5.535000  2.335000  5.795000  2.595000 ;
      RECT  5.535000  2.735000  5.795000  2.995000 ;
      RECT  5.535000  3.135000  5.795000  3.395000 ;
      RECT  5.535000  3.535000  5.795000  3.795000 ;
      RECT  5.535000  3.935000  5.795000  4.195000 ;
      RECT  5.535000  4.335000  5.795000  4.595000 ;
      RECT  5.535000  4.735000  5.795000  4.995000 ;
      RECT  5.535000  5.135000  5.795000  5.395000 ;
      RECT  5.535000  5.535000  5.795000  5.795000 ;
      RECT  5.535000  5.935000  5.795000  6.195000 ;
      RECT  5.535000  6.335000  5.795000  6.595000 ;
      RECT  5.535000  6.735000  5.795000  6.995000 ;
      RECT  5.535000  7.135000  5.795000  7.395000 ;
      RECT  5.535000  7.535000  5.795000  7.795000 ;
      RECT  5.535000  7.935000  5.795000  8.195000 ;
      RECT  5.535000  8.335000  5.795000  8.595000 ;
      RECT  5.535000  8.735000  5.795000  8.995000 ;
      RECT  5.535000  9.135000  5.795000  9.395000 ;
      RECT  5.535000  9.535000  5.795000  9.795000 ;
      RECT  5.535000  9.935000  5.795000 10.195000 ;
      RECT  5.535000 10.335000  5.795000 10.595000 ;
      RECT  5.935000  5.535000  6.195000  5.795000 ;
      RECT  5.990000  0.035000  6.250000  0.295000 ;
      RECT  5.990000 11.035000  6.250000 11.295000 ;
      RECT  6.335000  5.535000  6.595000  5.795000 ;
      RECT  6.390000  0.035000  6.650000  0.295000 ;
      RECT  6.390000 11.035000  6.650000 11.295000 ;
      RECT  6.735000  5.535000  6.995000  5.795000 ;
      RECT  6.790000  0.035000  7.050000  0.295000 ;
      RECT  6.790000 11.035000  7.050000 11.295000 ;
      RECT  7.135000  5.535000  7.395000  5.795000 ;
      RECT  7.190000  0.035000  7.450000  0.295000 ;
      RECT  7.190000 11.035000  7.450000 11.295000 ;
      RECT  7.535000  5.535000  7.795000  5.795000 ;
      RECT  7.590000  0.035000  7.850000  0.295000 ;
      RECT  7.590000 11.035000  7.850000 11.295000 ;
      RECT  7.935000  5.535000  8.195000  5.795000 ;
      RECT  7.990000  0.035000  8.250000  0.295000 ;
      RECT  7.990000 11.035000  8.250000 11.295000 ;
      RECT  8.335000  5.535000  8.595000  5.795000 ;
      RECT  8.390000  0.035000  8.650000  0.295000 ;
      RECT  8.390000 11.035000  8.650000 11.295000 ;
      RECT  8.735000  5.535000  8.995000  5.795000 ;
      RECT  8.790000  0.035000  9.050000  0.295000 ;
      RECT  8.790000 11.035000  9.050000 11.295000 ;
      RECT  9.135000  5.535000  9.395000  5.795000 ;
      RECT  9.190000  0.035000  9.450000  0.295000 ;
      RECT  9.190000 11.035000  9.450000 11.295000 ;
      RECT  9.535000  5.535000  9.795000  5.795000 ;
      RECT  9.590000  0.035000  9.850000  0.295000 ;
      RECT  9.590000 11.035000  9.850000 11.295000 ;
      RECT  9.935000  5.535000 10.195000  5.795000 ;
      RECT  9.990000  0.035000 10.250000  0.295000 ;
      RECT  9.990000 11.035000 10.250000 11.295000 ;
      RECT 10.335000  5.535000 10.595000  5.795000 ;
      RECT 10.390000  0.035000 10.650000  0.295000 ;
      RECT 10.390000 11.035000 10.650000 11.295000 ;
      RECT 10.790000  0.035000 11.050000  0.295000 ;
      RECT 10.790000 11.035000 11.050000 11.295000 ;
      RECT 11.035000  0.680000 11.295000  0.940000 ;
      RECT 11.035000  1.080000 11.295000  1.340000 ;
      RECT 11.035000  1.480000 11.295000  1.740000 ;
      RECT 11.035000  1.880000 11.295000  2.140000 ;
      RECT 11.035000  2.280000 11.295000  2.540000 ;
      RECT 11.035000  2.680000 11.295000  2.940000 ;
      RECT 11.035000  3.080000 11.295000  3.340000 ;
      RECT 11.035000  3.480000 11.295000  3.740000 ;
      RECT 11.035000  3.880000 11.295000  4.140000 ;
      RECT 11.035000  4.280000 11.295000  4.540000 ;
      RECT 11.035000  4.680000 11.295000  4.940000 ;
      RECT 11.035000  5.080000 11.295000  5.340000 ;
      RECT 11.035000  5.990000 11.295000  6.250000 ;
      RECT 11.035000  6.390000 11.295000  6.650000 ;
      RECT 11.035000  6.790000 11.295000  7.050000 ;
      RECT 11.035000  7.190000 11.295000  7.450000 ;
      RECT 11.035000  7.590000 11.295000  7.850000 ;
      RECT 11.035000  7.990000 11.295000  8.250000 ;
      RECT 11.035000  8.390000 11.295000  8.650000 ;
      RECT 11.035000  8.790000 11.295000  9.050000 ;
      RECT 11.035000  9.190000 11.295000  9.450000 ;
      RECT 11.035000  9.590000 11.295000  9.850000 ;
      RECT 11.035000  9.990000 11.295000 10.250000 ;
      RECT 11.035000 10.390000 11.295000 10.650000 ;
    LAYER via2 ;
      RECT  0.025000  0.390000  0.305000  0.670000 ;
      RECT  0.025000  1.020000  0.305000  1.300000 ;
      RECT  0.025000  1.650000  0.305000  1.930000 ;
      RECT  0.025000  2.280000  0.305000  2.560000 ;
      RECT  0.025000  2.910000  0.305000  3.190000 ;
      RECT  0.025000  3.540000  0.305000  3.820000 ;
      RECT  0.025000  4.170000  0.305000  4.450000 ;
      RECT  0.025000  4.800000  0.305000  5.080000 ;
      RECT  0.025000  6.250000  0.305000  6.530000 ;
      RECT  0.025000  6.880000  0.305000  7.160000 ;
      RECT  0.025000  7.510000  0.305000  7.790000 ;
      RECT  0.025000  8.140000  0.305000  8.420000 ;
      RECT  0.025000  8.770000  0.305000  9.050000 ;
      RECT  0.025000  9.400000  0.305000  9.680000 ;
      RECT  0.025000 10.030000  0.305000 10.310000 ;
      RECT  0.025000 10.660000  0.305000 10.940000 ;
      RECT  0.390000  0.025000  0.670000  0.305000 ;
      RECT  0.390000 11.025000  0.670000 11.305000 ;
      RECT  0.485000  5.525000  0.765000  5.805000 ;
      RECT  1.020000  0.025000  1.300000  0.305000 ;
      RECT  1.020000 11.025000  1.300000 11.305000 ;
      RECT  1.115000  5.525000  1.395000  5.805000 ;
      RECT  1.650000  0.025000  1.930000  0.305000 ;
      RECT  1.650000 11.025000  1.930000 11.305000 ;
      RECT  1.745000  5.525000  2.025000  5.805000 ;
      RECT  2.280000  0.025000  2.560000  0.305000 ;
      RECT  2.280000 11.025000  2.560000 11.305000 ;
      RECT  2.375000  5.525000  2.655000  5.805000 ;
      RECT  2.910000  0.025000  3.190000  0.305000 ;
      RECT  2.910000 11.025000  3.190000 11.305000 ;
      RECT  3.005000  5.525000  3.285000  5.805000 ;
      RECT  3.540000  0.025000  3.820000  0.305000 ;
      RECT  3.540000 11.025000  3.820000 11.305000 ;
      RECT  3.635000  5.525000  3.915000  5.805000 ;
      RECT  4.170000  0.025000  4.450000  0.305000 ;
      RECT  4.170000 11.025000  4.450000 11.305000 ;
      RECT  4.265000  5.525000  4.545000  5.805000 ;
      RECT  4.800000  0.025000  5.080000  0.305000 ;
      RECT  4.800000 11.025000  5.080000 11.305000 ;
      RECT  4.895000  5.525000  5.175000  5.805000 ;
      RECT  5.525000  0.485000  5.805000  0.765000 ;
      RECT  5.525000  1.115000  5.805000  1.395000 ;
      RECT  5.525000  1.745000  5.805000  2.025000 ;
      RECT  5.525000  2.375000  5.805000  2.655000 ;
      RECT  5.525000  3.005000  5.805000  3.285000 ;
      RECT  5.525000  3.635000  5.805000  3.915000 ;
      RECT  5.525000  4.265000  5.805000  4.545000 ;
      RECT  5.525000  4.895000  5.805000  5.175000 ;
      RECT  5.525000  5.525000  5.805000  5.805000 ;
      RECT  5.525000  6.155000  5.805000  6.435000 ;
      RECT  5.525000  6.785000  5.805000  7.065000 ;
      RECT  5.525000  7.415000  5.805000  7.695000 ;
      RECT  5.525000  8.045000  5.805000  8.325000 ;
      RECT  5.525000  8.675000  5.805000  8.955000 ;
      RECT  5.525000  9.305000  5.805000  9.585000 ;
      RECT  5.525000  9.935000  5.805000 10.215000 ;
      RECT  5.525000 10.565000  5.805000 10.845000 ;
      RECT  6.155000  5.525000  6.435000  5.805000 ;
      RECT  6.250000  0.025000  6.530000  0.305000 ;
      RECT  6.250000 11.025000  6.530000 11.305000 ;
      RECT  6.785000  5.525000  7.065000  5.805000 ;
      RECT  6.880000  0.025000  7.160000  0.305000 ;
      RECT  6.880000 11.025000  7.160000 11.305000 ;
      RECT  7.415000  5.525000  7.695000  5.805000 ;
      RECT  7.510000  0.025000  7.790000  0.305000 ;
      RECT  7.510000 11.025000  7.790000 11.305000 ;
      RECT  8.045000  5.525000  8.325000  5.805000 ;
      RECT  8.140000  0.025000  8.420000  0.305000 ;
      RECT  8.140000 11.025000  8.420000 11.305000 ;
      RECT  8.675000  5.525000  8.955000  5.805000 ;
      RECT  8.770000  0.025000  9.050000  0.305000 ;
      RECT  8.770000 11.025000  9.050000 11.305000 ;
      RECT  9.305000  5.525000  9.585000  5.805000 ;
      RECT  9.400000  0.025000  9.680000  0.305000 ;
      RECT  9.400000 11.025000  9.680000 11.305000 ;
      RECT  9.935000  5.525000 10.215000  5.805000 ;
      RECT 10.030000  0.025000 10.310000  0.305000 ;
      RECT 10.030000 11.025000 10.310000 11.305000 ;
      RECT 10.565000  5.525000 10.845000  5.805000 ;
      RECT 10.660000  0.025000 10.940000  0.305000 ;
      RECT 10.660000 11.025000 10.940000 11.305000 ;
      RECT 11.025000  0.390000 11.305000  0.670000 ;
      RECT 11.025000  1.020000 11.305000  1.300000 ;
      RECT 11.025000  1.650000 11.305000  1.930000 ;
      RECT 11.025000  2.280000 11.305000  2.560000 ;
      RECT 11.025000  2.910000 11.305000  3.190000 ;
      RECT 11.025000  3.540000 11.305000  3.820000 ;
      RECT 11.025000  4.170000 11.305000  4.450000 ;
      RECT 11.025000  4.800000 11.305000  5.080000 ;
      RECT 11.025000  6.250000 11.305000  6.530000 ;
      RECT 11.025000  6.880000 11.305000  7.160000 ;
      RECT 11.025000  7.510000 11.305000  7.790000 ;
      RECT 11.025000  8.140000 11.305000  8.420000 ;
      RECT 11.025000  8.770000 11.305000  9.050000 ;
      RECT 11.025000  9.400000 11.305000  9.680000 ;
      RECT 11.025000 10.030000 11.305000 10.310000 ;
      RECT 11.025000 10.660000 11.305000 10.940000 ;
    LAYER via3 ;
      RECT  0.005000  0.370000  0.325000  0.690000 ;
      RECT  0.005000  1.000000  0.325000  1.320000 ;
      RECT  0.005000  1.630000  0.325000  1.950000 ;
      RECT  0.005000  2.260000  0.325000  2.580000 ;
      RECT  0.005000  2.890000  0.325000  3.210000 ;
      RECT  0.005000  3.520000  0.325000  3.840000 ;
      RECT  0.005000  4.150000  0.325000  4.470000 ;
      RECT  0.005000  4.780000  0.325000  5.100000 ;
      RECT  0.005000  6.230000  0.325000  6.550000 ;
      RECT  0.005000  6.860000  0.325000  7.180000 ;
      RECT  0.005000  7.490000  0.325000  7.810000 ;
      RECT  0.005000  8.120000  0.325000  8.440000 ;
      RECT  0.005000  8.750000  0.325000  9.070000 ;
      RECT  0.005000  9.380000  0.325000  9.700000 ;
      RECT  0.005000 10.010000  0.325000 10.330000 ;
      RECT  0.005000 10.640000  0.325000 10.960000 ;
      RECT  0.370000  0.005000  0.690000  0.325000 ;
      RECT  0.370000 11.005000  0.690000 11.325000 ;
      RECT  1.000000  0.005000  1.320000  0.325000 ;
      RECT  1.000000 11.005000  1.320000 11.325000 ;
      RECT  1.095000  5.505000  1.415000  5.825000 ;
      RECT  1.630000  0.005000  1.950000  0.325000 ;
      RECT  1.630000 11.005000  1.950000 11.325000 ;
      RECT  1.725000  5.505000  2.045000  5.825000 ;
      RECT  2.260000  0.005000  2.580000  0.325000 ;
      RECT  2.260000 11.005000  2.580000 11.325000 ;
      RECT  2.355000  5.505000  2.675000  5.825000 ;
      RECT  2.890000  0.005000  3.210000  0.325000 ;
      RECT  2.890000 11.005000  3.210000 11.325000 ;
      RECT  2.985000  5.505000  3.305000  5.825000 ;
      RECT  3.520000  0.005000  3.840000  0.325000 ;
      RECT  3.520000 11.005000  3.840000 11.325000 ;
      RECT  3.615000  5.505000  3.935000  5.825000 ;
      RECT  4.150000  0.005000  4.470000  0.325000 ;
      RECT  4.150000 11.005000  4.470000 11.325000 ;
      RECT  4.245000  5.505000  4.565000  5.825000 ;
      RECT  4.780000  0.005000  5.100000  0.325000 ;
      RECT  4.780000 11.005000  5.100000 11.325000 ;
      RECT  4.875000  5.505000  5.195000  5.825000 ;
      RECT  5.505000  1.095000  5.825000  1.415000 ;
      RECT  5.505000  1.725000  5.825000  2.045000 ;
      RECT  5.505000  2.355000  5.825000  2.675000 ;
      RECT  5.505000  2.985000  5.825000  3.305000 ;
      RECT  5.505000  3.615000  5.825000  3.935000 ;
      RECT  5.505000  4.245000  5.825000  4.565000 ;
      RECT  5.505000  4.875000  5.825000  5.195000 ;
      RECT  5.505000  5.505000  5.825000  5.825000 ;
      RECT  5.505000  6.135000  5.825000  6.455000 ;
      RECT  5.505000  6.765000  5.825000  7.085000 ;
      RECT  5.505000  7.395000  5.825000  7.715000 ;
      RECT  5.505000  8.025000  5.825000  8.345000 ;
      RECT  5.505000  8.655000  5.825000  8.975000 ;
      RECT  5.505000  9.285000  5.825000  9.605000 ;
      RECT  5.505000  9.915000  5.825000 10.235000 ;
      RECT  6.135000  5.505000  6.455000  5.825000 ;
      RECT  6.230000  0.005000  6.550000  0.325000 ;
      RECT  6.230000 11.005000  6.550000 11.325000 ;
      RECT  6.765000  5.505000  7.085000  5.825000 ;
      RECT  6.860000  0.005000  7.180000  0.325000 ;
      RECT  6.860000 11.005000  7.180000 11.325000 ;
      RECT  7.395000  5.505000  7.715000  5.825000 ;
      RECT  7.490000  0.005000  7.810000  0.325000 ;
      RECT  7.490000 11.005000  7.810000 11.325000 ;
      RECT  8.025000  5.505000  8.345000  5.825000 ;
      RECT  8.120000  0.005000  8.440000  0.325000 ;
      RECT  8.120000 11.005000  8.440000 11.325000 ;
      RECT  8.655000  5.505000  8.975000  5.825000 ;
      RECT  8.750000  0.005000  9.070000  0.325000 ;
      RECT  8.750000 11.005000  9.070000 11.325000 ;
      RECT  9.285000  5.505000  9.605000  5.825000 ;
      RECT  9.380000  0.005000  9.700000  0.325000 ;
      RECT  9.380000 11.005000  9.700000 11.325000 ;
      RECT  9.915000  5.505000 10.235000  5.825000 ;
      RECT 10.010000  0.005000 10.330000  0.325000 ;
      RECT 10.010000 11.005000 10.330000 11.325000 ;
      RECT 10.640000  0.005000 10.960000  0.325000 ;
      RECT 10.640000 11.005000 10.960000 11.325000 ;
      RECT 11.005000  0.370000 11.325000  0.690000 ;
      RECT 11.005000  1.000000 11.325000  1.320000 ;
      RECT 11.005000  1.630000 11.325000  1.950000 ;
      RECT 11.005000  2.260000 11.325000  2.580000 ;
      RECT 11.005000  2.890000 11.325000  3.210000 ;
      RECT 11.005000  3.520000 11.325000  3.840000 ;
      RECT 11.005000  4.150000 11.325000  4.470000 ;
      RECT 11.005000  4.780000 11.325000  5.100000 ;
      RECT 11.005000  6.230000 11.325000  6.550000 ;
      RECT 11.005000  6.860000 11.325000  7.180000 ;
      RECT 11.005000  7.490000 11.325000  7.810000 ;
      RECT 11.005000  8.120000 11.325000  8.440000 ;
      RECT 11.005000  8.750000 11.325000  9.070000 ;
      RECT 11.005000  9.380000 11.325000  9.700000 ;
      RECT 11.005000 10.010000 11.325000 10.330000 ;
      RECT 11.005000 10.640000 11.325000 10.960000 ;
  END
END sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap
END LIBRARY
