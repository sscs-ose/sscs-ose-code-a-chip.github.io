MACRO PMOS_S_89058261_X6_Y5
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_89058261_X6_Y5 0 0 ;
  SIZE 6880 BY 31080 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 260 3150 24100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3300 4460 3580 28300 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3730 680 4010 30400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 30745 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 30745 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 30745 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 30745 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 30745 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 21505 ;
    LAYER M1 ;
      RECT 5465 21755 5715 22765 ;
    LAYER M1 ;
      RECT 5465 23855 5715 27385 ;
    LAYER M1 ;
      RECT 5465 27635 5715 28645 ;
    LAYER M1 ;
      RECT 5465 29735 5715 30745 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 5895 23855 6145 27385 ;
    LAYER M2 ;
      RECT 1120 280 5760 560 ;
    LAYER M2 ;
      RECT 1120 4480 5760 4760 ;
    LAYER M2 ;
      RECT 690 700 6190 980 ;
    LAYER M2 ;
      RECT 1120 6160 5760 6440 ;
    LAYER M2 ;
      RECT 1120 10360 5760 10640 ;
    LAYER M2 ;
      RECT 690 6580 6190 6860 ;
    LAYER M2 ;
      RECT 1120 12040 5760 12320 ;
    LAYER M2 ;
      RECT 1120 16240 5760 16520 ;
    LAYER M2 ;
      RECT 690 12460 6190 12740 ;
    LAYER M2 ;
      RECT 1120 17920 5760 18200 ;
    LAYER M2 ;
      RECT 1120 22120 5760 22400 ;
    LAYER M2 ;
      RECT 690 18340 6190 18620 ;
    LAYER M2 ;
      RECT 1120 23800 5760 24080 ;
    LAYER M2 ;
      RECT 1120 28000 5760 28280 ;
    LAYER M2 ;
      RECT 1120 30100 5760 30380 ;
    LAYER M2 ;
      RECT 690 24220 6190 24500 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 30155 1375 30325 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 30155 2235 30325 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 30155 3095 30325 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 30155 3955 30325 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 30155 4815 30325 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 17975 5675 18145 ;
    LAYER V1 ;
      RECT 5505 22175 5675 22345 ;
    LAYER V1 ;
      RECT 5505 23855 5675 24025 ;
    LAYER V1 ;
      RECT 5505 28055 5675 28225 ;
    LAYER V1 ;
      RECT 5505 30155 5675 30325 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 5935 18395 6105 18565 ;
    LAYER V1 ;
      RECT 5935 24275 6105 24445 ;
    LAYER V2 ;
      RECT 2935 345 3085 495 ;
    LAYER V2 ;
      RECT 2935 6225 3085 6375 ;
    LAYER V2 ;
      RECT 2935 12105 3085 12255 ;
    LAYER V2 ;
      RECT 2935 17985 3085 18135 ;
    LAYER V2 ;
      RECT 2935 23865 3085 24015 ;
    LAYER V2 ;
      RECT 3365 4545 3515 4695 ;
    LAYER V2 ;
      RECT 3365 10425 3515 10575 ;
    LAYER V2 ;
      RECT 3365 16305 3515 16455 ;
    LAYER V2 ;
      RECT 3365 22185 3515 22335 ;
    LAYER V2 ;
      RECT 3365 28065 3515 28215 ;
    LAYER V2 ;
      RECT 3795 765 3945 915 ;
    LAYER V2 ;
      RECT 3795 6645 3945 6795 ;
    LAYER V2 ;
      RECT 3795 12525 3945 12675 ;
    LAYER V2 ;
      RECT 3795 18405 3945 18555 ;
    LAYER V2 ;
      RECT 3795 24285 3945 24435 ;
    LAYER V2 ;
      RECT 3795 30165 3945 30315 ;
  END
END PMOS_S_89058261_X6_Y5
