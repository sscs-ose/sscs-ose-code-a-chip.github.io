* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
*  Typical Parameters
.param
+ dkisnpn1x1=1.0 dkbfnpn1x1=1.0
+ dkisnpn1x2=1.0 dkbfnpn1x2=1.0
+ dkisnpnpolyhv=1.0 dkbfnpnpolyhv=1.0
.include "sky130_fd_pr__npn_05v5_W1p00L1p00.model.spice"
.include "sky130_fd_pr__npn_05v5_W1p00L2p00.model.spice"
.include "../npn_11v0/sky130_fd_pr__npn_11v0_W1p00L1p00.model.spice"
