* SKY130 Spice File.
.param
+ tol_nfom = 0.0483u
+ tol_pfom = 0.042u
+ tol_nw = 0.0483u
+ tol_poly = 0.0287u
+ tol_li = 0.014u
+ tol_m1 = 0.0175u
+ tol_m2 = 0.0175u
+ tol_m3 = 0.0455u
+ tol_m4 = 0.0455u
+ tol_m5 = 0.119u
+ tol_rdl = 0.7u
.param
+ rcn=103.6
+ rcp=411
+ rdn=111.6
+ rdp=175.3
+ rdn_hv=105.6
+ rdp_hv=169.3
+ rp1=44
+ rnw=1378
+ rl1=10.31
+ rm1=0.111
+ rm2=0.111
+ rm3=0.0407
+ rm4=0.0407
+ rm5=0.02339
+ rrdl=0.0043
+ rcp1=61.28
+ rcl1=3.91
+ rcvia=2.75
+ rcvia2=1.373
+ rcvia3=1.373
+ rcvia4=0.1224
+ rcrdlcon=0.00496
+ rspwres=3512
* P+ Poly Preres Parameters
.param
+ crpf_precision=  8.84e-5   $ Units: farad/meter^2
+ crpfsw_precision_1_1 = 4.67e-11 $ Units: farad/meter
+ crpfsw_precision_2_1 = 5.02e-11 $ Units: farad/meter
+ crpfsw_precision_4_1 = 5.45e-11 $ Units: farad/meter
+ crpfsw_precision_8_2 = 5.96e-11 $ Units: farad/meter
+ crpfsw_precision_16_2 = 6.54e-11 $ Units: farad/meter
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/fast_70p.spice"
