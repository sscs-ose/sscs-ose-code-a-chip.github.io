# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15 ;
  ORIGIN  0.000000 -0.020000 ;
  SIZE  4.400000 BY  3.990000 ;
  PIN DRAIN
    ANTENNADIFFAREA  3.732400 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 2.200000 4.400000 3.480000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.806000 ;
    PORT
      LAYER met1 ;
        RECT 0.820000 0.040000 3.450000 0.330000 ;
        RECT 0.820000 3.700000 3.450000 3.990000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  3.551800 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.550000 4.400000 1.830000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.809100 ;
    PORT
      LAYER met1 ;
        RECT 0.130000 0.820000 0.420000 3.210000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.110000 0.215000 0.440000 3.815000 ;
      RECT 0.690000 0.490000 0.915000 3.540000 ;
      RECT 0.840000 0.100000 3.550000 0.270000 ;
      RECT 0.840000 3.760000 3.550000 3.930000 ;
      RECT 1.165000 0.490000 1.695000 3.540000 ;
      RECT 1.935000 0.490000 2.465000 3.540000 ;
      RECT 2.705000 0.490000 3.235000 3.540000 ;
      RECT 3.485000 0.490000 3.710000 3.540000 ;
      RECT 3.960000 0.215000 4.290000 3.815000 ;
    LAYER mcon ;
      RECT 0.190000 0.850000 0.360000 1.020000 ;
      RECT 0.190000 1.210000 0.360000 1.380000 ;
      RECT 0.190000 1.570000 0.360000 1.740000 ;
      RECT 0.190000 1.930000 0.360000 2.100000 ;
      RECT 0.190000 2.290000 0.360000 2.460000 ;
      RECT 0.190000 2.650000 0.360000 2.820000 ;
      RECT 0.190000 3.010000 0.360000 3.180000 ;
      RECT 0.735000 0.695000 0.905000 0.865000 ;
      RECT 0.735000 1.055000 0.905000 1.225000 ;
      RECT 0.735000 1.415000 0.905000 1.585000 ;
      RECT 0.735000 1.775000 0.905000 1.945000 ;
      RECT 0.735000 2.135000 0.905000 2.305000 ;
      RECT 0.735000 2.495000 0.905000 2.665000 ;
      RECT 0.735000 2.855000 0.905000 3.025000 ;
      RECT 0.735000 3.215000 0.905000 3.385000 ;
      RECT 0.850000 0.100000 1.020000 0.270000 ;
      RECT 0.850000 3.760000 1.020000 3.930000 ;
      RECT 1.165000 0.695000 1.695000 3.385000 ;
      RECT 1.330000 0.100000 1.500000 0.270000 ;
      RECT 1.330000 3.760000 1.500000 3.930000 ;
      RECT 1.810000 0.100000 1.980000 0.270000 ;
      RECT 1.810000 3.760000 1.980000 3.930000 ;
      RECT 1.935000 0.645000 2.465000 3.335000 ;
      RECT 2.290000 0.100000 2.460000 0.270000 ;
      RECT 2.290000 3.760000 2.460000 3.930000 ;
      RECT 2.705000 0.695000 3.235000 3.385000 ;
      RECT 2.770000 0.100000 2.940000 0.270000 ;
      RECT 2.770000 3.760000 2.940000 3.930000 ;
      RECT 3.250000 0.100000 3.420000 0.270000 ;
      RECT 3.250000 3.760000 3.420000 3.930000 ;
      RECT 3.495000 0.695000 3.665000 0.865000 ;
      RECT 3.495000 1.055000 3.665000 1.225000 ;
      RECT 3.495000 1.415000 3.665000 1.585000 ;
      RECT 3.495000 1.775000 3.665000 1.945000 ;
      RECT 3.495000 2.135000 3.665000 2.305000 ;
      RECT 3.495000 2.495000 3.665000 2.665000 ;
      RECT 3.495000 2.855000 3.665000 3.025000 ;
      RECT 3.495000 3.215000 3.665000 3.385000 ;
      RECT 4.040000 0.850000 4.210000 1.020000 ;
      RECT 4.040000 1.210000 4.210000 1.380000 ;
      RECT 4.040000 1.570000 4.210000 1.740000 ;
      RECT 4.040000 1.930000 4.210000 2.100000 ;
      RECT 4.040000 2.290000 4.210000 2.460000 ;
      RECT 4.040000 2.650000 4.210000 2.820000 ;
      RECT 4.040000 3.010000 4.210000 3.180000 ;
    LAYER met1 ;
      RECT 0.690000 0.510000 0.970000 3.520000 ;
      RECT 1.115000 0.510000 1.745000 3.520000 ;
      RECT 1.885000 0.510000 2.515000 3.520000 ;
      RECT 2.655000 0.510000 3.285000 3.520000 ;
      RECT 3.430000 0.510000 3.710000 3.520000 ;
      RECT 3.980000 0.820000 4.270000 3.210000 ;
    LAYER via ;
      RECT 0.700000 0.580000 0.960000 0.840000 ;
      RECT 0.700000 0.900000 0.960000 1.160000 ;
      RECT 0.700000 1.220000 0.960000 1.480000 ;
      RECT 0.700000 1.540000 0.960000 1.800000 ;
      RECT 1.140000 2.230000 1.720000 3.450000 ;
      RECT 1.910000 0.580000 2.490000 1.800000 ;
      RECT 2.680000 2.230000 3.260000 3.450000 ;
      RECT 3.440000 0.580000 3.700000 0.840000 ;
      RECT 3.440000 0.900000 3.700000 1.160000 ;
      RECT 3.440000 1.220000 3.700000 1.480000 ;
      RECT 3.440000 1.540000 3.700000 1.800000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15
END LIBRARY
