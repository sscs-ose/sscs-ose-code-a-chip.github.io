# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.620000 BY  4.030000 ;
  PIN BULK
    ANTENNADIFFAREA  1.745800 ;
    PORT
      LAYER li1 ;
        RECT 0.240000 0.660000 0.410000 3.370000 ;
        RECT 2.210000 0.660000 2.380000 3.370000 ;
      LAYER mcon ;
        RECT 0.240000 0.670000 0.410000 0.840000 ;
        RECT 0.240000 1.030000 0.410000 1.200000 ;
        RECT 0.240000 1.390000 0.410000 1.560000 ;
        RECT 0.240000 1.750000 0.410000 1.920000 ;
        RECT 0.240000 2.110000 0.410000 2.280000 ;
        RECT 0.240000 2.470000 0.410000 2.640000 ;
        RECT 0.240000 2.830000 0.410000 3.000000 ;
        RECT 0.240000 3.190000 0.410000 3.360000 ;
        RECT 2.210000 0.670000 2.380000 0.840000 ;
        RECT 2.210000 1.030000 2.380000 1.200000 ;
        RECT 2.210000 1.390000 2.380000 1.560000 ;
        RECT 2.210000 1.750000 2.380000 1.920000 ;
        RECT 2.210000 2.110000 2.380000 2.280000 ;
        RECT 2.210000 2.470000 2.380000 2.640000 ;
        RECT 2.210000 2.830000 2.380000 3.000000 ;
        RECT 2.210000 3.190000 2.380000 3.360000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.180000 0.610000 0.470000 3.420000 ;
        RECT 2.150000 0.610000 2.440000 3.420000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  0.842800 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 2.140000 2.570000 3.420000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.903000 ;
    PORT
      LAYER li1 ;
        RECT 0.805000 0.100000 1.815000 0.270000 ;
        RECT 0.805000 3.760000 1.815000 3.930000 ;
      LAYER mcon ;
        RECT 0.865000 0.100000 1.035000 0.270000 ;
        RECT 0.865000 3.760000 1.035000 3.930000 ;
        RECT 1.225000 0.100000 1.395000 0.270000 ;
        RECT 1.225000 3.760000 1.395000 3.930000 ;
        RECT 1.585000 0.100000 1.755000 0.270000 ;
        RECT 1.585000 3.760000 1.755000 3.930000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.805000 0.000000 1.815000 0.330000 ;
        RECT 0.805000 3.700000 1.815000 4.030000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.610000 2.570000 1.890000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.795000 0.490000 0.965000 3.540000 ;
      RECT 1.225000 0.490000 1.395000 3.540000 ;
      RECT 1.655000 0.490000 1.825000 3.540000 ;
    LAYER mcon ;
      RECT 0.795000 0.670000 0.965000 0.840000 ;
      RECT 0.795000 1.030000 0.965000 1.200000 ;
      RECT 0.795000 1.390000 0.965000 1.560000 ;
      RECT 0.795000 1.750000 0.965000 1.920000 ;
      RECT 0.795000 2.110000 0.965000 2.280000 ;
      RECT 0.795000 2.470000 0.965000 2.640000 ;
      RECT 0.795000 2.830000 0.965000 3.000000 ;
      RECT 0.795000 3.190000 0.965000 3.360000 ;
      RECT 1.225000 0.670000 1.395000 0.840000 ;
      RECT 1.225000 1.030000 1.395000 1.200000 ;
      RECT 1.225000 1.390000 1.395000 1.560000 ;
      RECT 1.225000 1.750000 1.395000 1.920000 ;
      RECT 1.225000 2.110000 1.395000 2.280000 ;
      RECT 1.225000 2.470000 1.395000 2.640000 ;
      RECT 1.225000 2.830000 1.395000 3.000000 ;
      RECT 1.225000 3.190000 1.395000 3.360000 ;
      RECT 1.655000 0.670000 1.825000 0.840000 ;
      RECT 1.655000 1.030000 1.825000 1.200000 ;
      RECT 1.655000 1.390000 1.825000 1.560000 ;
      RECT 1.655000 1.750000 1.825000 1.920000 ;
      RECT 1.655000 2.110000 1.825000 2.280000 ;
      RECT 1.655000 2.470000 1.825000 2.640000 ;
      RECT 1.655000 2.830000 1.825000 3.000000 ;
      RECT 1.655000 3.190000 1.825000 3.360000 ;
    LAYER met1 ;
      RECT 0.750000 0.610000 1.010000 3.420000 ;
      RECT 1.180000 0.610000 1.440000 3.420000 ;
      RECT 1.610000 0.610000 1.870000 3.420000 ;
    LAYER via ;
      RECT 0.750000 0.640000 1.010000 0.900000 ;
      RECT 0.750000 0.960000 1.010000 1.220000 ;
      RECT 0.750000 1.280000 1.010000 1.540000 ;
      RECT 0.750000 1.600000 1.010000 1.860000 ;
      RECT 1.180000 2.170000 1.440000 2.430000 ;
      RECT 1.180000 2.490000 1.440000 2.750000 ;
      RECT 1.180000 2.810000 1.440000 3.070000 ;
      RECT 1.180000 3.130000 1.440000 3.390000 ;
      RECT 1.610000 0.640000 1.870000 0.900000 ;
      RECT 1.610000 0.960000 1.870000 1.220000 ;
      RECT 1.610000 1.280000 1.870000 1.540000 ;
      RECT 1.610000 1.600000 1.870000 1.860000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15
END LIBRARY
