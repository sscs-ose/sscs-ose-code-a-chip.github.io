# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__esd_rf_nfet_20v0_iec_21vW60p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__esd_rf_nfet_20v0_iec_21vW60p00 ;
  ORIGIN  6.040000  5.910000 ;
  SIZE  13.58000 BY  41.82000 ;
  OBS
    LAYER li1 ;
      RECT -6.040000 -5.910000  7.540000 -4.470000 ;
      RECT -6.040000 -4.470000 -4.480000 34.350000 ;
      RECT -6.040000 34.350000  7.540000 35.910000 ;
      RECT -0.950000 -4.470000  2.445000 -3.255000 ;
      RECT -0.945000 -3.255000  2.445000 -3.245000 ;
      RECT  0.000000  0.000000  1.500000 30.000000 ;
      RECT  5.980000 -4.470000  7.540000 34.350000 ;
    LAYER mcon ;
      RECT -5.810000 -5.785000 -4.560000 35.785000 ;
      RECT -4.195000 -5.785000  5.695000 -4.535000 ;
      RECT -4.195000 34.535000  5.695000 35.785000 ;
      RECT  0.125000  0.155000  1.375000 29.845000 ;
      RECT  6.060000 -5.785000  7.310000 35.785000 ;
    LAYER met1 ;
      POLYGON -3.550000 -1.815000 -3.115000 -2.250000 -3.550000 -2.250000 ;
      POLYGON -3.550000 32.250000 -3.115000 32.250000 -3.550000 31.815000 ;
      POLYGON -3.115000 -2.250000 -1.945000 -3.420000 -3.115000 -3.420000 ;
      POLYGON -3.115000 33.415000 -1.950000 33.415000 -3.115000 32.250000 ;
      POLYGON -2.245000 -1.870000 -2.155000 -1.870000 -2.155000 -1.960000 ;
      POLYGON -2.155000 -1.960000 -1.865000 -1.960000 -1.865000 -2.250000 ;
      POLYGON -2.155000 31.960000 -2.155000 31.870000 -2.245000 31.870000 ;
      POLYGON -1.865000 32.250000 -1.865000 31.960000 -2.155000 31.960000 ;
      POLYGON  3.370000 -1.960000  3.660000 -1.960000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.660000 31.960000  3.370000 31.960000 ;
      POLYGON  3.445000 33.415000  4.610000 33.415000  4.610000 32.250000 ;
      POLYGON  3.660000 -1.870000  3.750000 -1.870000  3.660000 -1.960000 ;
      POLYGON  3.660000 31.960000  3.750000 31.870000  3.660000 31.870000 ;
      POLYGON  4.610000 32.250000  4.900000 32.250000  4.900000 31.960000 ;
      POLYGON  4.620000 -2.250000  4.620000 -3.420000  3.450000 -3.420000 ;
      POLYGON  4.900000 31.960000  5.050000 31.960000  5.050000 31.810000 ;
      POLYGON  4.910000 -1.960000  4.910000 -2.250000  4.620000 -2.250000 ;
      POLYGON  5.050000 -1.820000  5.050000 -1.960000  4.910000 -1.960000 ;
      RECT -6.040000 -5.910000  7.540000 -3.420000 ;
      RECT -6.040000 -3.420000 -3.115000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.550000 32.250000 ;
      RECT -6.040000 32.250000 -3.115000 33.415000 ;
      RECT -6.040000 33.415000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.155000 -1.960000  3.660000 -1.870000 ;
      RECT -2.155000 31.870000  3.660000 31.960000 ;
      RECT -1.865000 -2.250000  3.370000 -1.960000 ;
      RECT -1.865000 31.960000  3.370000 32.250000 ;
      RECT  4.610000 32.250000  7.540000 33.415000 ;
      RECT  4.620000 -3.420000  7.540000 -2.250000 ;
      RECT  4.900000 31.960000  7.540000 32.250000 ;
      RECT  4.910000 -2.250000  7.540000 -1.960000 ;
      RECT  5.050000 -1.960000  7.540000 31.960000 ;
    LAYER met2 ;
      POLYGON -3.550000 -1.815000 -3.115000 -2.250000 -3.550000 -2.250000 ;
      POLYGON -3.550000 32.165000 -3.200000 32.165000 -3.550000 31.815000 ;
      POLYGON -3.200000 33.415000 -1.950000 33.415000 -3.200000 32.165000 ;
      POLYGON -3.115000 -2.250000 -1.945000 -3.420000 -3.115000 -3.420000 ;
      POLYGON -2.245000 -1.870000 -2.130000 -1.870000 -2.130000 -1.985000 ;
      POLYGON -2.130000 -1.985000 -1.865000 -1.985000 -1.865000 -2.250000 ;
      POLYGON -2.130000 31.985000 -2.130000 31.870000 -2.245000 31.870000 ;
      POLYGON -1.950000 32.165000 -1.950000 31.985000 -2.130000 31.985000 ;
      POLYGON -1.865000 32.250000 -1.865000 32.165000 -1.950000 32.165000 ;
      POLYGON  3.370000 -1.985000  3.635000 -1.985000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.445000 32.175000  3.370000 32.175000 ;
      POLYGON  3.445000 32.175000  3.635000 31.985000  3.445000 31.985000 ;
      POLYGON  3.445000 33.415000  4.610000 33.415000  4.610000 32.250000 ;
      POLYGON  3.635000 -1.870000  3.750000 -1.870000  3.635000 -1.985000 ;
      POLYGON  3.635000 31.985000  3.750000 31.870000  3.635000 31.870000 ;
      POLYGON  4.610000 32.250000  4.685000 32.250000  4.685000 32.175000 ;
      POLYGON  4.620000 -2.250000  4.620000 -3.420000  3.450000 -3.420000 ;
      POLYGON  4.685000 32.175000  4.875000 32.175000  4.875000 31.985000 ;
      POLYGON  4.875000 31.985000  5.050000 31.985000  5.050000 31.810000 ;
      POLYGON  4.885000 -1.985000  4.885000 -2.250000  4.620000 -2.250000 ;
      POLYGON  5.050000 -1.820000  5.050000 -1.985000  4.885000 -1.985000 ;
      RECT -6.040000 -5.910000  7.540000 -3.420000 ;
      RECT -6.040000 -3.420000 -3.115000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.550000 32.165000 ;
      RECT -6.040000 32.165000 -3.200000 33.415000 ;
      RECT -6.040000 33.415000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.130000 -1.985000  3.635000 -1.870000 ;
      RECT -2.130000 31.870000  3.635000 31.985000 ;
      RECT -1.950000 31.985000  3.445000 32.165000 ;
      RECT -1.865000 -2.250000  3.370000 -1.985000 ;
      RECT -1.865000 32.165000  3.445000 32.175000 ;
      RECT -1.865000 32.175000  3.370000 32.250000 ;
      RECT  4.610000 32.250000  7.540000 33.415000 ;
      RECT  4.620000 -3.420000  7.540000 -2.250000 ;
      RECT  4.685000 32.175000  7.540000 32.250000 ;
      RECT  4.875000 31.985000  7.540000 32.175000 ;
      RECT  4.885000 -2.250000  7.540000 -1.985000 ;
      RECT  5.050000 -1.985000  7.540000 31.985000 ;
    LAYER met3 ;
      POLYGON -3.550000 -1.815000 -3.115000 -2.250000 -3.550000 -2.250000 ;
      POLYGON -3.550000 32.165000 -3.200000 32.165000 -3.550000 31.815000 ;
      POLYGON -3.200000 33.415000 -1.950000 33.415000 -3.200000 32.165000 ;
      POLYGON -3.115000 -2.250000 -1.945000 -3.420000 -3.115000 -3.420000 ;
      POLYGON -2.245000 -1.870000 -2.125000 -1.870000 -2.125000 -1.990000 ;
      POLYGON -2.125000 -1.990000 -1.865000 -1.990000 -1.865000 -2.250000 ;
      POLYGON -2.125000 31.990000 -2.125000 31.870000 -2.245000 31.870000 ;
      POLYGON -1.950000 32.165000 -1.950000 31.990000 -2.125000 31.990000 ;
      POLYGON -1.865000 32.250000 -1.865000 32.165000 -1.950000 32.165000 ;
      POLYGON  3.370000 -1.990000  3.630000 -1.990000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.445000 32.175000  3.370000 32.175000 ;
      POLYGON  3.445000 32.175000  3.630000 31.990000  3.445000 31.990000 ;
      POLYGON  3.445000 33.415000  4.610000 33.415000  4.610000 32.250000 ;
      POLYGON  3.630000 -1.870000  3.750000 -1.870000  3.630000 -1.990000 ;
      POLYGON  3.630000 31.990000  3.750000 31.870000  3.630000 31.870000 ;
      POLYGON  4.610000 32.250000  4.685000 32.250000  4.685000 32.175000 ;
      POLYGON  4.620000 -2.250000  4.620000 -3.420000  3.450000 -3.420000 ;
      POLYGON  4.685000 32.175000  4.870000 32.175000  4.870000 31.990000 ;
      POLYGON  4.870000 31.990000  5.050000 31.990000  5.050000 31.810000 ;
      POLYGON  4.880000 -1.990000  4.880000 -2.250000  4.620000 -2.250000 ;
      POLYGON  5.050000 -1.820000  5.050000 -1.990000  4.880000 -1.990000 ;
      RECT -6.040000 -5.910000  7.540000 -3.420000 ;
      RECT -6.040000 -3.420000 -3.115000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.550000 32.165000 ;
      RECT -6.040000 32.165000 -3.200000 33.415000 ;
      RECT -6.040000 33.415000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.125000 -1.990000  3.630000 -1.870000 ;
      RECT -2.125000 31.870000  3.630000 31.990000 ;
      RECT -1.950000 31.990000  3.445000 32.165000 ;
      RECT -1.865000 -2.250000  3.370000 -1.990000 ;
      RECT -1.865000 32.165000  3.445000 32.175000 ;
      RECT -1.865000 32.175000  3.370000 32.250000 ;
      RECT  4.610000 32.250000  7.540000 33.415000 ;
      RECT  4.620000 -3.420000  7.540000 -2.250000 ;
      RECT  4.685000 32.175000  7.540000 32.250000 ;
      RECT  4.870000 31.990000  7.540000 32.175000 ;
      RECT  4.880000 -2.250000  7.540000 -1.990000 ;
      RECT  5.050000 -1.990000  7.540000 31.990000 ;
    LAYER met4 ;
      POLYGON -3.550000 -1.815000 -3.115000 -2.250000 -3.550000 -2.250000 ;
      POLYGON -3.550000 32.165000 -3.200000 32.165000 -3.550000 31.815000 ;
      POLYGON -3.200000 33.415000 -1.950000 33.415000 -3.200000 32.165000 ;
      POLYGON -3.115000 -2.250000 -1.945000 -3.420000 -3.115000 -3.420000 ;
      POLYGON -2.245000 -1.870000 -2.150000 -1.870000 -2.150000 -1.965000 ;
      POLYGON -2.155000 31.960000 -2.155000 31.870000 -2.245000 31.870000 ;
      POLYGON -2.150000 -1.965000 -1.865000 -1.965000 -1.865000 -2.250000 ;
      POLYGON -1.950000 32.165000 -1.950000 31.960000 -2.155000 31.960000 ;
      POLYGON -1.865000 32.250000 -1.865000 32.165000 -1.950000 32.165000 ;
      POLYGON  3.370000 -1.965000  3.655000 -1.965000  3.370000 -2.250000 ;
      POLYGON  3.370000 32.250000  3.445000 32.175000  3.370000 32.175000 ;
      POLYGON  3.445000 32.175000  3.655000 31.965000  3.445000 31.965000 ;
      POLYGON  3.445000 33.415000  4.610000 33.415000  4.610000 32.250000 ;
      POLYGON  3.655000 -1.870000  3.750000 -1.870000  3.655000 -1.965000 ;
      POLYGON  3.655000 31.965000  3.750000 31.870000  3.655000 31.870000 ;
      POLYGON  4.610000 32.250000  4.685000 32.250000  4.685000 32.175000 ;
      POLYGON  4.620000 -2.250000  4.620000 -3.420000  3.450000 -3.420000 ;
      POLYGON  4.685000 32.175000  4.895000 32.175000  4.895000 31.965000 ;
      POLYGON  4.895000 31.965000  5.050000 31.965000  5.050000 31.810000 ;
      POLYGON  4.905000 -1.965000  4.905000 -2.250000  4.620000 -2.250000 ;
      POLYGON  5.050000 -1.820000  5.050000 -1.965000  4.905000 -1.965000 ;
      RECT -6.040000 -5.910000  7.540000 -3.420000 ;
      RECT -6.040000 -3.420000 -3.115000 -2.250000 ;
      RECT -6.040000 -2.250000 -3.550000 32.165000 ;
      RECT -6.040000 32.165000 -3.200000 33.415000 ;
      RECT -6.040000 33.415000  7.540000 35.910000 ;
      RECT -2.245000 -1.870000  3.750000 31.870000 ;
      RECT -2.155000 31.870000  3.655000 31.960000 ;
      RECT -2.150000 -1.965000  3.655000 -1.870000 ;
      RECT -1.950000 31.960000  3.655000 31.965000 ;
      RECT -1.950000 31.965000  3.445000 32.165000 ;
      RECT -1.865000 -2.250000  3.370000 -1.965000 ;
      RECT -1.865000 32.165000  3.445000 32.175000 ;
      RECT -1.865000 32.175000  3.370000 32.250000 ;
      RECT  4.610000 32.250000  7.540000 33.415000 ;
      RECT  4.620000 -3.420000  7.540000 -2.250000 ;
      RECT  4.685000 32.175000  7.540000 32.250000 ;
      RECT  4.895000 31.965000  7.540000 32.175000 ;
      RECT  4.905000 -2.250000  7.540000 -1.965000 ;
      RECT  5.050000 -1.965000  7.540000 31.965000 ;
    LAYER met5 ;
      RECT -6.040000 -5.910000 7.540000  4.090000 ;
      RECT -6.040000 25.910000 7.540000 35.910000 ;
      RECT -4.790000  4.090000 6.290000 25.910000 ;
    LAYER via ;
      RECT -5.930000 -5.760000 -3.750000 35.780000 ;
      RECT -3.380000 -5.760000  4.880000 -3.580000 ;
      RECT -3.380000 33.600000  4.880000 35.780000 ;
      RECT -1.940000 -1.930000  3.440000 31.930000 ;
      RECT  5.250000 -5.760000  7.430000 35.780000 ;
    LAYER via2 ;
      RECT -5.875000 -5.740000 -3.595000 35.740000 ;
      RECT -3.190000 -5.745000  4.690000 -3.465000 ;
      RECT -3.190000 33.460000  4.690000 35.740000 ;
      RECT -1.985000 -1.940000  3.495000 31.940000 ;
      RECT  5.095000 -5.740000  7.375000 35.740000 ;
    LAYER via3 ;
      RECT -5.900000 -5.760000 -3.580000 35.760000 ;
      RECT -3.210000 -5.770000  4.710000 -3.450000 ;
      RECT -3.210000 33.445000  4.710000 35.765000 ;
      RECT -2.005000 -1.960000  3.515000 31.960000 ;
      RECT  5.080000 -5.760000  7.400000 35.760000 ;
    LAYER via4 ;
      RECT -2.240000 -1.590000 3.740000 31.590000 ;
  END
END sky130_fd_pr__esd_rf_nfet_20v0_iec_21vW60p00
END LIBRARY
