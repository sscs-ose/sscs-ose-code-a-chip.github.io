* NGSPICE file created from Unnamed_e9e9e382.ext - technology: sky130A

.subckt ota AVSS AVDD INM INP VOUT NBC_10U NB_10U
X0 AVDD a_n14196_2392# a_n14196_2392# AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=49.1712 ps=283.36 w=1.88 l=3 M=4
X2 a_7567_n7591# a_7567_n7591# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X3 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=102.063 ps=586.58 w=4 l=2 M=23.235
X4 VOUT a_n793_n4248# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1 M=2
X5 a_7567_n7591# NB_10U a_4567_n7591# AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X6 a_n793_n4248# a_n3478_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X7 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=0 ps=0 w=3 l=4 M=4
X8 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0 ps=0 w=0.5 l=4 M=4
X9 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=0 ps=0 w=2.75 l=1 M=5.63636
X10 a_4567_n7591# NBC_10U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X11 a_n8111_n7591# NB_10U a_n14196_2392# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X12 NBC_10U NB_10U a_n2123_n7595# AVSS sky130_fd_pr__nfet_01v8 ad=0.68475 pd=4.48 as=1.6185 ps=9.08 w=4.15 l=2 M=2
X13 a_n7071_n377# INM a_n14274_2810# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X14 AVSS NBC_10U a_n2123_n7595# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X15 AVSS NBC_10U a_n8111_n7591# AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X16 a_n3478_1981# a_n2600_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X17 a_n2600_1981# AVSS a_n3478_1981# AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=4
X18 a_n511_n10433# NB_10U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=2
X19 a_n2600_1981# AVDD a_n3478_1981# AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0.195 ps=1.78 w=0.5 l=4
X20 a_4636_n502# a_7567_n7591# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X21 VOUT a_n331_9295# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X22 a_n511_n10433# NB_10U NB_10U AVSS sky130_fd_pr__nfet_01v8 ad=1.6185 pd=9.08 as=0.68475 ps=4.48 w=4.15 l=2 M=2
X23 AVSS a_n14274_2810# a_n7071_n377# AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=1.0725 ps=6.28 w=2.75 l=1
X24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1 M=4
X25 a_n331_9295# a_n2600_1981# AVDD AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.755 pd=9.78 as=1.755 ps=9.78 w=4.5 l=1 M=2
X26 AVDD a_n14196_2392# a_n14274_2810# AVDD sky130_fd_pr__pfet_01v8_lvt ad=0.7332 pd=4.54 as=0.7332 ps=4.54 w=1.88 l=3 M=2
X27 a_n331_9295# AVSS a_n2600_1981# AVDD sky130_fd_pr__pfet_01v8_lvt ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=4
X28 a_n331_9295# INP a_n7071_n377# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X29 a_n331_9295# AVDD a_n2600_1981# AVSS sky130_fd_pr__nfet_01v8_lvt ad=0.195 pd=1.78 as=0.195 ps=1.78 w=0.5 l=4
X30 a_n1678_n502# a_4636_n502# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=1.0725 pd=6.28 as=1.0725 ps=6.28 w=2.75 l=1
X31 a_n793_n4248# a_n793_n4248# AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1 M=2
X32 a_n3478_1981# INM a_n1678_n502# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
X33 a_4636_n502# INP a_n1678_n502# AVSS sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=1.56 ps=8.78 w=4 l=2
.ends

