* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 2
.param
+ sky130_fd_pr__pfet_01v8_mvt__toxe_mult = 0.948
+ sky130_fd_pr__pfet_01v8_mvt__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8_mvt__overlap_mult = 0.95436
+ sky130_fd_pr__pfet_01v8_mvt__ajunction_mult = 0.90161
+ sky130_fd_pr__pfet_01v8_mvt__pjunction_mult = 0.90587
+ sky130_fd_pr__pfet_01v8_mvt__wint_diff = -3.2175e-8
+ sky130_fd_pr__pfet_01v8_mvt__lint_diff = 1.7325e-8
+ sky130_fd_pr__pfet_01v8_mvt__dlc_diff = 1.7325e-8
+ sky130_fd_pr__pfet_01v8_mvt__dwc_diff = -3.2175e-8
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult = 0.85
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult = 0.75
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult = 0.75
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult_2 = 0.65
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult_2 = 0.65
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rs_mult = 1.0
*
* sky130_fd_pr__pfet_01v8_mvt, Bin 000, W = 1.68, L = 0.15
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_mvt__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__voff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__vsat_diff_0 = -14993.0
+ sky130_fd_pr__pfet_01v8_mvt__ua_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__u0_diff_0 = -0.00014433
+ sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__ub_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__k2_diff_0 = -0.32
+ sky130_fd_pr__pfet_01v8_mvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__vth0_diff_0 = 0.11281
+ sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__a0_diff_0 = 0.0
*
* sky130_fd_pr__pfet_01v8_mvt, Bin 001, W = 0.84, L = 0.15
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_mvt__a0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__voff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__vsat_diff_1 = -13854.0
+ sky130_fd_pr__pfet_01v8_mvt__ua_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__u0_diff_1 = -0.00018259
+ sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__ub_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__ags_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__k2_diff_1 = -0.26031
+ sky130_fd_pr__pfet_01v8_mvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_mvt__vth0_diff_1 = 0.23239
+ sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_1 = 0.0
.include "../pfet_01v8_mvt/sky130_fd_pr__pfet_01v8_mvt.pm3.spice"
