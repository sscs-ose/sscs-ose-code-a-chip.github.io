# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  6.670000 BY  6.940000 ;
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 3.595000 6.740000 5.955000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  10.099999 ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.000000 4.810000 0.685000 ;
        RECT 2.000000 6.255000 4.810000 6.940000 ;
      LAYER mcon ;
        RECT 2.060000 0.095000 4.750000 0.625000 ;
        RECT 2.060000 6.315000 4.750000 6.845000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.000000 0.000000 4.810000 0.685000 ;
        RECT 2.000000 6.255000 4.810000 6.940000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 0.985000 6.740000 3.345000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  5.050000 ;
    ANTENNAGATEAREA  2.525000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 0.985000 0.500000 5.955000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.310000 0.985000 6.605000 5.955000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 1.150000 6.015000 ;
      RECT 0.950000 0.485000 1.280000 0.815000 ;
      RECT 0.950000 0.815000 1.150000 0.925000 ;
      RECT 0.950000 6.015000 1.150000 6.125000 ;
      RECT 0.950000 6.125000 1.280000 6.455000 ;
      RECT 1.760000 0.925000 1.930000 6.015000 ;
      RECT 2.540000 0.925000 2.710000 6.015000 ;
      RECT 3.320000 0.925000 3.490000 6.015000 ;
      RECT 4.100000 0.925000 4.270000 6.015000 ;
      RECT 4.880000 0.925000 5.050000 6.015000 ;
      RECT 5.530000 0.485000 5.860000 0.815000 ;
      RECT 5.530000 6.125000 5.860000 6.455000 ;
      RECT 5.660000 0.815000 5.860000 0.925000 ;
      RECT 5.660000 0.925000 6.605000 6.015000 ;
      RECT 5.660000 6.015000 5.860000 6.125000 ;
    LAYER mcon ;
      RECT 0.300000 1.045000 0.470000 1.215000 ;
      RECT 0.300000 1.405000 0.470000 1.575000 ;
      RECT 0.300000 1.765000 0.470000 1.935000 ;
      RECT 0.300000 2.125000 0.470000 2.295000 ;
      RECT 0.300000 2.485000 0.470000 2.655000 ;
      RECT 0.300000 2.845000 0.470000 3.015000 ;
      RECT 0.300000 3.205000 0.470000 3.375000 ;
      RECT 0.300000 3.565000 0.470000 3.735000 ;
      RECT 0.300000 3.925000 0.470000 4.095000 ;
      RECT 0.300000 4.285000 0.470000 4.455000 ;
      RECT 0.300000 4.645000 0.470000 4.815000 ;
      RECT 0.300000 5.005000 0.470000 5.175000 ;
      RECT 0.300000 5.365000 0.470000 5.535000 ;
      RECT 0.300000 5.725000 0.470000 5.895000 ;
      RECT 1.760000 1.045000 1.930000 1.215000 ;
      RECT 1.760000 1.405000 1.930000 1.575000 ;
      RECT 1.760000 1.765000 1.930000 1.935000 ;
      RECT 1.760000 2.125000 1.930000 2.295000 ;
      RECT 1.760000 2.485000 1.930000 2.655000 ;
      RECT 1.760000 2.845000 1.930000 3.015000 ;
      RECT 1.760000 3.205000 1.930000 3.375000 ;
      RECT 1.760000 3.565000 1.930000 3.735000 ;
      RECT 1.760000 3.925000 1.930000 4.095000 ;
      RECT 1.760000 4.285000 1.930000 4.455000 ;
      RECT 1.760000 4.645000 1.930000 4.815000 ;
      RECT 1.760000 5.005000 1.930000 5.175000 ;
      RECT 1.760000 5.365000 1.930000 5.535000 ;
      RECT 1.760000 5.725000 1.930000 5.895000 ;
      RECT 2.540000 1.045000 2.710000 1.215000 ;
      RECT 2.540000 1.405000 2.710000 1.575000 ;
      RECT 2.540000 1.765000 2.710000 1.935000 ;
      RECT 2.540000 2.125000 2.710000 2.295000 ;
      RECT 2.540000 2.485000 2.710000 2.655000 ;
      RECT 2.540000 2.845000 2.710000 3.015000 ;
      RECT 2.540000 3.205000 2.710000 3.375000 ;
      RECT 2.540000 3.565000 2.710000 3.735000 ;
      RECT 2.540000 3.925000 2.710000 4.095000 ;
      RECT 2.540000 4.285000 2.710000 4.455000 ;
      RECT 2.540000 4.645000 2.710000 4.815000 ;
      RECT 2.540000 5.005000 2.710000 5.175000 ;
      RECT 2.540000 5.365000 2.710000 5.535000 ;
      RECT 2.540000 5.725000 2.710000 5.895000 ;
      RECT 3.320000 1.045000 3.490000 1.215000 ;
      RECT 3.320000 1.405000 3.490000 1.575000 ;
      RECT 3.320000 1.765000 3.490000 1.935000 ;
      RECT 3.320000 2.125000 3.490000 2.295000 ;
      RECT 3.320000 2.485000 3.490000 2.655000 ;
      RECT 3.320000 2.845000 3.490000 3.015000 ;
      RECT 3.320000 3.205000 3.490000 3.375000 ;
      RECT 3.320000 3.565000 3.490000 3.735000 ;
      RECT 3.320000 3.925000 3.490000 4.095000 ;
      RECT 3.320000 4.285000 3.490000 4.455000 ;
      RECT 3.320000 4.645000 3.490000 4.815000 ;
      RECT 3.320000 5.005000 3.490000 5.175000 ;
      RECT 3.320000 5.365000 3.490000 5.535000 ;
      RECT 3.320000 5.725000 3.490000 5.895000 ;
      RECT 4.100000 1.045000 4.270000 1.215000 ;
      RECT 4.100000 1.405000 4.270000 1.575000 ;
      RECT 4.100000 1.765000 4.270000 1.935000 ;
      RECT 4.100000 2.125000 4.270000 2.295000 ;
      RECT 4.100000 2.485000 4.270000 2.655000 ;
      RECT 4.100000 2.845000 4.270000 3.015000 ;
      RECT 4.100000 3.205000 4.270000 3.375000 ;
      RECT 4.100000 3.565000 4.270000 3.735000 ;
      RECT 4.100000 3.925000 4.270000 4.095000 ;
      RECT 4.100000 4.285000 4.270000 4.455000 ;
      RECT 4.100000 4.645000 4.270000 4.815000 ;
      RECT 4.100000 5.005000 4.270000 5.175000 ;
      RECT 4.100000 5.365000 4.270000 5.535000 ;
      RECT 4.100000 5.725000 4.270000 5.895000 ;
      RECT 4.880000 1.045000 5.050000 1.215000 ;
      RECT 4.880000 1.405000 5.050000 1.575000 ;
      RECT 4.880000 1.765000 5.050000 1.935000 ;
      RECT 4.880000 2.125000 5.050000 2.295000 ;
      RECT 4.880000 2.485000 5.050000 2.655000 ;
      RECT 4.880000 2.845000 5.050000 3.015000 ;
      RECT 4.880000 3.205000 5.050000 3.375000 ;
      RECT 4.880000 3.565000 5.050000 3.735000 ;
      RECT 4.880000 3.925000 5.050000 4.095000 ;
      RECT 4.880000 4.285000 5.050000 4.455000 ;
      RECT 4.880000 4.645000 5.050000 4.815000 ;
      RECT 4.880000 5.005000 5.050000 5.175000 ;
      RECT 4.880000 5.365000 5.050000 5.535000 ;
      RECT 4.880000 5.725000 5.050000 5.895000 ;
      RECT 6.340000 1.045000 6.510000 1.215000 ;
      RECT 6.340000 1.405000 6.510000 1.575000 ;
      RECT 6.340000 1.765000 6.510000 1.935000 ;
      RECT 6.340000 2.125000 6.510000 2.295000 ;
      RECT 6.340000 2.485000 6.510000 2.655000 ;
      RECT 6.340000 2.845000 6.510000 3.015000 ;
      RECT 6.340000 3.205000 6.510000 3.375000 ;
      RECT 6.340000 3.565000 6.510000 3.735000 ;
      RECT 6.340000 3.925000 6.510000 4.095000 ;
      RECT 6.340000 4.285000 6.510000 4.455000 ;
      RECT 6.340000 4.645000 6.510000 4.815000 ;
      RECT 6.340000 5.005000 6.510000 5.175000 ;
      RECT 6.340000 5.365000 6.510000 5.535000 ;
      RECT 6.340000 5.725000 6.510000 5.895000 ;
    LAYER met1 ;
      RECT 1.715000 0.985000 1.975000 5.955000 ;
      RECT 2.495000 0.985000 2.755000 5.955000 ;
      RECT 3.275000 0.985000 3.535000 5.955000 ;
      RECT 4.055000 0.985000 4.315000 5.955000 ;
      RECT 4.835000 0.985000 5.095000 5.955000 ;
    LAYER via ;
      RECT 1.715000 1.015000 1.975000 1.275000 ;
      RECT 1.715000 1.335000 1.975000 1.595000 ;
      RECT 1.715000 1.655000 1.975000 1.915000 ;
      RECT 1.715000 1.975000 1.975000 2.235000 ;
      RECT 1.715000 2.295000 1.975000 2.555000 ;
      RECT 1.715000 2.615000 1.975000 2.875000 ;
      RECT 1.715000 2.935000 1.975000 3.195000 ;
      RECT 2.495000 3.745000 2.755000 4.005000 ;
      RECT 2.495000 4.065000 2.755000 4.325000 ;
      RECT 2.495000 4.385000 2.755000 4.645000 ;
      RECT 2.495000 4.705000 2.755000 4.965000 ;
      RECT 2.495000 5.025000 2.755000 5.285000 ;
      RECT 2.495000 5.345000 2.755000 5.605000 ;
      RECT 2.495000 5.665000 2.755000 5.925000 ;
      RECT 3.275000 1.015000 3.535000 1.275000 ;
      RECT 3.275000 1.335000 3.535000 1.595000 ;
      RECT 3.275000 1.655000 3.535000 1.915000 ;
      RECT 3.275000 1.975000 3.535000 2.235000 ;
      RECT 3.275000 2.295000 3.535000 2.555000 ;
      RECT 3.275000 2.615000 3.535000 2.875000 ;
      RECT 3.275000 2.935000 3.535000 3.195000 ;
      RECT 4.055000 3.745000 4.315000 4.005000 ;
      RECT 4.055000 4.065000 4.315000 4.325000 ;
      RECT 4.055000 4.385000 4.315000 4.645000 ;
      RECT 4.055000 4.705000 4.315000 4.965000 ;
      RECT 4.055000 5.025000 4.315000 5.285000 ;
      RECT 4.055000 5.345000 4.315000 5.605000 ;
      RECT 4.055000 5.665000 4.315000 5.925000 ;
      RECT 4.835000 1.015000 5.095000 1.275000 ;
      RECT 4.835000 1.335000 5.095000 1.595000 ;
      RECT 4.835000 1.655000 5.095000 1.915000 ;
      RECT 4.835000 1.975000 5.095000 2.235000 ;
      RECT 4.835000 2.295000 5.095000 2.555000 ;
      RECT 4.835000 2.615000 5.095000 2.875000 ;
      RECT 4.835000 2.935000 5.095000 3.195000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50
END LIBRARY
