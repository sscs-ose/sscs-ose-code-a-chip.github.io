* NGSPICE file created from clockdiv.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

.subckt clockdiv VDD VSS clk outclkdiv1 outclkdiv2 outclkdiv4 rst_n
XFILLER_0_9_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I rst_n VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_clk clk clknet_0_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 rst_n net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_0_clk_I clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_8_ clknet_1_0__leaf_clk net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7_ _1_ net1 clknet_1_1__leaf_clk net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6_ _0_ net1 clknet_1_0__leaf_clk net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5_ net3 _0_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4_ _2_ _1_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3_ net4 net3 _2_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput2 net2 outclkdiv1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput3 net3 outclkdiv2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput4 net4 outclkdiv4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

