# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  11.35000 BY  8.980000 ;
  PIN DRAIN
    ANTENNADIFFAREA  9.926000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.890000 11.420000 6.090000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  35.450001 ;
    PORT
      LAYER met1 ;
        RECT 1.905000 0.000000 9.585000 0.685000 ;
        RECT 1.905000 8.295000 9.585000 8.980000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  11.91120 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.010000 11.420000 2.610000 ;
        RECT 0.070000 6.370000 11.420000 7.970000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  7.090000 ;
    ANTENNAGATEAREA  3.545000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.010000 0.500000 7.970000 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.990000 1.010000 11.285000 7.970000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT  0.205000 0.925000  1.150000 8.055000 ;
      RECT  0.950000 0.485000  1.280000 0.815000 ;
      RECT  0.950000 0.815000  1.150000 0.925000 ;
      RECT  0.950000 8.055000  1.150000 8.165000 ;
      RECT  0.950000 8.165000  1.280000 8.495000 ;
      RECT  1.760000 0.925000  1.930000 8.055000 ;
      RECT  1.925000 0.000000  9.565000 0.685000 ;
      RECT  1.925000 8.295000  9.565000 8.980000 ;
      RECT  2.540000 0.925000  2.710000 8.055000 ;
      RECT  3.320000 0.925000  3.490000 8.055000 ;
      RECT  4.100000 0.925000  4.270000 8.055000 ;
      RECT  4.880000 0.925000  5.050000 8.055000 ;
      RECT  5.660000 0.925000  5.830000 8.055000 ;
      RECT  6.440000 0.925000  6.610000 8.055000 ;
      RECT  7.220000 0.925000  7.390000 8.055000 ;
      RECT  8.000000 0.925000  8.170000 8.055000 ;
      RECT  8.780000 0.925000  8.950000 8.055000 ;
      RECT  9.560000 0.925000  9.730000 8.055000 ;
      RECT 10.210000 0.485000 10.540000 0.815000 ;
      RECT 10.210000 8.165000 10.540000 8.495000 ;
      RECT 10.340000 0.815000 10.540000 0.925000 ;
      RECT 10.340000 0.925000 11.285000 8.055000 ;
      RECT 10.340000 8.055000 10.540000 8.165000 ;
    LAYER mcon ;
      RECT  0.300000 1.165000  0.470000 1.335000 ;
      RECT  0.300000 1.525000  0.470000 1.695000 ;
      RECT  0.300000 1.885000  0.470000 2.055000 ;
      RECT  0.300000 2.245000  0.470000 2.415000 ;
      RECT  0.300000 2.605000  0.470000 2.775000 ;
      RECT  0.300000 2.965000  0.470000 3.135000 ;
      RECT  0.300000 3.325000  0.470000 3.495000 ;
      RECT  0.300000 3.685000  0.470000 3.855000 ;
      RECT  0.300000 4.045000  0.470000 4.215000 ;
      RECT  0.300000 4.405000  0.470000 4.575000 ;
      RECT  0.300000 4.765000  0.470000 4.935000 ;
      RECT  0.300000 5.125000  0.470000 5.295000 ;
      RECT  0.300000 5.485000  0.470000 5.655000 ;
      RECT  0.300000 5.845000  0.470000 6.015000 ;
      RECT  0.300000 6.205000  0.470000 6.375000 ;
      RECT  0.300000 6.565000  0.470000 6.735000 ;
      RECT  0.300000 6.925000  0.470000 7.095000 ;
      RECT  0.300000 7.285000  0.470000 7.455000 ;
      RECT  0.300000 7.645000  0.470000 7.815000 ;
      RECT  1.760000 1.165000  1.930000 1.335000 ;
      RECT  1.760000 1.525000  1.930000 1.695000 ;
      RECT  1.760000 1.885000  1.930000 2.055000 ;
      RECT  1.760000 2.245000  1.930000 2.415000 ;
      RECT  1.760000 2.605000  1.930000 2.775000 ;
      RECT  1.760000 2.965000  1.930000 3.135000 ;
      RECT  1.760000 3.325000  1.930000 3.495000 ;
      RECT  1.760000 3.685000  1.930000 3.855000 ;
      RECT  1.760000 4.045000  1.930000 4.215000 ;
      RECT  1.760000 4.405000  1.930000 4.575000 ;
      RECT  1.760000 4.765000  1.930000 4.935000 ;
      RECT  1.760000 5.125000  1.930000 5.295000 ;
      RECT  1.760000 5.485000  1.930000 5.655000 ;
      RECT  1.760000 5.845000  1.930000 6.015000 ;
      RECT  1.760000 6.205000  1.930000 6.375000 ;
      RECT  1.760000 6.565000  1.930000 6.735000 ;
      RECT  1.760000 6.925000  1.930000 7.095000 ;
      RECT  1.760000 7.285000  1.930000 7.455000 ;
      RECT  1.760000 7.645000  1.930000 7.815000 ;
      RECT  2.060000 0.095000  9.430000 0.625000 ;
      RECT  2.060000 8.355000  9.430000 8.885000 ;
      RECT  2.540000 1.165000  2.710000 1.335000 ;
      RECT  2.540000 1.525000  2.710000 1.695000 ;
      RECT  2.540000 1.885000  2.710000 2.055000 ;
      RECT  2.540000 2.245000  2.710000 2.415000 ;
      RECT  2.540000 2.605000  2.710000 2.775000 ;
      RECT  2.540000 2.965000  2.710000 3.135000 ;
      RECT  2.540000 3.325000  2.710000 3.495000 ;
      RECT  2.540000 3.685000  2.710000 3.855000 ;
      RECT  2.540000 4.045000  2.710000 4.215000 ;
      RECT  2.540000 4.405000  2.710000 4.575000 ;
      RECT  2.540000 4.765000  2.710000 4.935000 ;
      RECT  2.540000 5.125000  2.710000 5.295000 ;
      RECT  2.540000 5.485000  2.710000 5.655000 ;
      RECT  2.540000 5.845000  2.710000 6.015000 ;
      RECT  2.540000 6.205000  2.710000 6.375000 ;
      RECT  2.540000 6.565000  2.710000 6.735000 ;
      RECT  2.540000 6.925000  2.710000 7.095000 ;
      RECT  2.540000 7.285000  2.710000 7.455000 ;
      RECT  2.540000 7.645000  2.710000 7.815000 ;
      RECT  3.320000 1.165000  3.490000 1.335000 ;
      RECT  3.320000 1.525000  3.490000 1.695000 ;
      RECT  3.320000 1.885000  3.490000 2.055000 ;
      RECT  3.320000 2.245000  3.490000 2.415000 ;
      RECT  3.320000 2.605000  3.490000 2.775000 ;
      RECT  3.320000 2.965000  3.490000 3.135000 ;
      RECT  3.320000 3.325000  3.490000 3.495000 ;
      RECT  3.320000 3.685000  3.490000 3.855000 ;
      RECT  3.320000 4.045000  3.490000 4.215000 ;
      RECT  3.320000 4.405000  3.490000 4.575000 ;
      RECT  3.320000 4.765000  3.490000 4.935000 ;
      RECT  3.320000 5.125000  3.490000 5.295000 ;
      RECT  3.320000 5.485000  3.490000 5.655000 ;
      RECT  3.320000 5.845000  3.490000 6.015000 ;
      RECT  3.320000 6.205000  3.490000 6.375000 ;
      RECT  3.320000 6.565000  3.490000 6.735000 ;
      RECT  3.320000 6.925000  3.490000 7.095000 ;
      RECT  3.320000 7.285000  3.490000 7.455000 ;
      RECT  3.320000 7.645000  3.490000 7.815000 ;
      RECT  4.100000 1.165000  4.270000 1.335000 ;
      RECT  4.100000 1.525000  4.270000 1.695000 ;
      RECT  4.100000 1.885000  4.270000 2.055000 ;
      RECT  4.100000 2.245000  4.270000 2.415000 ;
      RECT  4.100000 2.605000  4.270000 2.775000 ;
      RECT  4.100000 2.965000  4.270000 3.135000 ;
      RECT  4.100000 3.325000  4.270000 3.495000 ;
      RECT  4.100000 3.685000  4.270000 3.855000 ;
      RECT  4.100000 4.045000  4.270000 4.215000 ;
      RECT  4.100000 4.405000  4.270000 4.575000 ;
      RECT  4.100000 4.765000  4.270000 4.935000 ;
      RECT  4.100000 5.125000  4.270000 5.295000 ;
      RECT  4.100000 5.485000  4.270000 5.655000 ;
      RECT  4.100000 5.845000  4.270000 6.015000 ;
      RECT  4.100000 6.205000  4.270000 6.375000 ;
      RECT  4.100000 6.565000  4.270000 6.735000 ;
      RECT  4.100000 6.925000  4.270000 7.095000 ;
      RECT  4.100000 7.285000  4.270000 7.455000 ;
      RECT  4.100000 7.645000  4.270000 7.815000 ;
      RECT  4.880000 1.165000  5.050000 1.335000 ;
      RECT  4.880000 1.525000  5.050000 1.695000 ;
      RECT  4.880000 1.885000  5.050000 2.055000 ;
      RECT  4.880000 2.245000  5.050000 2.415000 ;
      RECT  4.880000 2.605000  5.050000 2.775000 ;
      RECT  4.880000 2.965000  5.050000 3.135000 ;
      RECT  4.880000 3.325000  5.050000 3.495000 ;
      RECT  4.880000 3.685000  5.050000 3.855000 ;
      RECT  4.880000 4.045000  5.050000 4.215000 ;
      RECT  4.880000 4.405000  5.050000 4.575000 ;
      RECT  4.880000 4.765000  5.050000 4.935000 ;
      RECT  4.880000 5.125000  5.050000 5.295000 ;
      RECT  4.880000 5.485000  5.050000 5.655000 ;
      RECT  4.880000 5.845000  5.050000 6.015000 ;
      RECT  4.880000 6.205000  5.050000 6.375000 ;
      RECT  4.880000 6.565000  5.050000 6.735000 ;
      RECT  4.880000 6.925000  5.050000 7.095000 ;
      RECT  4.880000 7.285000  5.050000 7.455000 ;
      RECT  4.880000 7.645000  5.050000 7.815000 ;
      RECT  5.660000 1.165000  5.830000 1.335000 ;
      RECT  5.660000 1.525000  5.830000 1.695000 ;
      RECT  5.660000 1.885000  5.830000 2.055000 ;
      RECT  5.660000 2.245000  5.830000 2.415000 ;
      RECT  5.660000 2.605000  5.830000 2.775000 ;
      RECT  5.660000 2.965000  5.830000 3.135000 ;
      RECT  5.660000 3.325000  5.830000 3.495000 ;
      RECT  5.660000 3.685000  5.830000 3.855000 ;
      RECT  5.660000 4.045000  5.830000 4.215000 ;
      RECT  5.660000 4.405000  5.830000 4.575000 ;
      RECT  5.660000 4.765000  5.830000 4.935000 ;
      RECT  5.660000 5.125000  5.830000 5.295000 ;
      RECT  5.660000 5.485000  5.830000 5.655000 ;
      RECT  5.660000 5.845000  5.830000 6.015000 ;
      RECT  5.660000 6.205000  5.830000 6.375000 ;
      RECT  5.660000 6.565000  5.830000 6.735000 ;
      RECT  5.660000 6.925000  5.830000 7.095000 ;
      RECT  5.660000 7.285000  5.830000 7.455000 ;
      RECT  5.660000 7.645000  5.830000 7.815000 ;
      RECT  6.440000 1.165000  6.610000 1.335000 ;
      RECT  6.440000 1.525000  6.610000 1.695000 ;
      RECT  6.440000 1.885000  6.610000 2.055000 ;
      RECT  6.440000 2.245000  6.610000 2.415000 ;
      RECT  6.440000 2.605000  6.610000 2.775000 ;
      RECT  6.440000 2.965000  6.610000 3.135000 ;
      RECT  6.440000 3.325000  6.610000 3.495000 ;
      RECT  6.440000 3.685000  6.610000 3.855000 ;
      RECT  6.440000 4.045000  6.610000 4.215000 ;
      RECT  6.440000 4.405000  6.610000 4.575000 ;
      RECT  6.440000 4.765000  6.610000 4.935000 ;
      RECT  6.440000 5.125000  6.610000 5.295000 ;
      RECT  6.440000 5.485000  6.610000 5.655000 ;
      RECT  6.440000 5.845000  6.610000 6.015000 ;
      RECT  6.440000 6.205000  6.610000 6.375000 ;
      RECT  6.440000 6.565000  6.610000 6.735000 ;
      RECT  6.440000 6.925000  6.610000 7.095000 ;
      RECT  6.440000 7.285000  6.610000 7.455000 ;
      RECT  6.440000 7.645000  6.610000 7.815000 ;
      RECT  7.220000 1.165000  7.390000 1.335000 ;
      RECT  7.220000 1.525000  7.390000 1.695000 ;
      RECT  7.220000 1.885000  7.390000 2.055000 ;
      RECT  7.220000 2.245000  7.390000 2.415000 ;
      RECT  7.220000 2.605000  7.390000 2.775000 ;
      RECT  7.220000 2.965000  7.390000 3.135000 ;
      RECT  7.220000 3.325000  7.390000 3.495000 ;
      RECT  7.220000 3.685000  7.390000 3.855000 ;
      RECT  7.220000 4.045000  7.390000 4.215000 ;
      RECT  7.220000 4.405000  7.390000 4.575000 ;
      RECT  7.220000 4.765000  7.390000 4.935000 ;
      RECT  7.220000 5.125000  7.390000 5.295000 ;
      RECT  7.220000 5.485000  7.390000 5.655000 ;
      RECT  7.220000 5.845000  7.390000 6.015000 ;
      RECT  7.220000 6.205000  7.390000 6.375000 ;
      RECT  7.220000 6.565000  7.390000 6.735000 ;
      RECT  7.220000 6.925000  7.390000 7.095000 ;
      RECT  7.220000 7.285000  7.390000 7.455000 ;
      RECT  7.220000 7.645000  7.390000 7.815000 ;
      RECT  8.000000 1.165000  8.170000 1.335000 ;
      RECT  8.000000 1.525000  8.170000 1.695000 ;
      RECT  8.000000 1.885000  8.170000 2.055000 ;
      RECT  8.000000 2.245000  8.170000 2.415000 ;
      RECT  8.000000 2.605000  8.170000 2.775000 ;
      RECT  8.000000 2.965000  8.170000 3.135000 ;
      RECT  8.000000 3.325000  8.170000 3.495000 ;
      RECT  8.000000 3.685000  8.170000 3.855000 ;
      RECT  8.000000 4.045000  8.170000 4.215000 ;
      RECT  8.000000 4.405000  8.170000 4.575000 ;
      RECT  8.000000 4.765000  8.170000 4.935000 ;
      RECT  8.000000 5.125000  8.170000 5.295000 ;
      RECT  8.000000 5.485000  8.170000 5.655000 ;
      RECT  8.000000 5.845000  8.170000 6.015000 ;
      RECT  8.000000 6.205000  8.170000 6.375000 ;
      RECT  8.000000 6.565000  8.170000 6.735000 ;
      RECT  8.000000 6.925000  8.170000 7.095000 ;
      RECT  8.000000 7.285000  8.170000 7.455000 ;
      RECT  8.000000 7.645000  8.170000 7.815000 ;
      RECT  8.780000 1.165000  8.950000 1.335000 ;
      RECT  8.780000 1.525000  8.950000 1.695000 ;
      RECT  8.780000 1.885000  8.950000 2.055000 ;
      RECT  8.780000 2.245000  8.950000 2.415000 ;
      RECT  8.780000 2.605000  8.950000 2.775000 ;
      RECT  8.780000 2.965000  8.950000 3.135000 ;
      RECT  8.780000 3.325000  8.950000 3.495000 ;
      RECT  8.780000 3.685000  8.950000 3.855000 ;
      RECT  8.780000 4.045000  8.950000 4.215000 ;
      RECT  8.780000 4.405000  8.950000 4.575000 ;
      RECT  8.780000 4.765000  8.950000 4.935000 ;
      RECT  8.780000 5.125000  8.950000 5.295000 ;
      RECT  8.780000 5.485000  8.950000 5.655000 ;
      RECT  8.780000 5.845000  8.950000 6.015000 ;
      RECT  8.780000 6.205000  8.950000 6.375000 ;
      RECT  8.780000 6.565000  8.950000 6.735000 ;
      RECT  8.780000 6.925000  8.950000 7.095000 ;
      RECT  8.780000 7.285000  8.950000 7.455000 ;
      RECT  8.780000 7.645000  8.950000 7.815000 ;
      RECT  9.560000 1.165000  9.730000 1.335000 ;
      RECT  9.560000 1.525000  9.730000 1.695000 ;
      RECT  9.560000 1.885000  9.730000 2.055000 ;
      RECT  9.560000 2.245000  9.730000 2.415000 ;
      RECT  9.560000 2.605000  9.730000 2.775000 ;
      RECT  9.560000 2.965000  9.730000 3.135000 ;
      RECT  9.560000 3.325000  9.730000 3.495000 ;
      RECT  9.560000 3.685000  9.730000 3.855000 ;
      RECT  9.560000 4.045000  9.730000 4.215000 ;
      RECT  9.560000 4.405000  9.730000 4.575000 ;
      RECT  9.560000 4.765000  9.730000 4.935000 ;
      RECT  9.560000 5.125000  9.730000 5.295000 ;
      RECT  9.560000 5.485000  9.730000 5.655000 ;
      RECT  9.560000 5.845000  9.730000 6.015000 ;
      RECT  9.560000 6.205000  9.730000 6.375000 ;
      RECT  9.560000 6.565000  9.730000 6.735000 ;
      RECT  9.560000 6.925000  9.730000 7.095000 ;
      RECT  9.560000 7.285000  9.730000 7.455000 ;
      RECT  9.560000 7.645000  9.730000 7.815000 ;
      RECT 11.020000 1.165000 11.190000 1.335000 ;
      RECT 11.020000 1.525000 11.190000 1.695000 ;
      RECT 11.020000 1.885000 11.190000 2.055000 ;
      RECT 11.020000 2.245000 11.190000 2.415000 ;
      RECT 11.020000 2.605000 11.190000 2.775000 ;
      RECT 11.020000 2.965000 11.190000 3.135000 ;
      RECT 11.020000 3.325000 11.190000 3.495000 ;
      RECT 11.020000 3.685000 11.190000 3.855000 ;
      RECT 11.020000 4.045000 11.190000 4.215000 ;
      RECT 11.020000 4.405000 11.190000 4.575000 ;
      RECT 11.020000 4.765000 11.190000 4.935000 ;
      RECT 11.020000 5.125000 11.190000 5.295000 ;
      RECT 11.020000 5.485000 11.190000 5.655000 ;
      RECT 11.020000 5.845000 11.190000 6.015000 ;
      RECT 11.020000 6.205000 11.190000 6.375000 ;
      RECT 11.020000 6.565000 11.190000 6.735000 ;
      RECT 11.020000 6.925000 11.190000 7.095000 ;
      RECT 11.020000 7.285000 11.190000 7.455000 ;
      RECT 11.020000 7.645000 11.190000 7.815000 ;
    LAYER met1 ;
      RECT 1.715000 1.010000 1.975000 7.970000 ;
      RECT 2.495000 1.010000 2.755000 7.970000 ;
      RECT 3.275000 1.010000 3.535000 7.970000 ;
      RECT 4.055000 1.010000 4.315000 7.970000 ;
      RECT 4.835000 1.010000 5.095000 7.970000 ;
      RECT 5.615000 1.010000 5.875000 7.970000 ;
      RECT 6.395000 1.010000 6.655000 7.970000 ;
      RECT 7.175000 1.010000 7.435000 7.970000 ;
      RECT 7.955000 1.010000 8.215000 7.970000 ;
      RECT 8.735000 1.010000 8.995000 7.970000 ;
      RECT 9.515000 1.010000 9.775000 7.970000 ;
    LAYER via ;
      RECT 1.715000 1.040000 1.975000 1.300000 ;
      RECT 1.715000 1.360000 1.975000 1.620000 ;
      RECT 1.715000 1.680000 1.975000 1.940000 ;
      RECT 1.715000 2.000000 1.975000 2.260000 ;
      RECT 1.715000 2.320000 1.975000 2.580000 ;
      RECT 1.715000 6.400000 1.975000 6.660000 ;
      RECT 1.715000 6.720000 1.975000 6.980000 ;
      RECT 1.715000 7.040000 1.975000 7.300000 ;
      RECT 1.715000 7.360000 1.975000 7.620000 ;
      RECT 1.715000 7.680000 1.975000 7.940000 ;
      RECT 2.495000 2.920000 2.755000 3.180000 ;
      RECT 2.495000 3.240000 2.755000 3.500000 ;
      RECT 2.495000 3.560000 2.755000 3.820000 ;
      RECT 2.495000 3.880000 2.755000 4.140000 ;
      RECT 2.495000 4.200000 2.755000 4.460000 ;
      RECT 2.495000 4.520000 2.755000 4.780000 ;
      RECT 2.495000 4.840000 2.755000 5.100000 ;
      RECT 2.495000 5.160000 2.755000 5.420000 ;
      RECT 2.495000 5.480000 2.755000 5.740000 ;
      RECT 2.495000 5.800000 2.755000 6.060000 ;
      RECT 3.275000 1.040000 3.535000 1.300000 ;
      RECT 3.275000 1.360000 3.535000 1.620000 ;
      RECT 3.275000 1.680000 3.535000 1.940000 ;
      RECT 3.275000 2.000000 3.535000 2.260000 ;
      RECT 3.275000 2.320000 3.535000 2.580000 ;
      RECT 3.275000 6.400000 3.535000 6.660000 ;
      RECT 3.275000 6.720000 3.535000 6.980000 ;
      RECT 3.275000 7.040000 3.535000 7.300000 ;
      RECT 3.275000 7.360000 3.535000 7.620000 ;
      RECT 3.275000 7.680000 3.535000 7.940000 ;
      RECT 4.055000 2.920000 4.315000 3.180000 ;
      RECT 4.055000 3.240000 4.315000 3.500000 ;
      RECT 4.055000 3.560000 4.315000 3.820000 ;
      RECT 4.055000 3.880000 4.315000 4.140000 ;
      RECT 4.055000 4.200000 4.315000 4.460000 ;
      RECT 4.055000 4.520000 4.315000 4.780000 ;
      RECT 4.055000 4.840000 4.315000 5.100000 ;
      RECT 4.055000 5.160000 4.315000 5.420000 ;
      RECT 4.055000 5.480000 4.315000 5.740000 ;
      RECT 4.055000 5.800000 4.315000 6.060000 ;
      RECT 4.835000 1.040000 5.095000 1.300000 ;
      RECT 4.835000 1.360000 5.095000 1.620000 ;
      RECT 4.835000 1.680000 5.095000 1.940000 ;
      RECT 4.835000 2.000000 5.095000 2.260000 ;
      RECT 4.835000 2.320000 5.095000 2.580000 ;
      RECT 4.835000 6.400000 5.095000 6.660000 ;
      RECT 4.835000 6.720000 5.095000 6.980000 ;
      RECT 4.835000 7.040000 5.095000 7.300000 ;
      RECT 4.835000 7.360000 5.095000 7.620000 ;
      RECT 4.835000 7.680000 5.095000 7.940000 ;
      RECT 5.615000 2.920000 5.875000 3.180000 ;
      RECT 5.615000 3.240000 5.875000 3.500000 ;
      RECT 5.615000 3.560000 5.875000 3.820000 ;
      RECT 5.615000 3.880000 5.875000 4.140000 ;
      RECT 5.615000 4.200000 5.875000 4.460000 ;
      RECT 5.615000 4.520000 5.875000 4.780000 ;
      RECT 5.615000 4.840000 5.875000 5.100000 ;
      RECT 5.615000 5.160000 5.875000 5.420000 ;
      RECT 5.615000 5.480000 5.875000 5.740000 ;
      RECT 5.615000 5.800000 5.875000 6.060000 ;
      RECT 6.395000 1.040000 6.655000 1.300000 ;
      RECT 6.395000 1.360000 6.655000 1.620000 ;
      RECT 6.395000 1.680000 6.655000 1.940000 ;
      RECT 6.395000 2.000000 6.655000 2.260000 ;
      RECT 6.395000 2.320000 6.655000 2.580000 ;
      RECT 6.395000 6.400000 6.655000 6.660000 ;
      RECT 6.395000 6.720000 6.655000 6.980000 ;
      RECT 6.395000 7.040000 6.655000 7.300000 ;
      RECT 6.395000 7.360000 6.655000 7.620000 ;
      RECT 6.395000 7.680000 6.655000 7.940000 ;
      RECT 7.175000 2.920000 7.435000 3.180000 ;
      RECT 7.175000 3.240000 7.435000 3.500000 ;
      RECT 7.175000 3.560000 7.435000 3.820000 ;
      RECT 7.175000 3.880000 7.435000 4.140000 ;
      RECT 7.175000 4.200000 7.435000 4.460000 ;
      RECT 7.175000 4.520000 7.435000 4.780000 ;
      RECT 7.175000 4.840000 7.435000 5.100000 ;
      RECT 7.175000 5.160000 7.435000 5.420000 ;
      RECT 7.175000 5.480000 7.435000 5.740000 ;
      RECT 7.175000 5.800000 7.435000 6.060000 ;
      RECT 7.955000 1.040000 8.215000 1.300000 ;
      RECT 7.955000 1.360000 8.215000 1.620000 ;
      RECT 7.955000 1.680000 8.215000 1.940000 ;
      RECT 7.955000 2.000000 8.215000 2.260000 ;
      RECT 7.955000 2.320000 8.215000 2.580000 ;
      RECT 7.955000 6.400000 8.215000 6.660000 ;
      RECT 7.955000 6.720000 8.215000 6.980000 ;
      RECT 7.955000 7.040000 8.215000 7.300000 ;
      RECT 7.955000 7.360000 8.215000 7.620000 ;
      RECT 7.955000 7.680000 8.215000 7.940000 ;
      RECT 8.735000 2.920000 8.995000 3.180000 ;
      RECT 8.735000 3.240000 8.995000 3.500000 ;
      RECT 8.735000 3.560000 8.995000 3.820000 ;
      RECT 8.735000 3.880000 8.995000 4.140000 ;
      RECT 8.735000 4.200000 8.995000 4.460000 ;
      RECT 8.735000 4.520000 8.995000 4.780000 ;
      RECT 8.735000 4.840000 8.995000 5.100000 ;
      RECT 8.735000 5.160000 8.995000 5.420000 ;
      RECT 8.735000 5.480000 8.995000 5.740000 ;
      RECT 8.735000 5.800000 8.995000 6.060000 ;
      RECT 9.515000 1.040000 9.775000 1.300000 ;
      RECT 9.515000 1.360000 9.775000 1.620000 ;
      RECT 9.515000 1.680000 9.775000 1.940000 ;
      RECT 9.515000 2.000000 9.775000 2.260000 ;
      RECT 9.515000 2.320000 9.775000 2.580000 ;
      RECT 9.515000 6.400000 9.775000 6.660000 ;
      RECT 9.515000 6.720000 9.775000 6.980000 ;
      RECT 9.515000 7.040000 9.775000 7.300000 ;
      RECT 9.515000 7.360000 9.775000 7.620000 ;
      RECT 9.515000 7.680000 9.775000 7.940000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50
END LIBRARY
