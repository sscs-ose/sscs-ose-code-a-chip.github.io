# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4_top
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4_top ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.83000 BY  15.35000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT  0.000000  0.000000 16.830000  0.330000 ;
        RECT  0.000000  0.330000  0.330000  7.510000 ;
        RECT  0.000000  7.510000 16.830000  7.840000 ;
        RECT  0.000000  7.840000  0.330000 15.020000 ;
        RECT  0.000000 15.020000 16.830000 15.350000 ;
        RECT  1.320000  0.330000  1.710000  3.455000 ;
        RECT  1.320000  4.385000  1.710000  7.510000 ;
        RECT  1.320000  7.840000  1.710000 10.965000 ;
        RECT  1.320000 11.895000  1.710000 15.020000 ;
        RECT  2.700000  0.330000  3.090000  3.455000 ;
        RECT  2.700000  4.385000  3.090000  7.510000 ;
        RECT  2.700000  7.840000  3.090000 10.965000 ;
        RECT  2.700000 11.895000  3.090000 15.020000 ;
        RECT  4.095000  0.330000  4.485000  3.455000 ;
        RECT  4.095000  4.385000  4.485000  7.510000 ;
        RECT  4.095000  7.840000  4.485000 10.965000 ;
        RECT  4.095000 11.895000  4.485000 15.020000 ;
        RECT  5.490000  0.330000  5.880000  3.455000 ;
        RECT  5.490000  4.385000  5.880000  7.510000 ;
        RECT  5.490000  7.840000  5.880000 10.965000 ;
        RECT  5.490000 11.895000  5.880000 15.020000 ;
        RECT  6.870000  0.330000  7.260000  3.455000 ;
        RECT  6.870000  4.385000  7.260000  7.510000 ;
        RECT  6.870000  7.840000  7.260000 10.965000 ;
        RECT  6.870000 11.895000  7.260000 15.020000 ;
        RECT  8.250000  0.330000  8.580000  7.510000 ;
        RECT  8.250000  7.840000  8.580000 15.020000 ;
        RECT  9.570000  0.330000  9.960000  3.455000 ;
        RECT  9.570000  4.385000  9.960000  7.510000 ;
        RECT  9.570000  7.840000  9.960000 10.965000 ;
        RECT  9.570000 11.895000  9.960000 15.020000 ;
        RECT 10.950000  0.330000 11.340000  3.455000 ;
        RECT 10.950000  4.385000 11.340000  7.510000 ;
        RECT 10.950000  7.840000 11.340000 10.965000 ;
        RECT 10.950000 11.895000 11.340000 15.020000 ;
        RECT 12.345000  0.330000 12.735000  3.455000 ;
        RECT 12.345000  4.385000 12.735000  7.510000 ;
        RECT 12.345000  7.840000 12.735000 10.965000 ;
        RECT 12.345000 11.895000 12.735000 15.020000 ;
        RECT 13.740000  0.330000 14.130000  3.455000 ;
        RECT 13.740000  4.385000 14.130000  7.510000 ;
        RECT 13.740000  7.840000 14.130000 10.965000 ;
        RECT 13.740000 11.895000 14.130000 15.020000 ;
        RECT 15.120000  0.330000 15.510000  3.455000 ;
        RECT 15.120000  4.385000 15.510000  7.510000 ;
        RECT 15.120000  7.840000 15.510000 10.965000 ;
        RECT 15.120000 11.895000 15.510000 15.020000 ;
        RECT 16.500000  0.330000 16.830000  7.510000 ;
        RECT 16.500000  7.840000 16.830000 15.020000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT  0.630000  0.630000  1.020000  3.755000 ;
        RECT  0.630000  3.755000  7.950000  4.085000 ;
        RECT  0.630000  4.085000  1.020000  7.210000 ;
        RECT  0.630000  8.140000  1.020000 11.265000 ;
        RECT  0.630000 11.265000  7.950000 11.595000 ;
        RECT  0.630000 11.595000  1.020000 14.720000 ;
        RECT  2.010000  0.630000  2.400000  3.755000 ;
        RECT  2.010000  4.085000  2.400000  7.210000 ;
        RECT  2.010000  8.140000  2.400000 11.265000 ;
        RECT  2.010000 11.595000  2.400000 14.720000 ;
        RECT  3.390000  0.630000  3.780000  3.755000 ;
        RECT  3.390000  4.085000  3.780000  7.210000 ;
        RECT  3.390000  8.140000  3.780000 11.265000 ;
        RECT  3.390000 11.595000  3.780000 14.720000 ;
        RECT  4.800000  0.630000  5.190000  3.755000 ;
        RECT  4.800000  4.085000  5.190000  7.210000 ;
        RECT  4.800000  8.140000  5.190000 11.265000 ;
        RECT  4.800000 11.595000  5.190000 14.720000 ;
        RECT  6.180000  0.630000  6.570000  3.755000 ;
        RECT  6.180000  4.085000  6.570000  7.210000 ;
        RECT  6.180000  8.140000  6.570000 11.265000 ;
        RECT  6.180000 11.595000  6.570000 14.720000 ;
        RECT  7.560000  0.630000  7.950000  3.755000 ;
        RECT  7.560000  4.085000  7.950000  7.210000 ;
        RECT  7.560000  8.140000  7.950000 11.265000 ;
        RECT  7.560000 11.595000  7.950000 14.720000 ;
        RECT  8.880000  0.630000  9.270000  3.755000 ;
        RECT  8.880000  3.755000 16.200000  4.085000 ;
        RECT  8.880000  4.085000  9.270000  7.210000 ;
        RECT  8.880000  8.140000  9.270000 11.265000 ;
        RECT  8.880000 11.265000 16.200000 11.595000 ;
        RECT  8.880000 11.595000  9.270000 14.720000 ;
        RECT 10.260000  0.630000 10.650000  3.755000 ;
        RECT 10.260000  4.085000 10.650000  7.210000 ;
        RECT 10.260000  8.140000 10.650000 11.265000 ;
        RECT 10.260000 11.595000 10.650000 14.720000 ;
        RECT 11.640000  0.630000 12.030000  3.755000 ;
        RECT 11.640000  4.085000 12.030000  7.210000 ;
        RECT 11.640000  8.140000 12.030000 11.265000 ;
        RECT 11.640000 11.595000 12.030000 14.720000 ;
        RECT 13.050000  0.630000 13.440000  3.755000 ;
        RECT 13.050000  4.085000 13.440000  7.210000 ;
        RECT 13.050000  8.140000 13.440000 11.265000 ;
        RECT 13.050000 11.595000 13.440000 14.720000 ;
        RECT 14.430000  0.630000 14.820000  3.755000 ;
        RECT 14.430000  4.085000 14.820000  7.210000 ;
        RECT 14.430000  8.140000 14.820000 11.265000 ;
        RECT 14.430000 11.595000 14.820000 14.720000 ;
        RECT 15.810000  0.630000 16.200000  3.755000 ;
        RECT 15.810000  4.085000 16.200000  7.210000 ;
        RECT 15.810000  8.140000 16.200000 11.265000 ;
        RECT 15.810000 11.595000 16.200000 14.720000 ;
    END
  END C1
  PIN M5
    PORT
      LAYER met5 ;
        RECT 0.000000 0.000000 16.830000 15.350000 ;
    END
  END M5
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 5.895000 6.345000 5.945000 6.395000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 16.830000 15.350000 ;
    LAYER mcon ;
      RECT  0.080000  0.415000  0.250000  0.585000 ;
      RECT  0.080000  0.775000  0.250000  0.945000 ;
      RECT  0.080000  1.135000  0.250000  1.305000 ;
      RECT  0.080000  1.495000  0.250000  1.665000 ;
      RECT  0.080000  1.855000  0.250000  2.025000 ;
      RECT  0.080000  2.215000  0.250000  2.385000 ;
      RECT  0.080000  2.575000  0.250000  2.745000 ;
      RECT  0.080000  2.935000  0.250000  3.105000 ;
      RECT  0.080000  3.295000  0.250000  3.465000 ;
      RECT  0.080000  3.655000  0.250000  3.825000 ;
      RECT  0.080000  4.015000  0.250000  4.185000 ;
      RECT  0.080000  4.375000  0.250000  4.545000 ;
      RECT  0.080000  4.735000  0.250000  4.905000 ;
      RECT  0.080000  5.095000  0.250000  5.265000 ;
      RECT  0.080000  5.455000  0.250000  5.625000 ;
      RECT  0.080000  5.815000  0.250000  5.985000 ;
      RECT  0.080000  6.175000  0.250000  6.345000 ;
      RECT  0.080000  6.535000  0.250000  6.705000 ;
      RECT  0.080000  6.895000  0.250000  7.065000 ;
      RECT  0.080000  7.255000  0.250000  7.425000 ;
      RECT  0.080000  7.925000  0.250000  8.095000 ;
      RECT  0.080000  8.285000  0.250000  8.455000 ;
      RECT  0.080000  8.645000  0.250000  8.815000 ;
      RECT  0.080000  9.005000  0.250000  9.175000 ;
      RECT  0.080000  9.365000  0.250000  9.535000 ;
      RECT  0.080000  9.725000  0.250000  9.895000 ;
      RECT  0.080000 10.085000  0.250000 10.255000 ;
      RECT  0.080000 10.445000  0.250000 10.615000 ;
      RECT  0.080000 10.805000  0.250000 10.975000 ;
      RECT  0.080000 11.165000  0.250000 11.335000 ;
      RECT  0.080000 11.525000  0.250000 11.695000 ;
      RECT  0.080000 11.885000  0.250000 12.055000 ;
      RECT  0.080000 12.245000  0.250000 12.415000 ;
      RECT  0.080000 12.605000  0.250000 12.775000 ;
      RECT  0.080000 12.965000  0.250000 13.135000 ;
      RECT  0.080000 13.325000  0.250000 13.495000 ;
      RECT  0.080000 13.685000  0.250000 13.855000 ;
      RECT  0.080000 14.045000  0.250000 14.215000 ;
      RECT  0.080000 14.405000  0.250000 14.575000 ;
      RECT  0.080000 14.765000  0.250000 14.935000 ;
      RECT  0.425000  0.080000  0.595000  0.250000 ;
      RECT  0.425000  7.590000  0.595000  7.760000 ;
      RECT  0.425000 15.100000  0.595000 15.270000 ;
      RECT  0.785000  0.080000  0.955000  0.250000 ;
      RECT  0.785000  7.590000  0.955000  7.760000 ;
      RECT  0.785000 15.100000  0.955000 15.270000 ;
      RECT  1.145000  0.080000  1.315000  0.250000 ;
      RECT  1.145000  7.590000  1.315000  7.760000 ;
      RECT  1.145000 15.100000  1.315000 15.270000 ;
      RECT  1.505000  0.080000  1.675000  0.250000 ;
      RECT  1.505000  7.590000  1.675000  7.760000 ;
      RECT  1.505000 15.100000  1.675000 15.270000 ;
      RECT  1.865000  0.080000  2.035000  0.250000 ;
      RECT  1.865000  7.590000  2.035000  7.760000 ;
      RECT  1.865000 15.100000  2.035000 15.270000 ;
      RECT  2.225000  0.080000  2.395000  0.250000 ;
      RECT  2.225000  7.590000  2.395000  7.760000 ;
      RECT  2.225000 15.100000  2.395000 15.270000 ;
      RECT  2.585000  0.080000  2.755000  0.250000 ;
      RECT  2.585000  7.590000  2.755000  7.760000 ;
      RECT  2.585000 15.100000  2.755000 15.270000 ;
      RECT  2.945000  0.080000  3.115000  0.250000 ;
      RECT  2.945000  7.590000  3.115000  7.760000 ;
      RECT  2.945000 15.100000  3.115000 15.270000 ;
      RECT  3.305000  0.080000  3.475000  0.250000 ;
      RECT  3.305000  7.590000  3.475000  7.760000 ;
      RECT  3.305000 15.100000  3.475000 15.270000 ;
      RECT  3.665000  0.080000  3.835000  0.250000 ;
      RECT  3.665000  7.590000  3.835000  7.760000 ;
      RECT  3.665000 15.100000  3.835000 15.270000 ;
      RECT  4.025000  0.080000  4.195000  0.250000 ;
      RECT  4.025000  7.590000  4.195000  7.760000 ;
      RECT  4.025000 15.100000  4.195000 15.270000 ;
      RECT  4.385000  0.080000  4.555000  0.250000 ;
      RECT  4.385000  7.590000  4.555000  7.760000 ;
      RECT  4.385000 15.100000  4.555000 15.270000 ;
      RECT  4.745000  0.080000  4.915000  0.250000 ;
      RECT  4.745000  7.590000  4.915000  7.760000 ;
      RECT  4.745000 15.100000  4.915000 15.270000 ;
      RECT  5.105000  0.080000  5.275000  0.250000 ;
      RECT  5.105000  7.590000  5.275000  7.760000 ;
      RECT  5.105000 15.100000  5.275000 15.270000 ;
      RECT  5.465000  0.080000  5.635000  0.250000 ;
      RECT  5.465000  7.590000  5.635000  7.760000 ;
      RECT  5.465000 15.100000  5.635000 15.270000 ;
      RECT  5.825000  0.080000  5.995000  0.250000 ;
      RECT  5.825000  7.590000  5.995000  7.760000 ;
      RECT  5.825000 15.100000  5.995000 15.270000 ;
      RECT  6.185000  0.080000  6.355000  0.250000 ;
      RECT  6.185000  7.590000  6.355000  7.760000 ;
      RECT  6.185000 15.100000  6.355000 15.270000 ;
      RECT  6.545000  0.080000  6.715000  0.250000 ;
      RECT  6.545000  7.590000  6.715000  7.760000 ;
      RECT  6.545000 15.100000  6.715000 15.270000 ;
      RECT  6.905000  0.080000  7.075000  0.250000 ;
      RECT  6.905000  7.590000  7.075000  7.760000 ;
      RECT  6.905000 15.100000  7.075000 15.270000 ;
      RECT  7.265000  0.080000  7.435000  0.250000 ;
      RECT  7.265000  7.590000  7.435000  7.760000 ;
      RECT  7.265000 15.100000  7.435000 15.270000 ;
      RECT  7.625000  0.080000  7.795000  0.250000 ;
      RECT  7.625000  7.590000  7.795000  7.760000 ;
      RECT  7.625000 15.100000  7.795000 15.270000 ;
      RECT  7.985000  0.080000  8.155000  0.250000 ;
      RECT  7.985000  7.590000  8.155000  7.760000 ;
      RECT  7.985000 15.100000  8.155000 15.270000 ;
      RECT  8.330000  0.415000  8.500000  0.585000 ;
      RECT  8.330000  0.775000  8.500000  0.945000 ;
      RECT  8.330000  1.135000  8.500000  1.305000 ;
      RECT  8.330000  1.495000  8.500000  1.665000 ;
      RECT  8.330000  1.855000  8.500000  2.025000 ;
      RECT  8.330000  2.215000  8.500000  2.385000 ;
      RECT  8.330000  2.575000  8.500000  2.745000 ;
      RECT  8.330000  2.935000  8.500000  3.105000 ;
      RECT  8.330000  3.295000  8.500000  3.465000 ;
      RECT  8.330000  3.655000  8.500000  3.825000 ;
      RECT  8.330000  4.015000  8.500000  4.185000 ;
      RECT  8.330000  4.375000  8.500000  4.545000 ;
      RECT  8.330000  4.735000  8.500000  4.905000 ;
      RECT  8.330000  5.095000  8.500000  5.265000 ;
      RECT  8.330000  5.455000  8.500000  5.625000 ;
      RECT  8.330000  5.815000  8.500000  5.985000 ;
      RECT  8.330000  6.175000  8.500000  6.345000 ;
      RECT  8.330000  6.535000  8.500000  6.705000 ;
      RECT  8.330000  6.895000  8.500000  7.065000 ;
      RECT  8.330000  7.255000  8.500000  7.425000 ;
      RECT  8.330000  7.925000  8.500000  8.095000 ;
      RECT  8.330000  8.285000  8.500000  8.455000 ;
      RECT  8.330000  8.645000  8.500000  8.815000 ;
      RECT  8.330000  9.005000  8.500000  9.175000 ;
      RECT  8.330000  9.365000  8.500000  9.535000 ;
      RECT  8.330000  9.725000  8.500000  9.895000 ;
      RECT  8.330000 10.085000  8.500000 10.255000 ;
      RECT  8.330000 10.445000  8.500000 10.615000 ;
      RECT  8.330000 10.805000  8.500000 10.975000 ;
      RECT  8.330000 11.165000  8.500000 11.335000 ;
      RECT  8.330000 11.525000  8.500000 11.695000 ;
      RECT  8.330000 11.885000  8.500000 12.055000 ;
      RECT  8.330000 12.245000  8.500000 12.415000 ;
      RECT  8.330000 12.605000  8.500000 12.775000 ;
      RECT  8.330000 12.965000  8.500000 13.135000 ;
      RECT  8.330000 13.325000  8.500000 13.495000 ;
      RECT  8.330000 13.685000  8.500000 13.855000 ;
      RECT  8.330000 14.045000  8.500000 14.215000 ;
      RECT  8.330000 14.405000  8.500000 14.575000 ;
      RECT  8.330000 14.765000  8.500000 14.935000 ;
      RECT  8.675000  0.080000  8.845000  0.250000 ;
      RECT  8.675000  7.590000  8.845000  7.760000 ;
      RECT  8.675000 15.100000  8.845000 15.270000 ;
      RECT  9.035000  0.080000  9.205000  0.250000 ;
      RECT  9.035000  7.590000  9.205000  7.760000 ;
      RECT  9.035000 15.100000  9.205000 15.270000 ;
      RECT  9.395000  0.080000  9.565000  0.250000 ;
      RECT  9.395000  7.590000  9.565000  7.760000 ;
      RECT  9.395000 15.100000  9.565000 15.270000 ;
      RECT  9.755000  0.080000  9.925000  0.250000 ;
      RECT  9.755000  7.590000  9.925000  7.760000 ;
      RECT  9.755000 15.100000  9.925000 15.270000 ;
      RECT 10.115000  0.080000 10.285000  0.250000 ;
      RECT 10.115000  7.590000 10.285000  7.760000 ;
      RECT 10.115000 15.100000 10.285000 15.270000 ;
      RECT 10.475000  0.080000 10.645000  0.250000 ;
      RECT 10.475000  7.590000 10.645000  7.760000 ;
      RECT 10.475000 15.100000 10.645000 15.270000 ;
      RECT 10.835000  0.080000 11.005000  0.250000 ;
      RECT 10.835000  7.590000 11.005000  7.760000 ;
      RECT 10.835000 15.100000 11.005000 15.270000 ;
      RECT 11.195000  0.080000 11.365000  0.250000 ;
      RECT 11.195000  7.590000 11.365000  7.760000 ;
      RECT 11.195000 15.100000 11.365000 15.270000 ;
      RECT 11.555000  0.080000 11.725000  0.250000 ;
      RECT 11.555000  7.590000 11.725000  7.760000 ;
      RECT 11.555000 15.100000 11.725000 15.270000 ;
      RECT 11.915000  0.080000 12.085000  0.250000 ;
      RECT 11.915000  7.590000 12.085000  7.760000 ;
      RECT 11.915000 15.100000 12.085000 15.270000 ;
      RECT 12.275000  0.080000 12.445000  0.250000 ;
      RECT 12.275000  7.590000 12.445000  7.760000 ;
      RECT 12.275000 15.100000 12.445000 15.270000 ;
      RECT 12.635000  0.080000 12.805000  0.250000 ;
      RECT 12.635000  7.590000 12.805000  7.760000 ;
      RECT 12.635000 15.100000 12.805000 15.270000 ;
      RECT 12.995000  0.080000 13.165000  0.250000 ;
      RECT 12.995000  7.590000 13.165000  7.760000 ;
      RECT 12.995000 15.100000 13.165000 15.270000 ;
      RECT 13.355000  0.080000 13.525000  0.250000 ;
      RECT 13.355000  7.590000 13.525000  7.760000 ;
      RECT 13.355000 15.100000 13.525000 15.270000 ;
      RECT 13.715000  0.080000 13.885000  0.250000 ;
      RECT 13.715000  7.590000 13.885000  7.760000 ;
      RECT 13.715000 15.100000 13.885000 15.270000 ;
      RECT 14.075000  0.080000 14.245000  0.250000 ;
      RECT 14.075000  7.590000 14.245000  7.760000 ;
      RECT 14.075000 15.100000 14.245000 15.270000 ;
      RECT 14.435000  0.080000 14.605000  0.250000 ;
      RECT 14.435000  7.590000 14.605000  7.760000 ;
      RECT 14.435000 15.100000 14.605000 15.270000 ;
      RECT 14.795000  0.080000 14.965000  0.250000 ;
      RECT 14.795000  7.590000 14.965000  7.760000 ;
      RECT 14.795000 15.100000 14.965000 15.270000 ;
      RECT 15.155000  0.080000 15.325000  0.250000 ;
      RECT 15.155000  7.590000 15.325000  7.760000 ;
      RECT 15.155000 15.100000 15.325000 15.270000 ;
      RECT 15.515000  0.080000 15.685000  0.250000 ;
      RECT 15.515000  7.590000 15.685000  7.760000 ;
      RECT 15.515000 15.100000 15.685000 15.270000 ;
      RECT 15.875000  0.080000 16.045000  0.250000 ;
      RECT 15.875000  7.590000 16.045000  7.760000 ;
      RECT 15.875000 15.100000 16.045000 15.270000 ;
      RECT 16.235000  0.080000 16.405000  0.250000 ;
      RECT 16.235000  7.590000 16.405000  7.760000 ;
      RECT 16.235000 15.100000 16.405000 15.270000 ;
      RECT 16.580000  0.415000 16.750000  0.585000 ;
      RECT 16.580000  0.775000 16.750000  0.945000 ;
      RECT 16.580000  1.135000 16.750000  1.305000 ;
      RECT 16.580000  1.495000 16.750000  1.665000 ;
      RECT 16.580000  1.855000 16.750000  2.025000 ;
      RECT 16.580000  2.215000 16.750000  2.385000 ;
      RECT 16.580000  2.575000 16.750000  2.745000 ;
      RECT 16.580000  2.935000 16.750000  3.105000 ;
      RECT 16.580000  3.295000 16.750000  3.465000 ;
      RECT 16.580000  3.655000 16.750000  3.825000 ;
      RECT 16.580000  4.015000 16.750000  4.185000 ;
      RECT 16.580000  4.375000 16.750000  4.545000 ;
      RECT 16.580000  4.735000 16.750000  4.905000 ;
      RECT 16.580000  5.095000 16.750000  5.265000 ;
      RECT 16.580000  5.455000 16.750000  5.625000 ;
      RECT 16.580000  5.815000 16.750000  5.985000 ;
      RECT 16.580000  6.175000 16.750000  6.345000 ;
      RECT 16.580000  6.535000 16.750000  6.705000 ;
      RECT 16.580000  6.895000 16.750000  7.065000 ;
      RECT 16.580000  7.255000 16.750000  7.425000 ;
      RECT 16.580000  7.925000 16.750000  8.095000 ;
      RECT 16.580000  8.285000 16.750000  8.455000 ;
      RECT 16.580000  8.645000 16.750000  8.815000 ;
      RECT 16.580000  9.005000 16.750000  9.175000 ;
      RECT 16.580000  9.365000 16.750000  9.535000 ;
      RECT 16.580000  9.725000 16.750000  9.895000 ;
      RECT 16.580000 10.085000 16.750000 10.255000 ;
      RECT 16.580000 10.445000 16.750000 10.615000 ;
      RECT 16.580000 10.805000 16.750000 10.975000 ;
      RECT 16.580000 11.165000 16.750000 11.335000 ;
      RECT 16.580000 11.525000 16.750000 11.695000 ;
      RECT 16.580000 11.885000 16.750000 12.055000 ;
      RECT 16.580000 12.245000 16.750000 12.415000 ;
      RECT 16.580000 12.605000 16.750000 12.775000 ;
      RECT 16.580000 12.965000 16.750000 13.135000 ;
      RECT 16.580000 13.325000 16.750000 13.495000 ;
      RECT 16.580000 13.685000 16.750000 13.855000 ;
      RECT 16.580000 14.045000 16.750000 14.215000 ;
      RECT 16.580000 14.405000 16.750000 14.575000 ;
      RECT 16.580000 14.765000 16.750000 14.935000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 16.830000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  7.510000 ;
      RECT  0.000000  7.510000 16.830000  7.840000 ;
      RECT  0.000000  7.840000  0.330000 15.020000 ;
      RECT  0.000000 15.020000 16.830000 15.350000 ;
      RECT  0.495000  0.470000  0.635000  3.760000 ;
      RECT  0.495000  3.760000  8.085000  4.080000 ;
      RECT  0.495000  4.080000  0.635000  7.370000 ;
      RECT  0.495000  7.980000  0.635000 11.270000 ;
      RECT  0.495000 11.270000  8.085000 11.590000 ;
      RECT  0.495000 11.590000  0.635000 14.880000 ;
      RECT  0.775000  0.330000  0.915000  3.620000 ;
      RECT  0.775000  4.220000  0.915000  7.510000 ;
      RECT  0.775000  7.840000  0.915000 11.130000 ;
      RECT  0.775000 11.730000  0.915000 15.020000 ;
      RECT  1.055000  0.470000  1.195000  3.760000 ;
      RECT  1.055000  4.080000  1.195000  7.370000 ;
      RECT  1.055000  7.980000  1.195000 11.270000 ;
      RECT  1.055000 11.590000  1.195000 14.880000 ;
      RECT  1.335000  0.330000  1.475000  3.620000 ;
      RECT  1.335000  4.220000  1.475000  7.510000 ;
      RECT  1.335000  7.840000  1.475000 11.130000 ;
      RECT  1.335000 11.730000  1.475000 15.020000 ;
      RECT  1.615000  0.470000  1.755000  3.760000 ;
      RECT  1.615000  4.080000  1.755000  7.370000 ;
      RECT  1.615000  7.980000  1.755000 11.270000 ;
      RECT  1.615000 11.590000  1.755000 14.880000 ;
      RECT  1.895000  0.330000  2.035000  3.620000 ;
      RECT  1.895000  4.220000  2.035000  7.510000 ;
      RECT  1.895000  7.840000  2.035000 11.130000 ;
      RECT  1.895000 11.730000  2.035000 15.020000 ;
      RECT  2.175000  0.470000  2.315000  3.760000 ;
      RECT  2.175000  4.080000  2.315000  7.370000 ;
      RECT  2.175000  7.980000  2.315000 11.270000 ;
      RECT  2.175000 11.590000  2.315000 14.880000 ;
      RECT  2.455000  0.330000  2.595000  3.620000 ;
      RECT  2.455000  4.220000  2.595000  7.510000 ;
      RECT  2.455000  7.840000  2.595000 11.130000 ;
      RECT  2.455000 11.730000  2.595000 15.020000 ;
      RECT  2.735000  0.470000  2.875000  3.760000 ;
      RECT  2.735000  4.080000  2.875000  7.370000 ;
      RECT  2.735000  7.980000  2.875000 11.270000 ;
      RECT  2.735000 11.590000  2.875000 14.880000 ;
      RECT  3.015000  0.330000  3.155000  3.620000 ;
      RECT  3.015000  4.220000  3.155000  7.510000 ;
      RECT  3.015000  7.840000  3.155000 11.130000 ;
      RECT  3.015000 11.730000  3.155000 15.020000 ;
      RECT  3.295000  0.470000  3.435000  3.760000 ;
      RECT  3.295000  4.080000  3.435000  7.370000 ;
      RECT  3.295000  7.980000  3.435000 11.270000 ;
      RECT  3.295000 11.590000  3.435000 14.880000 ;
      RECT  3.575000  0.330000  3.715000  3.620000 ;
      RECT  3.575000  4.220000  3.715000  7.510000 ;
      RECT  3.575000  7.840000  3.715000 11.130000 ;
      RECT  3.575000 11.730000  3.715000 15.020000 ;
      RECT  3.855000  0.470000  3.995000  3.760000 ;
      RECT  3.855000  4.080000  3.995000  7.370000 ;
      RECT  3.855000  7.980000  3.995000 11.270000 ;
      RECT  3.855000 11.590000  3.995000 14.880000 ;
      RECT  4.155000  0.470000  4.425000  3.760000 ;
      RECT  4.155000  4.080000  4.425000  7.370000 ;
      RECT  4.155000  7.980000  4.425000 11.270000 ;
      RECT  4.155000 11.590000  4.425000 14.880000 ;
      RECT  4.585000  0.470000  4.725000  3.760000 ;
      RECT  4.585000  4.080000  4.725000  7.370000 ;
      RECT  4.585000  7.980000  4.725000 11.270000 ;
      RECT  4.585000 11.590000  4.725000 14.880000 ;
      RECT  4.865000  0.330000  5.005000  3.620000 ;
      RECT  4.865000  4.220000  5.005000  7.510000 ;
      RECT  4.865000  7.840000  5.005000 11.130000 ;
      RECT  4.865000 11.730000  5.005000 15.020000 ;
      RECT  5.145000  0.470000  5.285000  3.760000 ;
      RECT  5.145000  4.080000  5.285000  7.370000 ;
      RECT  5.145000  7.980000  5.285000 11.270000 ;
      RECT  5.145000 11.590000  5.285000 14.880000 ;
      RECT  5.425000  0.330000  5.565000  3.620000 ;
      RECT  5.425000  4.220000  5.565000  7.510000 ;
      RECT  5.425000  7.840000  5.565000 11.130000 ;
      RECT  5.425000 11.730000  5.565000 15.020000 ;
      RECT  5.705000  0.470000  5.845000  3.760000 ;
      RECT  5.705000  4.080000  5.845000  7.370000 ;
      RECT  5.705000  7.980000  5.845000 11.270000 ;
      RECT  5.705000 11.590000  5.845000 14.880000 ;
      RECT  5.985000  0.330000  6.125000  3.620000 ;
      RECT  5.985000  4.220000  6.125000  7.510000 ;
      RECT  5.985000  7.840000  6.125000 11.130000 ;
      RECT  5.985000 11.730000  6.125000 15.020000 ;
      RECT  6.265000  0.470000  6.405000  3.760000 ;
      RECT  6.265000  4.080000  6.405000  7.370000 ;
      RECT  6.265000  7.980000  6.405000 11.270000 ;
      RECT  6.265000 11.590000  6.405000 14.880000 ;
      RECT  6.545000  0.330000  6.685000  3.620000 ;
      RECT  6.545000  4.220000  6.685000  7.510000 ;
      RECT  6.545000  7.840000  6.685000 11.130000 ;
      RECT  6.545000 11.730000  6.685000 15.020000 ;
      RECT  6.825000  0.470000  6.965000  3.760000 ;
      RECT  6.825000  4.080000  6.965000  7.370000 ;
      RECT  6.825000  7.980000  6.965000 11.270000 ;
      RECT  6.825000 11.590000  6.965000 14.880000 ;
      RECT  7.105000  0.330000  7.245000  3.620000 ;
      RECT  7.105000  4.220000  7.245000  7.510000 ;
      RECT  7.105000  7.840000  7.245000 11.130000 ;
      RECT  7.105000 11.730000  7.245000 15.020000 ;
      RECT  7.385000  0.470000  7.525000  3.760000 ;
      RECT  7.385000  4.080000  7.525000  7.370000 ;
      RECT  7.385000  7.980000  7.525000 11.270000 ;
      RECT  7.385000 11.590000  7.525000 14.880000 ;
      RECT  7.665000  0.330000  7.805000  3.620000 ;
      RECT  7.665000  4.220000  7.805000  7.510000 ;
      RECT  7.665000  7.840000  7.805000 11.130000 ;
      RECT  7.665000 11.730000  7.805000 15.020000 ;
      RECT  7.945000  0.470000  8.085000  3.760000 ;
      RECT  7.945000  4.080000  8.085000  7.370000 ;
      RECT  7.945000  7.980000  8.085000 11.270000 ;
      RECT  7.945000 11.590000  8.085000 14.880000 ;
      RECT  8.250000  0.330000  8.580000  7.510000 ;
      RECT  8.250000  7.840000  8.580000 15.020000 ;
      RECT  8.745000  0.470000  8.885000  3.760000 ;
      RECT  8.745000  3.760000 16.335000  4.080000 ;
      RECT  8.745000  4.080000  8.885000  7.370000 ;
      RECT  8.745000  7.980000  8.885000 11.270000 ;
      RECT  8.745000 11.270000 16.335000 11.590000 ;
      RECT  8.745000 11.590000  8.885000 14.880000 ;
      RECT  9.025000  0.330000  9.165000  3.620000 ;
      RECT  9.025000  4.220000  9.165000  7.510000 ;
      RECT  9.025000  7.840000  9.165000 11.130000 ;
      RECT  9.025000 11.730000  9.165000 15.020000 ;
      RECT  9.305000  0.470000  9.445000  3.760000 ;
      RECT  9.305000  4.080000  9.445000  7.370000 ;
      RECT  9.305000  7.980000  9.445000 11.270000 ;
      RECT  9.305000 11.590000  9.445000 14.880000 ;
      RECT  9.585000  0.330000  9.725000  3.620000 ;
      RECT  9.585000  4.220000  9.725000  7.510000 ;
      RECT  9.585000  7.840000  9.725000 11.130000 ;
      RECT  9.585000 11.730000  9.725000 15.020000 ;
      RECT  9.865000  0.470000 10.005000  3.760000 ;
      RECT  9.865000  4.080000 10.005000  7.370000 ;
      RECT  9.865000  7.980000 10.005000 11.270000 ;
      RECT  9.865000 11.590000 10.005000 14.880000 ;
      RECT 10.145000  0.330000 10.285000  3.620000 ;
      RECT 10.145000  4.220000 10.285000  7.510000 ;
      RECT 10.145000  7.840000 10.285000 11.130000 ;
      RECT 10.145000 11.730000 10.285000 15.020000 ;
      RECT 10.425000  0.470000 10.565000  3.760000 ;
      RECT 10.425000  4.080000 10.565000  7.370000 ;
      RECT 10.425000  7.980000 10.565000 11.270000 ;
      RECT 10.425000 11.590000 10.565000 14.880000 ;
      RECT 10.705000  0.330000 10.845000  3.620000 ;
      RECT 10.705000  4.220000 10.845000  7.510000 ;
      RECT 10.705000  7.840000 10.845000 11.130000 ;
      RECT 10.705000 11.730000 10.845000 15.020000 ;
      RECT 10.985000  0.470000 11.125000  3.760000 ;
      RECT 10.985000  4.080000 11.125000  7.370000 ;
      RECT 10.985000  7.980000 11.125000 11.270000 ;
      RECT 10.985000 11.590000 11.125000 14.880000 ;
      RECT 11.265000  0.330000 11.405000  3.620000 ;
      RECT 11.265000  4.220000 11.405000  7.510000 ;
      RECT 11.265000  7.840000 11.405000 11.130000 ;
      RECT 11.265000 11.730000 11.405000 15.020000 ;
      RECT 11.545000  0.470000 11.685000  3.760000 ;
      RECT 11.545000  4.080000 11.685000  7.370000 ;
      RECT 11.545000  7.980000 11.685000 11.270000 ;
      RECT 11.545000 11.590000 11.685000 14.880000 ;
      RECT 11.825000  0.330000 11.965000  3.620000 ;
      RECT 11.825000  4.220000 11.965000  7.510000 ;
      RECT 11.825000  7.840000 11.965000 11.130000 ;
      RECT 11.825000 11.730000 11.965000 15.020000 ;
      RECT 12.105000  0.470000 12.245000  3.760000 ;
      RECT 12.105000  4.080000 12.245000  7.370000 ;
      RECT 12.105000  7.980000 12.245000 11.270000 ;
      RECT 12.105000 11.590000 12.245000 14.880000 ;
      RECT 12.405000  0.470000 12.675000  3.760000 ;
      RECT 12.405000  4.080000 12.675000  7.370000 ;
      RECT 12.405000  7.980000 12.675000 11.270000 ;
      RECT 12.405000 11.590000 12.675000 14.880000 ;
      RECT 12.835000  0.470000 12.975000  3.760000 ;
      RECT 12.835000  4.080000 12.975000  7.370000 ;
      RECT 12.835000  7.980000 12.975000 11.270000 ;
      RECT 12.835000 11.590000 12.975000 14.880000 ;
      RECT 13.115000  0.330000 13.255000  3.620000 ;
      RECT 13.115000  4.220000 13.255000  7.510000 ;
      RECT 13.115000  7.840000 13.255000 11.130000 ;
      RECT 13.115000 11.730000 13.255000 15.020000 ;
      RECT 13.395000  0.470000 13.535000  3.760000 ;
      RECT 13.395000  4.080000 13.535000  7.370000 ;
      RECT 13.395000  7.980000 13.535000 11.270000 ;
      RECT 13.395000 11.590000 13.535000 14.880000 ;
      RECT 13.675000  0.330000 13.815000  3.620000 ;
      RECT 13.675000  4.220000 13.815000  7.510000 ;
      RECT 13.675000  7.840000 13.815000 11.130000 ;
      RECT 13.675000 11.730000 13.815000 15.020000 ;
      RECT 13.955000  0.470000 14.095000  3.760000 ;
      RECT 13.955000  4.080000 14.095000  7.370000 ;
      RECT 13.955000  7.980000 14.095000 11.270000 ;
      RECT 13.955000 11.590000 14.095000 14.880000 ;
      RECT 14.235000  0.330000 14.375000  3.620000 ;
      RECT 14.235000  4.220000 14.375000  7.510000 ;
      RECT 14.235000  7.840000 14.375000 11.130000 ;
      RECT 14.235000 11.730000 14.375000 15.020000 ;
      RECT 14.515000  0.470000 14.655000  3.760000 ;
      RECT 14.515000  4.080000 14.655000  7.370000 ;
      RECT 14.515000  7.980000 14.655000 11.270000 ;
      RECT 14.515000 11.590000 14.655000 14.880000 ;
      RECT 14.795000  0.330000 14.935000  3.620000 ;
      RECT 14.795000  4.220000 14.935000  7.510000 ;
      RECT 14.795000  7.840000 14.935000 11.130000 ;
      RECT 14.795000 11.730000 14.935000 15.020000 ;
      RECT 15.075000  0.470000 15.215000  3.760000 ;
      RECT 15.075000  4.080000 15.215000  7.370000 ;
      RECT 15.075000  7.980000 15.215000 11.270000 ;
      RECT 15.075000 11.590000 15.215000 14.880000 ;
      RECT 15.355000  0.330000 15.495000  3.620000 ;
      RECT 15.355000  4.220000 15.495000  7.510000 ;
      RECT 15.355000  7.840000 15.495000 11.130000 ;
      RECT 15.355000 11.730000 15.495000 15.020000 ;
      RECT 15.635000  0.470000 15.775000  3.760000 ;
      RECT 15.635000  4.080000 15.775000  7.370000 ;
      RECT 15.635000  7.980000 15.775000 11.270000 ;
      RECT 15.635000 11.590000 15.775000 14.880000 ;
      RECT 15.915000  0.330000 16.055000  3.620000 ;
      RECT 15.915000  4.220000 16.055000  7.510000 ;
      RECT 15.915000  7.840000 16.055000 11.130000 ;
      RECT 15.915000 11.730000 16.055000 15.020000 ;
      RECT 16.195000  0.470000 16.335000  3.760000 ;
      RECT 16.195000  4.080000 16.335000  7.370000 ;
      RECT 16.195000  7.980000 16.335000 11.270000 ;
      RECT 16.195000 11.590000 16.335000 14.880000 ;
      RECT 16.500000  0.330000 16.830000  7.510000 ;
      RECT 16.500000  7.840000 16.830000 15.020000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  4.015000  0.330000 ;
      RECT  0.000000  0.330000  0.330000  0.750000 ;
      RECT  0.000000  0.750000  4.010000  0.890000 ;
      RECT  0.000000  0.890000  0.330000  1.310000 ;
      RECT  0.000000  1.310000  4.010000  1.450000 ;
      RECT  0.000000  1.450000  0.330000  1.870000 ;
      RECT  0.000000  1.870000  4.010000  2.010000 ;
      RECT  0.000000  2.010000  0.330000  2.430000 ;
      RECT  0.000000  2.430000  4.010000  2.570000 ;
      RECT  0.000000  2.570000  0.330000  2.990000 ;
      RECT  0.000000  2.990000  4.010000  3.130000 ;
      RECT  0.000000  3.130000  0.330000  3.645000 ;
      RECT  0.000000  3.785000 16.830000  4.055000 ;
      RECT  0.000000  4.195000  0.330000  4.710000 ;
      RECT  0.000000  4.710000  4.010000  4.850000 ;
      RECT  0.000000  4.850000  0.330000  5.270000 ;
      RECT  0.000000  5.270000  4.010000  5.410000 ;
      RECT  0.000000  5.410000  0.330000  5.830000 ;
      RECT  0.000000  5.830000  4.010000  5.970000 ;
      RECT  0.000000  5.970000  0.330000  6.390000 ;
      RECT  0.000000  6.390000  4.010000  6.530000 ;
      RECT  0.000000  6.530000  0.330000  6.950000 ;
      RECT  0.000000  6.950000  4.010000  7.090000 ;
      RECT  0.000000  7.090000  0.330000  7.510000 ;
      RECT  0.000000  7.510000  4.015000  7.840000 ;
      RECT  0.000000  7.840000  0.330000  8.260000 ;
      RECT  0.000000  8.260000  4.010000  8.400000 ;
      RECT  0.000000  8.400000  0.330000  8.820000 ;
      RECT  0.000000  8.820000  4.010000  8.960000 ;
      RECT  0.000000  8.960000  0.330000  9.380000 ;
      RECT  0.000000  9.380000  4.010000  9.520000 ;
      RECT  0.000000  9.520000  0.330000  9.940000 ;
      RECT  0.000000  9.940000  4.010000 10.080000 ;
      RECT  0.000000 10.080000  0.330000 10.500000 ;
      RECT  0.000000 10.500000  4.010000 10.640000 ;
      RECT  0.000000 10.640000  0.330000 11.155000 ;
      RECT  0.000000 11.295000 16.830000 11.565000 ;
      RECT  0.000000 11.705000  0.330000 12.220000 ;
      RECT  0.000000 12.220000  4.010000 12.360000 ;
      RECT  0.000000 12.360000  0.330000 12.780000 ;
      RECT  0.000000 12.780000  4.010000 12.920000 ;
      RECT  0.000000 12.920000  0.330000 13.340000 ;
      RECT  0.000000 13.340000  4.010000 13.480000 ;
      RECT  0.000000 13.480000  0.330000 13.900000 ;
      RECT  0.000000 13.900000  4.010000 14.040000 ;
      RECT  0.000000 14.040000  0.330000 14.460000 ;
      RECT  0.000000 14.460000  4.010000 14.600000 ;
      RECT  0.000000 14.600000  0.330000 15.020000 ;
      RECT  0.000000 15.020000  4.015000 15.350000 ;
      RECT  0.370000  3.780000  8.210000  3.785000 ;
      RECT  0.370000  4.055000  8.210000  4.060000 ;
      RECT  0.370000 11.290000  8.210000 11.295000 ;
      RECT  0.370000 11.565000  8.210000 11.570000 ;
      RECT  0.470000  0.470000  8.110000  0.610000 ;
      RECT  0.470000  1.030000  8.110000  1.170000 ;
      RECT  0.470000  1.590000  8.110000  1.730000 ;
      RECT  0.470000  2.150000  8.110000  2.290000 ;
      RECT  0.470000  2.710000  8.110000  2.850000 ;
      RECT  0.470000  3.270000  8.110000  3.640000 ;
      RECT  0.470000  4.200000  8.110000  4.570000 ;
      RECT  0.470000  4.990000  8.110000  5.130000 ;
      RECT  0.470000  5.550000  8.110000  5.690000 ;
      RECT  0.470000  6.110000  8.110000  6.250000 ;
      RECT  0.470000  6.670000  8.110000  6.810000 ;
      RECT  0.470000  7.230000  8.110000  7.370000 ;
      RECT  0.470000  7.980000  8.110000  8.120000 ;
      RECT  0.470000  8.540000  8.110000  8.680000 ;
      RECT  0.470000  9.100000  8.110000  9.240000 ;
      RECT  0.470000  9.660000  8.110000  9.800000 ;
      RECT  0.470000 10.220000  8.110000 10.360000 ;
      RECT  0.470000 10.780000  8.110000 11.150000 ;
      RECT  0.470000 11.710000  8.110000 12.080000 ;
      RECT  0.470000 12.500000  8.110000 12.640000 ;
      RECT  0.470000 13.060000  8.110000 13.200000 ;
      RECT  0.470000 13.620000  8.110000 13.760000 ;
      RECT  0.470000 14.180000  8.110000 14.320000 ;
      RECT  0.470000 14.740000  8.110000 14.880000 ;
      RECT  4.150000  0.610000  4.430000  1.030000 ;
      RECT  4.150000  1.170000  4.430000  1.590000 ;
      RECT  4.150000  1.730000  4.430000  2.150000 ;
      RECT  4.150000  2.290000  4.430000  2.710000 ;
      RECT  4.150000  2.850000  4.430000  3.270000 ;
      RECT  4.150000  3.640000  4.430000  3.780000 ;
      RECT  4.150000  4.060000  4.430000  4.200000 ;
      RECT  4.150000  4.570000  4.430000  4.990000 ;
      RECT  4.150000  5.130000  4.430000  5.550000 ;
      RECT  4.150000  5.690000  4.430000  6.110000 ;
      RECT  4.150000  6.250000  4.430000  6.670000 ;
      RECT  4.150000  6.810000  4.430000  7.230000 ;
      RECT  4.150000  8.120000  4.430000  8.540000 ;
      RECT  4.150000  8.680000  4.430000  9.100000 ;
      RECT  4.150000  9.240000  4.430000  9.660000 ;
      RECT  4.150000  9.800000  4.430000 10.220000 ;
      RECT  4.150000 10.360000  4.430000 10.780000 ;
      RECT  4.150000 11.150000  4.430000 11.290000 ;
      RECT  4.150000 11.570000  4.430000 11.710000 ;
      RECT  4.150000 12.080000  4.430000 12.500000 ;
      RECT  4.150000 12.640000  4.430000 13.060000 ;
      RECT  4.150000 13.200000  4.430000 13.620000 ;
      RECT  4.150000 13.760000  4.430000 14.180000 ;
      RECT  4.150000 14.320000  4.430000 14.740000 ;
      RECT  4.155000  0.000000  4.425000  0.470000 ;
      RECT  4.155000  7.370000  4.425000  7.980000 ;
      RECT  4.155000 14.880000  4.425000 15.350000 ;
      RECT  4.565000  0.000000 12.265000  0.330000 ;
      RECT  4.565000  7.510000 12.265000  7.840000 ;
      RECT  4.565000 15.020000 12.265000 15.350000 ;
      RECT  4.570000  0.750000 12.260000  0.890000 ;
      RECT  4.570000  1.310000 12.260000  1.450000 ;
      RECT  4.570000  1.870000 12.260000  2.010000 ;
      RECT  4.570000  2.430000 12.260000  2.570000 ;
      RECT  4.570000  2.990000 12.260000  3.130000 ;
      RECT  4.570000  4.710000 12.260000  4.850000 ;
      RECT  4.570000  5.270000 12.260000  5.410000 ;
      RECT  4.570000  5.830000 12.260000  5.970000 ;
      RECT  4.570000  6.390000 12.260000  6.530000 ;
      RECT  4.570000  6.950000 12.260000  7.090000 ;
      RECT  4.570000  8.260000 12.260000  8.400000 ;
      RECT  4.570000  8.820000 12.260000  8.960000 ;
      RECT  4.570000  9.380000 12.260000  9.520000 ;
      RECT  4.570000  9.940000 12.260000 10.080000 ;
      RECT  4.570000 10.500000 12.260000 10.640000 ;
      RECT  4.570000 12.220000 12.260000 12.360000 ;
      RECT  4.570000 12.780000 12.260000 12.920000 ;
      RECT  4.570000 13.340000 12.260000 13.480000 ;
      RECT  4.570000 13.900000 12.260000 14.040000 ;
      RECT  4.570000 14.460000 12.260000 14.600000 ;
      RECT  8.250000  0.330000  8.580000  0.750000 ;
      RECT  8.250000  0.890000  8.580000  1.310000 ;
      RECT  8.250000  1.450000  8.580000  1.870000 ;
      RECT  8.250000  2.010000  8.580000  2.430000 ;
      RECT  8.250000  2.570000  8.580000  2.990000 ;
      RECT  8.250000  3.130000  8.580000  3.645000 ;
      RECT  8.250000  4.195000  8.580000  4.710000 ;
      RECT  8.250000  4.850000  8.580000  5.270000 ;
      RECT  8.250000  5.410000  8.580000  5.830000 ;
      RECT  8.250000  5.970000  8.580000  6.390000 ;
      RECT  8.250000  6.530000  8.580000  6.950000 ;
      RECT  8.250000  7.090000  8.580000  7.510000 ;
      RECT  8.250000  7.840000  8.580000  8.260000 ;
      RECT  8.250000  8.400000  8.580000  8.820000 ;
      RECT  8.250000  8.960000  8.580000  9.380000 ;
      RECT  8.250000  9.520000  8.580000  9.940000 ;
      RECT  8.250000 10.080000  8.580000 10.500000 ;
      RECT  8.250000 10.640000  8.580000 11.155000 ;
      RECT  8.250000 11.705000  8.580000 12.220000 ;
      RECT  8.250000 12.360000  8.580000 12.780000 ;
      RECT  8.250000 12.920000  8.580000 13.340000 ;
      RECT  8.250000 13.480000  8.580000 13.900000 ;
      RECT  8.250000 14.040000  8.580000 14.460000 ;
      RECT  8.250000 14.600000  8.580000 15.020000 ;
      RECT  8.620000  3.780000 16.460000  3.785000 ;
      RECT  8.620000  4.055000 16.460000  4.060000 ;
      RECT  8.620000 11.290000 16.460000 11.295000 ;
      RECT  8.620000 11.565000 16.460000 11.570000 ;
      RECT  8.720000  0.470000 16.360000  0.610000 ;
      RECT  8.720000  1.030000 16.360000  1.170000 ;
      RECT  8.720000  1.590000 16.360000  1.730000 ;
      RECT  8.720000  2.150000 16.360000  2.290000 ;
      RECT  8.720000  2.710000 16.360000  2.850000 ;
      RECT  8.720000  3.270000 16.360000  3.640000 ;
      RECT  8.720000  4.200000 16.360000  4.570000 ;
      RECT  8.720000  4.990000 16.360000  5.130000 ;
      RECT  8.720000  5.550000 16.360000  5.690000 ;
      RECT  8.720000  6.110000 16.360000  6.250000 ;
      RECT  8.720000  6.670000 16.360000  6.810000 ;
      RECT  8.720000  7.230000 16.360000  7.370000 ;
      RECT  8.720000  7.980000 16.360000  8.120000 ;
      RECT  8.720000  8.540000 16.360000  8.680000 ;
      RECT  8.720000  9.100000 16.360000  9.240000 ;
      RECT  8.720000  9.660000 16.360000  9.800000 ;
      RECT  8.720000 10.220000 16.360000 10.360000 ;
      RECT  8.720000 10.780000 16.360000 11.150000 ;
      RECT  8.720000 11.710000 16.360000 12.080000 ;
      RECT  8.720000 12.500000 16.360000 12.640000 ;
      RECT  8.720000 13.060000 16.360000 13.200000 ;
      RECT  8.720000 13.620000 16.360000 13.760000 ;
      RECT  8.720000 14.180000 16.360000 14.320000 ;
      RECT  8.720000 14.740000 16.360000 14.880000 ;
      RECT 12.400000  0.610000 12.680000  1.030000 ;
      RECT 12.400000  1.170000 12.680000  1.590000 ;
      RECT 12.400000  1.730000 12.680000  2.150000 ;
      RECT 12.400000  2.290000 12.680000  2.710000 ;
      RECT 12.400000  2.850000 12.680000  3.270000 ;
      RECT 12.400000  3.640000 12.680000  3.780000 ;
      RECT 12.400000  4.060000 12.680000  4.200000 ;
      RECT 12.400000  4.570000 12.680000  4.990000 ;
      RECT 12.400000  5.130000 12.680000  5.550000 ;
      RECT 12.400000  5.690000 12.680000  6.110000 ;
      RECT 12.400000  6.250000 12.680000  6.670000 ;
      RECT 12.400000  6.810000 12.680000  7.230000 ;
      RECT 12.400000  8.120000 12.680000  8.540000 ;
      RECT 12.400000  8.680000 12.680000  9.100000 ;
      RECT 12.400000  9.240000 12.680000  9.660000 ;
      RECT 12.400000  9.800000 12.680000 10.220000 ;
      RECT 12.400000 10.360000 12.680000 10.780000 ;
      RECT 12.400000 11.150000 12.680000 11.290000 ;
      RECT 12.400000 11.570000 12.680000 11.710000 ;
      RECT 12.400000 12.080000 12.680000 12.500000 ;
      RECT 12.400000 12.640000 12.680000 13.060000 ;
      RECT 12.400000 13.200000 12.680000 13.620000 ;
      RECT 12.400000 13.760000 12.680000 14.180000 ;
      RECT 12.400000 14.320000 12.680000 14.740000 ;
      RECT 12.405000  0.000000 12.675000  0.470000 ;
      RECT 12.405000  7.370000 12.675000  7.980000 ;
      RECT 12.405000 14.880000 12.675000 15.350000 ;
      RECT 12.815000  0.000000 16.830000  0.330000 ;
      RECT 12.815000  7.510000 16.830000  7.840000 ;
      RECT 12.815000 15.020000 16.830000 15.350000 ;
      RECT 12.820000  0.750000 16.830000  0.890000 ;
      RECT 12.820000  1.310000 16.830000  1.450000 ;
      RECT 12.820000  1.870000 16.830000  2.010000 ;
      RECT 12.820000  2.430000 16.830000  2.570000 ;
      RECT 12.820000  2.990000 16.830000  3.130000 ;
      RECT 12.820000  4.710000 16.830000  4.850000 ;
      RECT 12.820000  5.270000 16.830000  5.410000 ;
      RECT 12.820000  5.830000 16.830000  5.970000 ;
      RECT 12.820000  6.390000 16.830000  6.530000 ;
      RECT 12.820000  6.950000 16.830000  7.090000 ;
      RECT 12.820000  8.260000 16.830000  8.400000 ;
      RECT 12.820000  8.820000 16.830000  8.960000 ;
      RECT 12.820000  9.380000 16.830000  9.520000 ;
      RECT 12.820000  9.940000 16.830000 10.080000 ;
      RECT 12.820000 10.500000 16.830000 10.640000 ;
      RECT 12.820000 12.220000 16.830000 12.360000 ;
      RECT 12.820000 12.780000 16.830000 12.920000 ;
      RECT 12.820000 13.340000 16.830000 13.480000 ;
      RECT 12.820000 13.900000 16.830000 14.040000 ;
      RECT 12.820000 14.460000 16.830000 14.600000 ;
      RECT 16.500000  0.330000 16.830000  0.750000 ;
      RECT 16.500000  0.890000 16.830000  1.310000 ;
      RECT 16.500000  1.450000 16.830000  1.870000 ;
      RECT 16.500000  2.010000 16.830000  2.430000 ;
      RECT 16.500000  2.570000 16.830000  2.990000 ;
      RECT 16.500000  3.130000 16.830000  3.645000 ;
      RECT 16.500000  4.195000 16.830000  4.710000 ;
      RECT 16.500000  4.850000 16.830000  5.270000 ;
      RECT 16.500000  5.410000 16.830000  5.830000 ;
      RECT 16.500000  5.970000 16.830000  6.390000 ;
      RECT 16.500000  6.530000 16.830000  6.950000 ;
      RECT 16.500000  7.090000 16.830000  7.510000 ;
      RECT 16.500000  7.840000 16.830000  8.260000 ;
      RECT 16.500000  8.400000 16.830000  8.820000 ;
      RECT 16.500000  8.960000 16.830000  9.380000 ;
      RECT 16.500000  9.520000 16.830000  9.940000 ;
      RECT 16.500000 10.080000 16.830000 10.500000 ;
      RECT 16.500000 10.640000 16.830000 11.155000 ;
      RECT 16.500000 11.705000 16.830000 12.220000 ;
      RECT 16.500000 12.360000 16.830000 12.780000 ;
      RECT 16.500000 12.920000 16.830000 13.340000 ;
      RECT 16.500000 13.480000 16.830000 13.900000 ;
      RECT 16.500000 14.040000 16.830000 14.460000 ;
      RECT 16.500000 14.600000 16.830000 15.020000 ;
    LAYER met4 ;
      RECT  0.315000  0.315000  2.325000  2.325000 ;
      RECT  0.315000  2.920000  2.325000  4.930000 ;
      RECT  0.315000  5.515000  2.325000  7.525000 ;
      RECT  0.315000  7.825000  2.325000  9.835000 ;
      RECT  0.315000 10.430000  2.325000 12.440000 ;
      RECT  0.315000 13.025000  2.325000 15.035000 ;
      RECT  3.290000  0.315000  5.300000  2.325000 ;
      RECT  3.290000  2.920000  5.300000  4.930000 ;
      RECT  3.290000  5.515000  5.300000  7.525000 ;
      RECT  3.290000  7.825000  5.300000  9.835000 ;
      RECT  3.290000 10.430000  5.300000 12.440000 ;
      RECT  3.290000 13.025000  5.300000 15.035000 ;
      RECT  6.255000  0.315000  8.265000  2.325000 ;
      RECT  6.255000  2.920000  8.265000  4.930000 ;
      RECT  6.255000  5.515000  8.265000  7.525000 ;
      RECT  6.255000  7.825000  8.265000  9.835000 ;
      RECT  6.255000 10.430000  8.265000 12.440000 ;
      RECT  6.255000 13.025000  8.265000 15.035000 ;
      RECT  8.565000  0.315000 10.575000  2.325000 ;
      RECT  8.565000  2.920000 10.575000  4.930000 ;
      RECT  8.565000  5.515000 10.575000  7.525000 ;
      RECT  8.565000  7.825000 10.575000  9.835000 ;
      RECT  8.565000 10.430000 10.575000 12.440000 ;
      RECT  8.565000 13.025000 10.575000 15.035000 ;
      RECT 11.540000  0.315000 13.550000  2.325000 ;
      RECT 11.540000  2.920000 13.550000  4.930000 ;
      RECT 11.540000  5.515000 13.550000  7.525000 ;
      RECT 11.540000  7.825000 13.550000  9.835000 ;
      RECT 11.540000 10.430000 13.550000 12.440000 ;
      RECT 11.540000 13.025000 13.550000 15.035000 ;
      RECT 14.505000  0.315000 16.515000  2.325000 ;
      RECT 14.505000  2.920000 16.515000  4.930000 ;
      RECT 14.505000  5.515000 16.515000  7.525000 ;
      RECT 14.505000  7.825000 16.515000  9.835000 ;
      RECT 14.505000 10.430000 16.515000 12.440000 ;
      RECT 14.505000 13.025000 16.515000 15.035000 ;
    LAYER pwell ;
      RECT  4.470000  4.105000  4.590000  4.360000 ;
      RECT  4.470000 11.615000  4.590000 11.870000 ;
      RECT 12.720000  4.105000 12.840000  4.360000 ;
      RECT 12.720000 11.615000 12.840000 11.870000 ;
    LAYER via ;
      RECT  0.035000  0.265000  0.295000  0.525000 ;
      RECT  0.035000  0.585000  0.295000  0.845000 ;
      RECT  0.035000  0.905000  0.295000  1.165000 ;
      RECT  0.035000  1.225000  0.295000  1.485000 ;
      RECT  0.035000  1.545000  0.295000  1.805000 ;
      RECT  0.035000  1.865000  0.295000  2.125000 ;
      RECT  0.035000  2.185000  0.295000  2.445000 ;
      RECT  0.035000  2.505000  0.295000  2.765000 ;
      RECT  0.035000  2.825000  0.295000  3.085000 ;
      RECT  0.035000  3.145000  0.295000  3.405000 ;
      RECT  0.035000  4.435000  0.295000  4.695000 ;
      RECT  0.035000  4.755000  0.295000  5.015000 ;
      RECT  0.035000  5.075000  0.295000  5.335000 ;
      RECT  0.035000  5.395000  0.295000  5.655000 ;
      RECT  0.035000  5.715000  0.295000  5.975000 ;
      RECT  0.035000  6.035000  0.295000  6.295000 ;
      RECT  0.035000  6.355000  0.295000  6.615000 ;
      RECT  0.035000  6.675000  0.295000  6.935000 ;
      RECT  0.035000  6.995000  0.295000  7.255000 ;
      RECT  0.035000  7.315000  0.295000  7.575000 ;
      RECT  0.035000  7.775000  0.295000  8.035000 ;
      RECT  0.035000  8.095000  0.295000  8.355000 ;
      RECT  0.035000  8.415000  0.295000  8.675000 ;
      RECT  0.035000  8.735000  0.295000  8.995000 ;
      RECT  0.035000  9.055000  0.295000  9.315000 ;
      RECT  0.035000  9.375000  0.295000  9.635000 ;
      RECT  0.035000  9.695000  0.295000  9.955000 ;
      RECT  0.035000 10.015000  0.295000 10.275000 ;
      RECT  0.035000 10.335000  0.295000 10.595000 ;
      RECT  0.035000 10.655000  0.295000 10.915000 ;
      RECT  0.035000 11.945000  0.295000 12.205000 ;
      RECT  0.035000 12.265000  0.295000 12.525000 ;
      RECT  0.035000 12.585000  0.295000 12.845000 ;
      RECT  0.035000 12.905000  0.295000 13.165000 ;
      RECT  0.035000 13.225000  0.295000 13.485000 ;
      RECT  0.035000 13.545000  0.295000 13.805000 ;
      RECT  0.035000 13.865000  0.295000 14.125000 ;
      RECT  0.035000 14.185000  0.295000 14.445000 ;
      RECT  0.035000 14.505000  0.295000 14.765000 ;
      RECT  0.035000 14.825000  0.295000 15.085000 ;
      RECT  0.440000  0.035000  0.700000  0.295000 ;
      RECT  0.440000  7.545000  0.700000  7.805000 ;
      RECT  0.440000 15.055000  0.700000 15.315000 ;
      RECT  0.525000  3.790000  0.785000  4.050000 ;
      RECT  0.525000 11.300000  0.785000 11.560000 ;
      RECT  0.760000  0.035000  1.020000  0.295000 ;
      RECT  0.760000  7.545000  1.020000  7.805000 ;
      RECT  0.760000 15.055000  1.020000 15.315000 ;
      RECT  0.845000  3.790000  1.105000  4.050000 ;
      RECT  0.845000 11.300000  1.105000 11.560000 ;
      RECT  1.080000  0.035000  1.340000  0.295000 ;
      RECT  1.080000  7.545000  1.340000  7.805000 ;
      RECT  1.080000 15.055000  1.340000 15.315000 ;
      RECT  1.165000  3.790000  1.425000  4.050000 ;
      RECT  1.165000 11.300000  1.425000 11.560000 ;
      RECT  1.400000  0.035000  1.660000  0.295000 ;
      RECT  1.400000  7.545000  1.660000  7.805000 ;
      RECT  1.400000 15.055000  1.660000 15.315000 ;
      RECT  1.485000  3.790000  1.745000  4.050000 ;
      RECT  1.485000 11.300000  1.745000 11.560000 ;
      RECT  1.720000  0.035000  1.980000  0.295000 ;
      RECT  1.720000  7.545000  1.980000  7.805000 ;
      RECT  1.720000 15.055000  1.980000 15.315000 ;
      RECT  1.805000  3.790000  2.065000  4.050000 ;
      RECT  1.805000 11.300000  2.065000 11.560000 ;
      RECT  2.040000  0.035000  2.300000  0.295000 ;
      RECT  2.040000  7.545000  2.300000  7.805000 ;
      RECT  2.040000 15.055000  2.300000 15.315000 ;
      RECT  2.125000  3.790000  2.385000  4.050000 ;
      RECT  2.125000 11.300000  2.385000 11.560000 ;
      RECT  2.360000  0.035000  2.620000  0.295000 ;
      RECT  2.360000  7.545000  2.620000  7.805000 ;
      RECT  2.360000 15.055000  2.620000 15.315000 ;
      RECT  2.445000  3.790000  2.705000  4.050000 ;
      RECT  2.445000 11.300000  2.705000 11.560000 ;
      RECT  2.680000  0.035000  2.940000  0.295000 ;
      RECT  2.680000  7.545000  2.940000  7.805000 ;
      RECT  2.680000 15.055000  2.940000 15.315000 ;
      RECT  2.765000  3.790000  3.025000  4.050000 ;
      RECT  2.765000 11.300000  3.025000 11.560000 ;
      RECT  3.000000  0.035000  3.260000  0.295000 ;
      RECT  3.000000  7.545000  3.260000  7.805000 ;
      RECT  3.000000 15.055000  3.260000 15.315000 ;
      RECT  3.085000  3.790000  3.345000  4.050000 ;
      RECT  3.085000 11.300000  3.345000 11.560000 ;
      RECT  3.320000  0.035000  3.580000  0.295000 ;
      RECT  3.320000  7.545000  3.580000  7.805000 ;
      RECT  3.320000 15.055000  3.580000 15.315000 ;
      RECT  3.405000  3.790000  3.665000  4.050000 ;
      RECT  3.405000 11.300000  3.665000 11.560000 ;
      RECT  3.640000  0.035000  3.900000  0.295000 ;
      RECT  3.640000  7.545000  3.900000  7.805000 ;
      RECT  3.640000 15.055000  3.900000 15.315000 ;
      RECT  3.725000  3.790000  3.985000  4.050000 ;
      RECT  3.725000 11.300000  3.985000 11.560000 ;
      RECT  4.160000  0.500000  4.420000  0.760000 ;
      RECT  4.160000  0.820000  4.420000  1.080000 ;
      RECT  4.160000  1.140000  4.420000  1.400000 ;
      RECT  4.160000  1.460000  4.420000  1.720000 ;
      RECT  4.160000  1.780000  4.420000  2.040000 ;
      RECT  4.160000  2.100000  4.420000  2.360000 ;
      RECT  4.160000  2.420000  4.420000  2.680000 ;
      RECT  4.160000  2.740000  4.420000  3.000000 ;
      RECT  4.160000  3.060000  4.420000  3.320000 ;
      RECT  4.160000  3.380000  4.420000  3.640000 ;
      RECT  4.160000  4.200000  4.420000  4.460000 ;
      RECT  4.160000  4.520000  4.420000  4.780000 ;
      RECT  4.160000  4.840000  4.420000  5.100000 ;
      RECT  4.160000  5.160000  4.420000  5.420000 ;
      RECT  4.160000  5.480000  4.420000  5.740000 ;
      RECT  4.160000  5.800000  4.420000  6.060000 ;
      RECT  4.160000  6.120000  4.420000  6.380000 ;
      RECT  4.160000  6.440000  4.420000  6.700000 ;
      RECT  4.160000  6.760000  4.420000  7.020000 ;
      RECT  4.160000  7.080000  4.420000  7.340000 ;
      RECT  4.160000  8.010000  4.420000  8.270000 ;
      RECT  4.160000  8.330000  4.420000  8.590000 ;
      RECT  4.160000  8.650000  4.420000  8.910000 ;
      RECT  4.160000  8.970000  4.420000  9.230000 ;
      RECT  4.160000  9.290000  4.420000  9.550000 ;
      RECT  4.160000  9.610000  4.420000  9.870000 ;
      RECT  4.160000  9.930000  4.420000 10.190000 ;
      RECT  4.160000 10.250000  4.420000 10.510000 ;
      RECT  4.160000 10.570000  4.420000 10.830000 ;
      RECT  4.160000 10.890000  4.420000 11.150000 ;
      RECT  4.160000 11.710000  4.420000 11.970000 ;
      RECT  4.160000 12.030000  4.420000 12.290000 ;
      RECT  4.160000 12.350000  4.420000 12.610000 ;
      RECT  4.160000 12.670000  4.420000 12.930000 ;
      RECT  4.160000 12.990000  4.420000 13.250000 ;
      RECT  4.160000 13.310000  4.420000 13.570000 ;
      RECT  4.160000 13.630000  4.420000 13.890000 ;
      RECT  4.160000 13.950000  4.420000 14.210000 ;
      RECT  4.160000 14.270000  4.420000 14.530000 ;
      RECT  4.160000 14.590000  4.420000 14.850000 ;
      RECT  4.595000  3.790000  4.855000  4.050000 ;
      RECT  4.595000 11.300000  4.855000 11.560000 ;
      RECT  4.710000  0.035000  4.970000  0.295000 ;
      RECT  4.710000  7.545000  4.970000  7.805000 ;
      RECT  4.710000 15.055000  4.970000 15.315000 ;
      RECT  4.915000  3.790000  5.175000  4.050000 ;
      RECT  4.915000 11.300000  5.175000 11.560000 ;
      RECT  5.030000  0.035000  5.290000  0.295000 ;
      RECT  5.030000  7.545000  5.290000  7.805000 ;
      RECT  5.030000 15.055000  5.290000 15.315000 ;
      RECT  5.235000  3.790000  5.495000  4.050000 ;
      RECT  5.235000 11.300000  5.495000 11.560000 ;
      RECT  5.350000  0.035000  5.610000  0.295000 ;
      RECT  5.350000  7.545000  5.610000  7.805000 ;
      RECT  5.350000 15.055000  5.610000 15.315000 ;
      RECT  5.555000  3.790000  5.815000  4.050000 ;
      RECT  5.555000 11.300000  5.815000 11.560000 ;
      RECT  5.670000  0.035000  5.930000  0.295000 ;
      RECT  5.670000  7.545000  5.930000  7.805000 ;
      RECT  5.670000 15.055000  5.930000 15.315000 ;
      RECT  5.875000  3.790000  6.135000  4.050000 ;
      RECT  5.875000 11.300000  6.135000 11.560000 ;
      RECT  5.990000  0.035000  6.250000  0.295000 ;
      RECT  5.990000  7.545000  6.250000  7.805000 ;
      RECT  5.990000 15.055000  6.250000 15.315000 ;
      RECT  6.195000  3.790000  6.455000  4.050000 ;
      RECT  6.195000 11.300000  6.455000 11.560000 ;
      RECT  6.310000  0.035000  6.570000  0.295000 ;
      RECT  6.310000  7.545000  6.570000  7.805000 ;
      RECT  6.310000 15.055000  6.570000 15.315000 ;
      RECT  6.515000  3.790000  6.775000  4.050000 ;
      RECT  6.515000 11.300000  6.775000 11.560000 ;
      RECT  6.630000  0.035000  6.890000  0.295000 ;
      RECT  6.630000  7.545000  6.890000  7.805000 ;
      RECT  6.630000 15.055000  6.890000 15.315000 ;
      RECT  6.835000  3.790000  7.095000  4.050000 ;
      RECT  6.835000 11.300000  7.095000 11.560000 ;
      RECT  6.950000  0.035000  7.210000  0.295000 ;
      RECT  6.950000  7.545000  7.210000  7.805000 ;
      RECT  6.950000 15.055000  7.210000 15.315000 ;
      RECT  7.155000  3.790000  7.415000  4.050000 ;
      RECT  7.155000 11.300000  7.415000 11.560000 ;
      RECT  7.270000  0.035000  7.530000  0.295000 ;
      RECT  7.270000  7.545000  7.530000  7.805000 ;
      RECT  7.270000 15.055000  7.530000 15.315000 ;
      RECT  7.475000  3.790000  7.735000  4.050000 ;
      RECT  7.475000 11.300000  7.735000 11.560000 ;
      RECT  7.590000  0.035000  7.850000  0.295000 ;
      RECT  7.590000  7.545000  7.850000  7.805000 ;
      RECT  7.590000 15.055000  7.850000 15.315000 ;
      RECT  7.795000  3.790000  8.055000  4.050000 ;
      RECT  7.795000 11.300000  8.055000 11.560000 ;
      RECT  7.910000  0.035000  8.170000  0.295000 ;
      RECT  7.910000  7.545000  8.170000  7.805000 ;
      RECT  7.910000 15.055000  8.170000 15.315000 ;
      RECT  8.285000  0.265000  8.545000  0.525000 ;
      RECT  8.285000  0.585000  8.545000  0.845000 ;
      RECT  8.285000  0.905000  8.545000  1.165000 ;
      RECT  8.285000  1.225000  8.545000  1.485000 ;
      RECT  8.285000  1.545000  8.545000  1.805000 ;
      RECT  8.285000  1.865000  8.545000  2.125000 ;
      RECT  8.285000  2.185000  8.545000  2.445000 ;
      RECT  8.285000  2.505000  8.545000  2.765000 ;
      RECT  8.285000  2.825000  8.545000  3.085000 ;
      RECT  8.285000  3.145000  8.545000  3.405000 ;
      RECT  8.285000  4.435000  8.545000  4.695000 ;
      RECT  8.285000  4.755000  8.545000  5.015000 ;
      RECT  8.285000  5.075000  8.545000  5.335000 ;
      RECT  8.285000  5.395000  8.545000  5.655000 ;
      RECT  8.285000  5.715000  8.545000  5.975000 ;
      RECT  8.285000  6.035000  8.545000  6.295000 ;
      RECT  8.285000  6.355000  8.545000  6.615000 ;
      RECT  8.285000  6.675000  8.545000  6.935000 ;
      RECT  8.285000  6.995000  8.545000  7.255000 ;
      RECT  8.285000  7.315000  8.545000  7.575000 ;
      RECT  8.285000  7.775000  8.545000  8.035000 ;
      RECT  8.285000  8.095000  8.545000  8.355000 ;
      RECT  8.285000  8.415000  8.545000  8.675000 ;
      RECT  8.285000  8.735000  8.545000  8.995000 ;
      RECT  8.285000  9.055000  8.545000  9.315000 ;
      RECT  8.285000  9.375000  8.545000  9.635000 ;
      RECT  8.285000  9.695000  8.545000  9.955000 ;
      RECT  8.285000 10.015000  8.545000 10.275000 ;
      RECT  8.285000 10.335000  8.545000 10.595000 ;
      RECT  8.285000 10.655000  8.545000 10.915000 ;
      RECT  8.285000 11.945000  8.545000 12.205000 ;
      RECT  8.285000 12.265000  8.545000 12.525000 ;
      RECT  8.285000 12.585000  8.545000 12.845000 ;
      RECT  8.285000 12.905000  8.545000 13.165000 ;
      RECT  8.285000 13.225000  8.545000 13.485000 ;
      RECT  8.285000 13.545000  8.545000 13.805000 ;
      RECT  8.285000 13.865000  8.545000 14.125000 ;
      RECT  8.285000 14.185000  8.545000 14.445000 ;
      RECT  8.285000 14.505000  8.545000 14.765000 ;
      RECT  8.285000 14.825000  8.545000 15.085000 ;
      RECT  8.690000  0.035000  8.950000  0.295000 ;
      RECT  8.690000  7.545000  8.950000  7.805000 ;
      RECT  8.690000 15.055000  8.950000 15.315000 ;
      RECT  8.775000  3.790000  9.035000  4.050000 ;
      RECT  8.775000 11.300000  9.035000 11.560000 ;
      RECT  9.010000  0.035000  9.270000  0.295000 ;
      RECT  9.010000  7.545000  9.270000  7.805000 ;
      RECT  9.010000 15.055000  9.270000 15.315000 ;
      RECT  9.095000  3.790000  9.355000  4.050000 ;
      RECT  9.095000 11.300000  9.355000 11.560000 ;
      RECT  9.330000  0.035000  9.590000  0.295000 ;
      RECT  9.330000  7.545000  9.590000  7.805000 ;
      RECT  9.330000 15.055000  9.590000 15.315000 ;
      RECT  9.415000  3.790000  9.675000  4.050000 ;
      RECT  9.415000 11.300000  9.675000 11.560000 ;
      RECT  9.650000  0.035000  9.910000  0.295000 ;
      RECT  9.650000  7.545000  9.910000  7.805000 ;
      RECT  9.650000 15.055000  9.910000 15.315000 ;
      RECT  9.735000  3.790000  9.995000  4.050000 ;
      RECT  9.735000 11.300000  9.995000 11.560000 ;
      RECT  9.970000  0.035000 10.230000  0.295000 ;
      RECT  9.970000  7.545000 10.230000  7.805000 ;
      RECT  9.970000 15.055000 10.230000 15.315000 ;
      RECT 10.055000  3.790000 10.315000  4.050000 ;
      RECT 10.055000 11.300000 10.315000 11.560000 ;
      RECT 10.290000  0.035000 10.550000  0.295000 ;
      RECT 10.290000  7.545000 10.550000  7.805000 ;
      RECT 10.290000 15.055000 10.550000 15.315000 ;
      RECT 10.375000  3.790000 10.635000  4.050000 ;
      RECT 10.375000 11.300000 10.635000 11.560000 ;
      RECT 10.610000  0.035000 10.870000  0.295000 ;
      RECT 10.610000  7.545000 10.870000  7.805000 ;
      RECT 10.610000 15.055000 10.870000 15.315000 ;
      RECT 10.695000  3.790000 10.955000  4.050000 ;
      RECT 10.695000 11.300000 10.955000 11.560000 ;
      RECT 10.930000  0.035000 11.190000  0.295000 ;
      RECT 10.930000  7.545000 11.190000  7.805000 ;
      RECT 10.930000 15.055000 11.190000 15.315000 ;
      RECT 11.015000  3.790000 11.275000  4.050000 ;
      RECT 11.015000 11.300000 11.275000 11.560000 ;
      RECT 11.250000  0.035000 11.510000  0.295000 ;
      RECT 11.250000  7.545000 11.510000  7.805000 ;
      RECT 11.250000 15.055000 11.510000 15.315000 ;
      RECT 11.335000  3.790000 11.595000  4.050000 ;
      RECT 11.335000 11.300000 11.595000 11.560000 ;
      RECT 11.570000  0.035000 11.830000  0.295000 ;
      RECT 11.570000  7.545000 11.830000  7.805000 ;
      RECT 11.570000 15.055000 11.830000 15.315000 ;
      RECT 11.655000  3.790000 11.915000  4.050000 ;
      RECT 11.655000 11.300000 11.915000 11.560000 ;
      RECT 11.890000  0.035000 12.150000  0.295000 ;
      RECT 11.890000  7.545000 12.150000  7.805000 ;
      RECT 11.890000 15.055000 12.150000 15.315000 ;
      RECT 11.975000  3.790000 12.235000  4.050000 ;
      RECT 11.975000 11.300000 12.235000 11.560000 ;
      RECT 12.410000  0.500000 12.670000  0.760000 ;
      RECT 12.410000  0.820000 12.670000  1.080000 ;
      RECT 12.410000  1.140000 12.670000  1.400000 ;
      RECT 12.410000  1.460000 12.670000  1.720000 ;
      RECT 12.410000  1.780000 12.670000  2.040000 ;
      RECT 12.410000  2.100000 12.670000  2.360000 ;
      RECT 12.410000  2.420000 12.670000  2.680000 ;
      RECT 12.410000  2.740000 12.670000  3.000000 ;
      RECT 12.410000  3.060000 12.670000  3.320000 ;
      RECT 12.410000  3.380000 12.670000  3.640000 ;
      RECT 12.410000  4.200000 12.670000  4.460000 ;
      RECT 12.410000  4.520000 12.670000  4.780000 ;
      RECT 12.410000  4.840000 12.670000  5.100000 ;
      RECT 12.410000  5.160000 12.670000  5.420000 ;
      RECT 12.410000  5.480000 12.670000  5.740000 ;
      RECT 12.410000  5.800000 12.670000  6.060000 ;
      RECT 12.410000  6.120000 12.670000  6.380000 ;
      RECT 12.410000  6.440000 12.670000  6.700000 ;
      RECT 12.410000  6.760000 12.670000  7.020000 ;
      RECT 12.410000  7.080000 12.670000  7.340000 ;
      RECT 12.410000  8.010000 12.670000  8.270000 ;
      RECT 12.410000  8.330000 12.670000  8.590000 ;
      RECT 12.410000  8.650000 12.670000  8.910000 ;
      RECT 12.410000  8.970000 12.670000  9.230000 ;
      RECT 12.410000  9.290000 12.670000  9.550000 ;
      RECT 12.410000  9.610000 12.670000  9.870000 ;
      RECT 12.410000  9.930000 12.670000 10.190000 ;
      RECT 12.410000 10.250000 12.670000 10.510000 ;
      RECT 12.410000 10.570000 12.670000 10.830000 ;
      RECT 12.410000 10.890000 12.670000 11.150000 ;
      RECT 12.410000 11.710000 12.670000 11.970000 ;
      RECT 12.410000 12.030000 12.670000 12.290000 ;
      RECT 12.410000 12.350000 12.670000 12.610000 ;
      RECT 12.410000 12.670000 12.670000 12.930000 ;
      RECT 12.410000 12.990000 12.670000 13.250000 ;
      RECT 12.410000 13.310000 12.670000 13.570000 ;
      RECT 12.410000 13.630000 12.670000 13.890000 ;
      RECT 12.410000 13.950000 12.670000 14.210000 ;
      RECT 12.410000 14.270000 12.670000 14.530000 ;
      RECT 12.410000 14.590000 12.670000 14.850000 ;
      RECT 12.845000  3.790000 13.105000  4.050000 ;
      RECT 12.845000 11.300000 13.105000 11.560000 ;
      RECT 12.960000  0.035000 13.220000  0.295000 ;
      RECT 12.960000  7.545000 13.220000  7.805000 ;
      RECT 12.960000 15.055000 13.220000 15.315000 ;
      RECT 13.165000  3.790000 13.425000  4.050000 ;
      RECT 13.165000 11.300000 13.425000 11.560000 ;
      RECT 13.280000  0.035000 13.540000  0.295000 ;
      RECT 13.280000  7.545000 13.540000  7.805000 ;
      RECT 13.280000 15.055000 13.540000 15.315000 ;
      RECT 13.485000  3.790000 13.745000  4.050000 ;
      RECT 13.485000 11.300000 13.745000 11.560000 ;
      RECT 13.600000  0.035000 13.860000  0.295000 ;
      RECT 13.600000  7.545000 13.860000  7.805000 ;
      RECT 13.600000 15.055000 13.860000 15.315000 ;
      RECT 13.805000  3.790000 14.065000  4.050000 ;
      RECT 13.805000 11.300000 14.065000 11.560000 ;
      RECT 13.920000  0.035000 14.180000  0.295000 ;
      RECT 13.920000  7.545000 14.180000  7.805000 ;
      RECT 13.920000 15.055000 14.180000 15.315000 ;
      RECT 14.125000  3.790000 14.385000  4.050000 ;
      RECT 14.125000 11.300000 14.385000 11.560000 ;
      RECT 14.240000  0.035000 14.500000  0.295000 ;
      RECT 14.240000  7.545000 14.500000  7.805000 ;
      RECT 14.240000 15.055000 14.500000 15.315000 ;
      RECT 14.445000  3.790000 14.705000  4.050000 ;
      RECT 14.445000 11.300000 14.705000 11.560000 ;
      RECT 14.560000  0.035000 14.820000  0.295000 ;
      RECT 14.560000  7.545000 14.820000  7.805000 ;
      RECT 14.560000 15.055000 14.820000 15.315000 ;
      RECT 14.765000  3.790000 15.025000  4.050000 ;
      RECT 14.765000 11.300000 15.025000 11.560000 ;
      RECT 14.880000  0.035000 15.140000  0.295000 ;
      RECT 14.880000  7.545000 15.140000  7.805000 ;
      RECT 14.880000 15.055000 15.140000 15.315000 ;
      RECT 15.085000  3.790000 15.345000  4.050000 ;
      RECT 15.085000 11.300000 15.345000 11.560000 ;
      RECT 15.200000  0.035000 15.460000  0.295000 ;
      RECT 15.200000  7.545000 15.460000  7.805000 ;
      RECT 15.200000 15.055000 15.460000 15.315000 ;
      RECT 15.405000  3.790000 15.665000  4.050000 ;
      RECT 15.405000 11.300000 15.665000 11.560000 ;
      RECT 15.520000  0.035000 15.780000  0.295000 ;
      RECT 15.520000  7.545000 15.780000  7.805000 ;
      RECT 15.520000 15.055000 15.780000 15.315000 ;
      RECT 15.725000  3.790000 15.985000  4.050000 ;
      RECT 15.725000 11.300000 15.985000 11.560000 ;
      RECT 15.840000  0.035000 16.100000  0.295000 ;
      RECT 15.840000  7.545000 16.100000  7.805000 ;
      RECT 15.840000 15.055000 16.100000 15.315000 ;
      RECT 16.045000  3.790000 16.305000  4.050000 ;
      RECT 16.045000 11.300000 16.305000 11.560000 ;
      RECT 16.160000  0.035000 16.420000  0.295000 ;
      RECT 16.160000  7.545000 16.420000  7.805000 ;
      RECT 16.160000 15.055000 16.420000 15.315000 ;
      RECT 16.535000  0.265000 16.795000  0.525000 ;
      RECT 16.535000  0.585000 16.795000  0.845000 ;
      RECT 16.535000  0.905000 16.795000  1.165000 ;
      RECT 16.535000  1.225000 16.795000  1.485000 ;
      RECT 16.535000  1.545000 16.795000  1.805000 ;
      RECT 16.535000  1.865000 16.795000  2.125000 ;
      RECT 16.535000  2.185000 16.795000  2.445000 ;
      RECT 16.535000  2.505000 16.795000  2.765000 ;
      RECT 16.535000  2.825000 16.795000  3.085000 ;
      RECT 16.535000  3.145000 16.795000  3.405000 ;
      RECT 16.535000  4.435000 16.795000  4.695000 ;
      RECT 16.535000  4.755000 16.795000  5.015000 ;
      RECT 16.535000  5.075000 16.795000  5.335000 ;
      RECT 16.535000  5.395000 16.795000  5.655000 ;
      RECT 16.535000  5.715000 16.795000  5.975000 ;
      RECT 16.535000  6.035000 16.795000  6.295000 ;
      RECT 16.535000  6.355000 16.795000  6.615000 ;
      RECT 16.535000  6.675000 16.795000  6.935000 ;
      RECT 16.535000  6.995000 16.795000  7.255000 ;
      RECT 16.535000  7.315000 16.795000  7.575000 ;
      RECT 16.535000  7.775000 16.795000  8.035000 ;
      RECT 16.535000  8.095000 16.795000  8.355000 ;
      RECT 16.535000  8.415000 16.795000  8.675000 ;
      RECT 16.535000  8.735000 16.795000  8.995000 ;
      RECT 16.535000  9.055000 16.795000  9.315000 ;
      RECT 16.535000  9.375000 16.795000  9.635000 ;
      RECT 16.535000  9.695000 16.795000  9.955000 ;
      RECT 16.535000 10.015000 16.795000 10.275000 ;
      RECT 16.535000 10.335000 16.795000 10.595000 ;
      RECT 16.535000 10.655000 16.795000 10.915000 ;
      RECT 16.535000 11.945000 16.795000 12.205000 ;
      RECT 16.535000 12.265000 16.795000 12.525000 ;
      RECT 16.535000 12.585000 16.795000 12.845000 ;
      RECT 16.535000 12.905000 16.795000 13.165000 ;
      RECT 16.535000 13.225000 16.795000 13.485000 ;
      RECT 16.535000 13.545000 16.795000 13.805000 ;
      RECT 16.535000 13.865000 16.795000 14.125000 ;
      RECT 16.535000 14.185000 16.795000 14.445000 ;
      RECT 16.535000 14.505000 16.795000 14.765000 ;
      RECT 16.535000 14.825000 16.795000 15.085000 ;
    LAYER via2 ;
      RECT  0.025000  0.520000  0.305000  0.800000 ;
      RECT  0.025000  0.920000  0.305000  1.200000 ;
      RECT  0.025000  1.320000  0.305000  1.600000 ;
      RECT  0.025000  1.720000  0.305000  2.000000 ;
      RECT  0.025000  2.120000  0.305000  2.400000 ;
      RECT  0.025000  2.520000  0.305000  2.800000 ;
      RECT  0.025000  2.920000  0.305000  3.200000 ;
      RECT  0.025000  3.320000  0.305000  3.600000 ;
      RECT  0.025000  4.240000  0.305000  4.520000 ;
      RECT  0.025000  4.640000  0.305000  4.920000 ;
      RECT  0.025000  5.040000  0.305000  5.320000 ;
      RECT  0.025000  5.440000  0.305000  5.720000 ;
      RECT  0.025000  5.840000  0.305000  6.120000 ;
      RECT  0.025000  6.240000  0.305000  6.520000 ;
      RECT  0.025000  6.640000  0.305000  6.920000 ;
      RECT  0.025000  7.040000  0.305000  7.320000 ;
      RECT  0.025000  8.030000  0.305000  8.310000 ;
      RECT  0.025000  8.430000  0.305000  8.710000 ;
      RECT  0.025000  8.830000  0.305000  9.110000 ;
      RECT  0.025000  9.230000  0.305000  9.510000 ;
      RECT  0.025000  9.630000  0.305000  9.910000 ;
      RECT  0.025000 10.030000  0.305000 10.310000 ;
      RECT  0.025000 10.430000  0.305000 10.710000 ;
      RECT  0.025000 10.830000  0.305000 11.110000 ;
      RECT  0.025000 11.750000  0.305000 12.030000 ;
      RECT  0.025000 12.150000  0.305000 12.430000 ;
      RECT  0.025000 12.550000  0.305000 12.830000 ;
      RECT  0.025000 12.950000  0.305000 13.230000 ;
      RECT  0.025000 13.350000  0.305000 13.630000 ;
      RECT  0.025000 13.750000  0.305000 14.030000 ;
      RECT  0.025000 14.150000  0.305000 14.430000 ;
      RECT  0.025000 14.550000  0.305000 14.830000 ;
      RECT  0.490000  0.025000  0.770000  0.305000 ;
      RECT  0.490000  7.535000  0.770000  7.815000 ;
      RECT  0.490000 15.045000  0.770000 15.325000 ;
      RECT  0.890000  0.025000  1.170000  0.305000 ;
      RECT  0.890000  7.535000  1.170000  7.815000 ;
      RECT  0.890000 15.045000  1.170000 15.325000 ;
      RECT  0.950000  3.780000  1.230000  4.060000 ;
      RECT  0.950000 11.290000  1.230000 11.570000 ;
      RECT  1.290000  0.025000  1.570000  0.305000 ;
      RECT  1.290000  7.535000  1.570000  7.815000 ;
      RECT  1.290000 15.045000  1.570000 15.325000 ;
      RECT  1.350000  3.780000  1.630000  4.060000 ;
      RECT  1.350000 11.290000  1.630000 11.570000 ;
      RECT  1.690000  0.025000  1.970000  0.305000 ;
      RECT  1.690000  7.535000  1.970000  7.815000 ;
      RECT  1.690000 15.045000  1.970000 15.325000 ;
      RECT  1.750000  3.780000  2.030000  4.060000 ;
      RECT  1.750000 11.290000  2.030000 11.570000 ;
      RECT  2.090000  0.025000  2.370000  0.305000 ;
      RECT  2.090000  7.535000  2.370000  7.815000 ;
      RECT  2.090000 15.045000  2.370000 15.325000 ;
      RECT  2.150000  3.780000  2.430000  4.060000 ;
      RECT  2.150000 11.290000  2.430000 11.570000 ;
      RECT  2.490000  0.025000  2.770000  0.305000 ;
      RECT  2.490000  7.535000  2.770000  7.815000 ;
      RECT  2.490000 15.045000  2.770000 15.325000 ;
      RECT  2.550000  3.780000  2.830000  4.060000 ;
      RECT  2.550000 11.290000  2.830000 11.570000 ;
      RECT  2.890000  0.025000  3.170000  0.305000 ;
      RECT  2.890000  7.535000  3.170000  7.815000 ;
      RECT  2.890000 15.045000  3.170000 15.325000 ;
      RECT  2.950000  3.780000  3.230000  4.060000 ;
      RECT  2.950000 11.290000  3.230000 11.570000 ;
      RECT  3.290000  0.025000  3.570000  0.305000 ;
      RECT  3.290000  7.535000  3.570000  7.815000 ;
      RECT  3.290000 15.045000  3.570000 15.325000 ;
      RECT  3.350000  3.780000  3.630000  4.060000 ;
      RECT  3.350000 11.290000  3.630000 11.570000 ;
      RECT  3.690000  0.025000  3.970000  0.305000 ;
      RECT  3.690000  7.535000  3.970000  7.815000 ;
      RECT  3.690000 15.045000  3.970000 15.325000 ;
      RECT  3.750000  3.780000  4.030000  4.060000 ;
      RECT  3.750000 11.290000  4.030000 11.570000 ;
      RECT  4.150000  3.780000  4.430000  4.060000 ;
      RECT  4.150000 11.290000  4.430000 11.570000 ;
      RECT  4.550000  3.780000  4.830000  4.060000 ;
      RECT  4.550000 11.290000  4.830000 11.570000 ;
      RECT  4.610000  0.025000  4.890000  0.305000 ;
      RECT  4.610000  7.535000  4.890000  7.815000 ;
      RECT  4.610000 15.045000  4.890000 15.325000 ;
      RECT  4.950000  3.780000  5.230000  4.060000 ;
      RECT  4.950000 11.290000  5.230000 11.570000 ;
      RECT  5.010000  0.025000  5.290000  0.305000 ;
      RECT  5.010000  7.535000  5.290000  7.815000 ;
      RECT  5.010000 15.045000  5.290000 15.325000 ;
      RECT  5.350000  3.780000  5.630000  4.060000 ;
      RECT  5.350000 11.290000  5.630000 11.570000 ;
      RECT  5.410000  0.025000  5.690000  0.305000 ;
      RECT  5.410000  7.535000  5.690000  7.815000 ;
      RECT  5.410000 15.045000  5.690000 15.325000 ;
      RECT  5.750000  3.780000  6.030000  4.060000 ;
      RECT  5.750000 11.290000  6.030000 11.570000 ;
      RECT  5.810000  0.025000  6.090000  0.305000 ;
      RECT  5.810000  7.535000  6.090000  7.815000 ;
      RECT  5.810000 15.045000  6.090000 15.325000 ;
      RECT  6.150000  3.780000  6.430000  4.060000 ;
      RECT  6.150000 11.290000  6.430000 11.570000 ;
      RECT  6.210000  0.025000  6.490000  0.305000 ;
      RECT  6.210000  7.535000  6.490000  7.815000 ;
      RECT  6.210000 15.045000  6.490000 15.325000 ;
      RECT  6.550000  3.780000  6.830000  4.060000 ;
      RECT  6.550000 11.290000  6.830000 11.570000 ;
      RECT  6.610000  0.025000  6.890000  0.305000 ;
      RECT  6.610000  7.535000  6.890000  7.815000 ;
      RECT  6.610000 15.045000  6.890000 15.325000 ;
      RECT  6.950000  3.780000  7.230000  4.060000 ;
      RECT  6.950000 11.290000  7.230000 11.570000 ;
      RECT  7.010000  0.025000  7.290000  0.305000 ;
      RECT  7.010000  7.535000  7.290000  7.815000 ;
      RECT  7.010000 15.045000  7.290000 15.325000 ;
      RECT  7.350000  3.780000  7.630000  4.060000 ;
      RECT  7.350000 11.290000  7.630000 11.570000 ;
      RECT  7.410000  0.025000  7.690000  0.305000 ;
      RECT  7.410000  7.535000  7.690000  7.815000 ;
      RECT  7.410000 15.045000  7.690000 15.325000 ;
      RECT  7.810000  0.025000  8.090000  0.305000 ;
      RECT  7.810000  7.535000  8.090000  7.815000 ;
      RECT  7.810000 15.045000  8.090000 15.325000 ;
      RECT  8.275000  0.520000  8.555000  0.800000 ;
      RECT  8.275000  0.920000  8.555000  1.200000 ;
      RECT  8.275000  1.320000  8.555000  1.600000 ;
      RECT  8.275000  1.720000  8.555000  2.000000 ;
      RECT  8.275000  2.120000  8.555000  2.400000 ;
      RECT  8.275000  2.520000  8.555000  2.800000 ;
      RECT  8.275000  2.920000  8.555000  3.200000 ;
      RECT  8.275000  3.320000  8.555000  3.600000 ;
      RECT  8.275000  4.240000  8.555000  4.520000 ;
      RECT  8.275000  4.640000  8.555000  4.920000 ;
      RECT  8.275000  5.040000  8.555000  5.320000 ;
      RECT  8.275000  5.440000  8.555000  5.720000 ;
      RECT  8.275000  5.840000  8.555000  6.120000 ;
      RECT  8.275000  6.240000  8.555000  6.520000 ;
      RECT  8.275000  6.640000  8.555000  6.920000 ;
      RECT  8.275000  7.040000  8.555000  7.320000 ;
      RECT  8.275000  8.030000  8.555000  8.310000 ;
      RECT  8.275000  8.430000  8.555000  8.710000 ;
      RECT  8.275000  8.830000  8.555000  9.110000 ;
      RECT  8.275000  9.230000  8.555000  9.510000 ;
      RECT  8.275000  9.630000  8.555000  9.910000 ;
      RECT  8.275000 10.030000  8.555000 10.310000 ;
      RECT  8.275000 10.430000  8.555000 10.710000 ;
      RECT  8.275000 10.830000  8.555000 11.110000 ;
      RECT  8.275000 11.750000  8.555000 12.030000 ;
      RECT  8.275000 12.150000  8.555000 12.430000 ;
      RECT  8.275000 12.550000  8.555000 12.830000 ;
      RECT  8.275000 12.950000  8.555000 13.230000 ;
      RECT  8.275000 13.350000  8.555000 13.630000 ;
      RECT  8.275000 13.750000  8.555000 14.030000 ;
      RECT  8.275000 14.150000  8.555000 14.430000 ;
      RECT  8.275000 14.550000  8.555000 14.830000 ;
      RECT  8.740000  0.025000  9.020000  0.305000 ;
      RECT  8.740000  7.535000  9.020000  7.815000 ;
      RECT  8.740000 15.045000  9.020000 15.325000 ;
      RECT  9.140000  0.025000  9.420000  0.305000 ;
      RECT  9.140000  7.535000  9.420000  7.815000 ;
      RECT  9.140000 15.045000  9.420000 15.325000 ;
      RECT  9.200000  3.780000  9.480000  4.060000 ;
      RECT  9.200000 11.290000  9.480000 11.570000 ;
      RECT  9.540000  0.025000  9.820000  0.305000 ;
      RECT  9.540000  7.535000  9.820000  7.815000 ;
      RECT  9.540000 15.045000  9.820000 15.325000 ;
      RECT  9.600000  3.780000  9.880000  4.060000 ;
      RECT  9.600000 11.290000  9.880000 11.570000 ;
      RECT  9.940000  0.025000 10.220000  0.305000 ;
      RECT  9.940000  7.535000 10.220000  7.815000 ;
      RECT  9.940000 15.045000 10.220000 15.325000 ;
      RECT 10.000000  3.780000 10.280000  4.060000 ;
      RECT 10.000000 11.290000 10.280000 11.570000 ;
      RECT 10.340000  0.025000 10.620000  0.305000 ;
      RECT 10.340000  7.535000 10.620000  7.815000 ;
      RECT 10.340000 15.045000 10.620000 15.325000 ;
      RECT 10.400000  3.780000 10.680000  4.060000 ;
      RECT 10.400000 11.290000 10.680000 11.570000 ;
      RECT 10.740000  0.025000 11.020000  0.305000 ;
      RECT 10.740000  7.535000 11.020000  7.815000 ;
      RECT 10.740000 15.045000 11.020000 15.325000 ;
      RECT 10.800000  3.780000 11.080000  4.060000 ;
      RECT 10.800000 11.290000 11.080000 11.570000 ;
      RECT 11.140000  0.025000 11.420000  0.305000 ;
      RECT 11.140000  7.535000 11.420000  7.815000 ;
      RECT 11.140000 15.045000 11.420000 15.325000 ;
      RECT 11.200000  3.780000 11.480000  4.060000 ;
      RECT 11.200000 11.290000 11.480000 11.570000 ;
      RECT 11.540000  0.025000 11.820000  0.305000 ;
      RECT 11.540000  7.535000 11.820000  7.815000 ;
      RECT 11.540000 15.045000 11.820000 15.325000 ;
      RECT 11.600000  3.780000 11.880000  4.060000 ;
      RECT 11.600000 11.290000 11.880000 11.570000 ;
      RECT 11.940000  0.025000 12.220000  0.305000 ;
      RECT 11.940000  7.535000 12.220000  7.815000 ;
      RECT 11.940000 15.045000 12.220000 15.325000 ;
      RECT 12.000000  3.780000 12.280000  4.060000 ;
      RECT 12.000000 11.290000 12.280000 11.570000 ;
      RECT 12.400000  3.780000 12.680000  4.060000 ;
      RECT 12.400000 11.290000 12.680000 11.570000 ;
      RECT 12.800000  3.780000 13.080000  4.060000 ;
      RECT 12.800000 11.290000 13.080000 11.570000 ;
      RECT 12.860000  0.025000 13.140000  0.305000 ;
      RECT 12.860000  7.535000 13.140000  7.815000 ;
      RECT 12.860000 15.045000 13.140000 15.325000 ;
      RECT 13.200000  3.780000 13.480000  4.060000 ;
      RECT 13.200000 11.290000 13.480000 11.570000 ;
      RECT 13.260000  0.025000 13.540000  0.305000 ;
      RECT 13.260000  7.535000 13.540000  7.815000 ;
      RECT 13.260000 15.045000 13.540000 15.325000 ;
      RECT 13.600000  3.780000 13.880000  4.060000 ;
      RECT 13.600000 11.290000 13.880000 11.570000 ;
      RECT 13.660000  0.025000 13.940000  0.305000 ;
      RECT 13.660000  7.535000 13.940000  7.815000 ;
      RECT 13.660000 15.045000 13.940000 15.325000 ;
      RECT 14.000000  3.780000 14.280000  4.060000 ;
      RECT 14.000000 11.290000 14.280000 11.570000 ;
      RECT 14.060000  0.025000 14.340000  0.305000 ;
      RECT 14.060000  7.535000 14.340000  7.815000 ;
      RECT 14.060000 15.045000 14.340000 15.325000 ;
      RECT 14.400000  3.780000 14.680000  4.060000 ;
      RECT 14.400000 11.290000 14.680000 11.570000 ;
      RECT 14.460000  0.025000 14.740000  0.305000 ;
      RECT 14.460000  7.535000 14.740000  7.815000 ;
      RECT 14.460000 15.045000 14.740000 15.325000 ;
      RECT 14.800000  3.780000 15.080000  4.060000 ;
      RECT 14.800000 11.290000 15.080000 11.570000 ;
      RECT 14.860000  0.025000 15.140000  0.305000 ;
      RECT 14.860000  7.535000 15.140000  7.815000 ;
      RECT 14.860000 15.045000 15.140000 15.325000 ;
      RECT 15.200000  3.780000 15.480000  4.060000 ;
      RECT 15.200000 11.290000 15.480000 11.570000 ;
      RECT 15.260000  0.025000 15.540000  0.305000 ;
      RECT 15.260000  7.535000 15.540000  7.815000 ;
      RECT 15.260000 15.045000 15.540000 15.325000 ;
      RECT 15.600000  3.780000 15.880000  4.060000 ;
      RECT 15.600000 11.290000 15.880000 11.570000 ;
      RECT 15.660000  0.025000 15.940000  0.305000 ;
      RECT 15.660000  7.535000 15.940000  7.815000 ;
      RECT 15.660000 15.045000 15.940000 15.325000 ;
      RECT 16.060000  0.025000 16.340000  0.305000 ;
      RECT 16.060000  7.535000 16.340000  7.815000 ;
      RECT 16.060000 15.045000 16.340000 15.325000 ;
      RECT 16.525000  0.520000 16.805000  0.800000 ;
      RECT 16.525000  0.920000 16.805000  1.200000 ;
      RECT 16.525000  1.320000 16.805000  1.600000 ;
      RECT 16.525000  1.720000 16.805000  2.000000 ;
      RECT 16.525000  2.120000 16.805000  2.400000 ;
      RECT 16.525000  2.520000 16.805000  2.800000 ;
      RECT 16.525000  2.920000 16.805000  3.200000 ;
      RECT 16.525000  3.320000 16.805000  3.600000 ;
      RECT 16.525000  4.240000 16.805000  4.520000 ;
      RECT 16.525000  4.640000 16.805000  4.920000 ;
      RECT 16.525000  5.040000 16.805000  5.320000 ;
      RECT 16.525000  5.440000 16.805000  5.720000 ;
      RECT 16.525000  5.840000 16.805000  6.120000 ;
      RECT 16.525000  6.240000 16.805000  6.520000 ;
      RECT 16.525000  6.640000 16.805000  6.920000 ;
      RECT 16.525000  7.040000 16.805000  7.320000 ;
      RECT 16.525000  8.030000 16.805000  8.310000 ;
      RECT 16.525000  8.430000 16.805000  8.710000 ;
      RECT 16.525000  8.830000 16.805000  9.110000 ;
      RECT 16.525000  9.230000 16.805000  9.510000 ;
      RECT 16.525000  9.630000 16.805000  9.910000 ;
      RECT 16.525000 10.030000 16.805000 10.310000 ;
      RECT 16.525000 10.430000 16.805000 10.710000 ;
      RECT 16.525000 10.830000 16.805000 11.110000 ;
      RECT 16.525000 11.750000 16.805000 12.030000 ;
      RECT 16.525000 12.150000 16.805000 12.430000 ;
      RECT 16.525000 12.550000 16.805000 12.830000 ;
      RECT 16.525000 12.950000 16.805000 13.230000 ;
      RECT 16.525000 13.350000 16.805000 13.630000 ;
      RECT 16.525000 13.750000 16.805000 14.030000 ;
      RECT 16.525000 14.150000 16.805000 14.430000 ;
      RECT 16.525000 14.550000 16.805000 14.830000 ;
  END
END sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4_top
END LIBRARY
