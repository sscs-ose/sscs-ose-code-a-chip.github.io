# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_20v0_withptap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_20v0_withptap ;
  ORIGIN  5.700000  5.910000 ;
  SIZE  12.15000 BY  41.82000 ;
  OBS
    LAYER li1 ;
      RECT -5.700000 -5.910000  6.450000 -5.500000 ;
      RECT -5.700000 -5.500000 -5.290000 35.500000 ;
      RECT -5.700000 35.500000  6.450000 35.910000 ;
      RECT -4.810000  0.045000 -4.480000 29.955000 ;
      RECT -1.480000 -4.285000  2.300000 -3.215000 ;
      RECT  0.040000  0.215000  0.710000 29.785000 ;
      RECT  5.230000  0.045000  5.560000 29.955000 ;
      RECT  6.040000 -5.500000  6.450000 35.500000 ;
    LAYER mcon ;
      RECT -5.580000 -5.425000 -5.410000 -5.255000 ;
      RECT -5.580000 -5.065000 -5.410000 -4.895000 ;
      RECT -5.580000 -4.705000 -5.410000 -4.535000 ;
      RECT -5.580000 -4.345000 -5.410000 -4.175000 ;
      RECT -5.580000 -3.985000 -5.410000 -3.815000 ;
      RECT -5.580000 -3.625000 -5.410000 -3.455000 ;
      RECT -5.580000 -3.265000 -5.410000 -3.095000 ;
      RECT -5.580000 -2.905000 -5.410000 -2.735000 ;
      RECT -5.580000 -2.545000 -5.410000 -2.375000 ;
      RECT -5.580000 -2.185000 -5.410000 -2.015000 ;
      RECT -5.580000 -1.825000 -5.410000 -1.655000 ;
      RECT -5.580000 -1.465000 -5.410000 -1.295000 ;
      RECT -5.580000 -1.105000 -5.410000 -0.935000 ;
      RECT -5.580000 -0.745000 -5.410000 -0.575000 ;
      RECT -5.580000 -0.385000 -5.410000 -0.215000 ;
      RECT -5.580000 -0.025000 -5.410000  0.145000 ;
      RECT -5.580000  0.335000 -5.410000  0.505000 ;
      RECT -5.580000  0.695000 -5.410000  0.865000 ;
      RECT -5.580000  1.055000 -5.410000  1.225000 ;
      RECT -5.580000  1.415000 -5.410000  1.585000 ;
      RECT -5.580000  1.775000 -5.410000  1.945000 ;
      RECT -5.580000  2.135000 -5.410000  2.305000 ;
      RECT -5.580000  2.495000 -5.410000  2.665000 ;
      RECT -5.580000  2.855000 -5.410000  3.025000 ;
      RECT -5.580000  3.215000 -5.410000  3.385000 ;
      RECT -5.580000  3.575000 -5.410000  3.745000 ;
      RECT -5.580000  3.935000 -5.410000  4.105000 ;
      RECT -5.580000  4.295000 -5.410000  4.465000 ;
      RECT -5.580000  4.655000 -5.410000  4.825000 ;
      RECT -5.580000  5.015000 -5.410000  5.185000 ;
      RECT -5.580000  5.375000 -5.410000  5.545000 ;
      RECT -5.580000  5.735000 -5.410000  5.905000 ;
      RECT -5.580000  6.095000 -5.410000  6.265000 ;
      RECT -5.580000  6.455000 -5.410000  6.625000 ;
      RECT -5.580000  6.815000 -5.410000  6.985000 ;
      RECT -5.580000  7.175000 -5.410000  7.345000 ;
      RECT -5.580000  7.535000 -5.410000  7.705000 ;
      RECT -5.580000  7.895000 -5.410000  8.065000 ;
      RECT -5.580000  8.255000 -5.410000  8.425000 ;
      RECT -5.580000  8.615000 -5.410000  8.785000 ;
      RECT -5.580000  8.975000 -5.410000  9.145000 ;
      RECT -5.580000  9.335000 -5.410000  9.505000 ;
      RECT -5.580000  9.695000 -5.410000  9.865000 ;
      RECT -5.580000 10.055000 -5.410000 10.225000 ;
      RECT -5.580000 10.415000 -5.410000 10.585000 ;
      RECT -5.580000 10.775000 -5.410000 10.945000 ;
      RECT -5.580000 11.135000 -5.410000 11.305000 ;
      RECT -5.580000 11.495000 -5.410000 11.665000 ;
      RECT -5.580000 11.855000 -5.410000 12.025000 ;
      RECT -5.580000 12.215000 -5.410000 12.385000 ;
      RECT -5.580000 12.575000 -5.410000 12.745000 ;
      RECT -5.580000 12.935000 -5.410000 13.105000 ;
      RECT -5.580000 13.295000 -5.410000 13.465000 ;
      RECT -5.580000 13.655000 -5.410000 13.825000 ;
      RECT -5.580000 14.015000 -5.410000 14.185000 ;
      RECT -5.580000 14.375000 -5.410000 14.545000 ;
      RECT -5.580000 14.735000 -5.410000 14.905000 ;
      RECT -5.580000 15.095000 -5.410000 15.265000 ;
      RECT -5.580000 15.455000 -5.410000 15.625000 ;
      RECT -5.580000 15.815000 -5.410000 15.985000 ;
      RECT -5.580000 16.175000 -5.410000 16.345000 ;
      RECT -5.580000 16.535000 -5.410000 16.705000 ;
      RECT -5.580000 16.895000 -5.410000 17.065000 ;
      RECT -5.580000 17.255000 -5.410000 17.425000 ;
      RECT -5.580000 17.615000 -5.410000 17.785000 ;
      RECT -5.580000 17.975000 -5.410000 18.145000 ;
      RECT -5.580000 18.335000 -5.410000 18.505000 ;
      RECT -5.580000 18.695000 -5.410000 18.865000 ;
      RECT -5.580000 19.055000 -5.410000 19.225000 ;
      RECT -5.580000 19.415000 -5.410000 19.585000 ;
      RECT -5.580000 19.775000 -5.410000 19.945000 ;
      RECT -5.580000 20.135000 -5.410000 20.305000 ;
      RECT -5.580000 20.495000 -5.410000 20.665000 ;
      RECT -5.580000 20.855000 -5.410000 21.025000 ;
      RECT -5.580000 21.215000 -5.410000 21.385000 ;
      RECT -5.580000 21.575000 -5.410000 21.745000 ;
      RECT -5.580000 21.935000 -5.410000 22.105000 ;
      RECT -5.580000 22.295000 -5.410000 22.465000 ;
      RECT -5.580000 22.655000 -5.410000 22.825000 ;
      RECT -5.580000 23.015000 -5.410000 23.185000 ;
      RECT -5.580000 23.375000 -5.410000 23.545000 ;
      RECT -5.580000 23.735000 -5.410000 23.905000 ;
      RECT -5.580000 24.095000 -5.410000 24.265000 ;
      RECT -5.580000 24.455000 -5.410000 24.625000 ;
      RECT -5.580000 24.815000 -5.410000 24.985000 ;
      RECT -5.580000 25.175000 -5.410000 25.345000 ;
      RECT -5.580000 25.535000 -5.410000 25.705000 ;
      RECT -5.580000 25.895000 -5.410000 26.065000 ;
      RECT -5.580000 26.255000 -5.410000 26.425000 ;
      RECT -5.580000 26.615000 -5.410000 26.785000 ;
      RECT -5.580000 26.975000 -5.410000 27.145000 ;
      RECT -5.580000 27.335000 -5.410000 27.505000 ;
      RECT -5.580000 27.695000 -5.410000 27.865000 ;
      RECT -5.580000 28.055000 -5.410000 28.225000 ;
      RECT -5.580000 28.415000 -5.410000 28.585000 ;
      RECT -5.580000 28.775000 -5.410000 28.945000 ;
      RECT -5.580000 29.135000 -5.410000 29.305000 ;
      RECT -5.580000 29.495000 -5.410000 29.665000 ;
      RECT -5.580000 29.855000 -5.410000 30.025000 ;
      RECT -5.580000 30.215000 -5.410000 30.385000 ;
      RECT -5.580000 30.575000 -5.410000 30.745000 ;
      RECT -5.580000 30.935000 -5.410000 31.105000 ;
      RECT -5.580000 31.295000 -5.410000 31.465000 ;
      RECT -5.580000 31.655000 -5.410000 31.825000 ;
      RECT -5.580000 32.015000 -5.410000 32.185000 ;
      RECT -5.580000 32.375000 -5.410000 32.545000 ;
      RECT -5.580000 32.735000 -5.410000 32.905000 ;
      RECT -5.580000 33.095000 -5.410000 33.265000 ;
      RECT -5.580000 33.455000 -5.410000 33.625000 ;
      RECT -5.580000 33.815000 -5.410000 33.985000 ;
      RECT -5.580000 34.175000 -5.410000 34.345000 ;
      RECT -5.580000 34.535000 -5.410000 34.705000 ;
      RECT -5.580000 34.895000 -5.410000 35.065000 ;
      RECT -5.580000 35.255000 -5.410000 35.425000 ;
      RECT -4.930000 -5.790000 -4.760000 -5.620000 ;
      RECT -4.930000 35.620000 -4.760000 35.790000 ;
      RECT -4.730000  0.155000 -4.560000  0.325000 ;
      RECT -4.730000  0.515000 -4.560000  0.685000 ;
      RECT -4.730000  0.875000 -4.560000  1.045000 ;
      RECT -4.730000  1.235000 -4.560000  1.405000 ;
      RECT -4.730000  1.595000 -4.560000  1.765000 ;
      RECT -4.730000  1.955000 -4.560000  2.125000 ;
      RECT -4.730000  2.315000 -4.560000  2.485000 ;
      RECT -4.730000  2.675000 -4.560000  2.845000 ;
      RECT -4.730000  3.035000 -4.560000  3.205000 ;
      RECT -4.730000  3.395000 -4.560000  3.565000 ;
      RECT -4.730000  3.755000 -4.560000  3.925000 ;
      RECT -4.730000  4.115000 -4.560000  4.285000 ;
      RECT -4.730000  4.475000 -4.560000  4.645000 ;
      RECT -4.730000  4.835000 -4.560000  5.005000 ;
      RECT -4.730000  5.195000 -4.560000  5.365000 ;
      RECT -4.730000  5.555000 -4.560000  5.725000 ;
      RECT -4.730000  5.915000 -4.560000  6.085000 ;
      RECT -4.730000  6.275000 -4.560000  6.445000 ;
      RECT -4.730000  6.635000 -4.560000  6.805000 ;
      RECT -4.730000  6.995000 -4.560000  7.165000 ;
      RECT -4.730000  7.355000 -4.560000  7.525000 ;
      RECT -4.730000  7.715000 -4.560000  7.885000 ;
      RECT -4.730000  8.075000 -4.560000  8.245000 ;
      RECT -4.730000  8.435000 -4.560000  8.605000 ;
      RECT -4.730000  8.795000 -4.560000  8.965000 ;
      RECT -4.730000  9.155000 -4.560000  9.325000 ;
      RECT -4.730000  9.515000 -4.560000  9.685000 ;
      RECT -4.730000  9.875000 -4.560000 10.045000 ;
      RECT -4.730000 10.235000 -4.560000 10.405000 ;
      RECT -4.730000 10.595000 -4.560000 10.765000 ;
      RECT -4.730000 10.955000 -4.560000 11.125000 ;
      RECT -4.730000 11.315000 -4.560000 11.485000 ;
      RECT -4.730000 11.675000 -4.560000 11.845000 ;
      RECT -4.730000 12.035000 -4.560000 12.205000 ;
      RECT -4.730000 12.395000 -4.560000 12.565000 ;
      RECT -4.730000 12.755000 -4.560000 12.925000 ;
      RECT -4.730000 13.115000 -4.560000 13.285000 ;
      RECT -4.730000 13.475000 -4.560000 13.645000 ;
      RECT -4.730000 13.835000 -4.560000 14.005000 ;
      RECT -4.730000 14.195000 -4.560000 14.365000 ;
      RECT -4.730000 14.555000 -4.560000 14.725000 ;
      RECT -4.730000 14.915000 -4.560000 15.085000 ;
      RECT -4.730000 15.275000 -4.560000 15.445000 ;
      RECT -4.730000 15.635000 -4.560000 15.805000 ;
      RECT -4.730000 15.995000 -4.560000 16.165000 ;
      RECT -4.730000 16.355000 -4.560000 16.525000 ;
      RECT -4.730000 16.715000 -4.560000 16.885000 ;
      RECT -4.730000 17.075000 -4.560000 17.245000 ;
      RECT -4.730000 17.435000 -4.560000 17.605000 ;
      RECT -4.730000 17.795000 -4.560000 17.965000 ;
      RECT -4.730000 18.155000 -4.560000 18.325000 ;
      RECT -4.730000 18.515000 -4.560000 18.685000 ;
      RECT -4.730000 18.875000 -4.560000 19.045000 ;
      RECT -4.730000 19.235000 -4.560000 19.405000 ;
      RECT -4.730000 19.595000 -4.560000 19.765000 ;
      RECT -4.730000 19.955000 -4.560000 20.125000 ;
      RECT -4.730000 20.315000 -4.560000 20.485000 ;
      RECT -4.730000 20.675000 -4.560000 20.845000 ;
      RECT -4.730000 21.035000 -4.560000 21.205000 ;
      RECT -4.730000 21.395000 -4.560000 21.565000 ;
      RECT -4.730000 21.755000 -4.560000 21.925000 ;
      RECT -4.730000 22.115000 -4.560000 22.285000 ;
      RECT -4.730000 22.475000 -4.560000 22.645000 ;
      RECT -4.730000 22.835000 -4.560000 23.005000 ;
      RECT -4.730000 23.195000 -4.560000 23.365000 ;
      RECT -4.730000 23.555000 -4.560000 23.725000 ;
      RECT -4.730000 23.915000 -4.560000 24.085000 ;
      RECT -4.730000 24.275000 -4.560000 24.445000 ;
      RECT -4.730000 24.635000 -4.560000 24.805000 ;
      RECT -4.730000 24.995000 -4.560000 25.165000 ;
      RECT -4.730000 25.355000 -4.560000 25.525000 ;
      RECT -4.730000 25.715000 -4.560000 25.885000 ;
      RECT -4.730000 26.075000 -4.560000 26.245000 ;
      RECT -4.730000 26.435000 -4.560000 26.605000 ;
      RECT -4.730000 26.795000 -4.560000 26.965000 ;
      RECT -4.730000 27.155000 -4.560000 27.325000 ;
      RECT -4.730000 27.515000 -4.560000 27.685000 ;
      RECT -4.730000 27.875000 -4.560000 28.045000 ;
      RECT -4.730000 28.235000 -4.560000 28.405000 ;
      RECT -4.730000 28.595000 -4.560000 28.765000 ;
      RECT -4.730000 28.955000 -4.560000 29.125000 ;
      RECT -4.730000 29.315000 -4.560000 29.485000 ;
      RECT -4.730000 29.675000 -4.560000 29.845000 ;
      RECT -4.570000 -5.790000 -4.400000 -5.620000 ;
      RECT -4.570000 35.620000 -4.400000 35.790000 ;
      RECT -4.210000 -5.790000 -4.040000 -5.620000 ;
      RECT -4.210000 35.620000 -4.040000 35.790000 ;
      RECT -3.850000 -5.790000 -3.680000 -5.620000 ;
      RECT -3.850000 35.620000 -3.680000 35.790000 ;
      RECT -3.490000 -5.790000 -3.320000 -5.620000 ;
      RECT -3.490000 35.620000 -3.320000 35.790000 ;
      RECT -3.130000 -5.790000 -2.960000 -5.620000 ;
      RECT -3.130000 35.620000 -2.960000 35.790000 ;
      RECT -2.770000 -5.790000 -2.600000 -5.620000 ;
      RECT -2.770000 35.620000 -2.600000 35.790000 ;
      RECT -2.410000 -5.790000 -2.240000 -5.620000 ;
      RECT -2.410000 35.620000 -2.240000 35.790000 ;
      RECT -2.050000 -5.790000 -1.880000 -5.620000 ;
      RECT -2.050000 35.620000 -1.880000 35.790000 ;
      RECT -1.690000 -5.790000 -1.520000 -5.620000 ;
      RECT -1.690000 35.620000 -1.520000 35.790000 ;
      RECT -1.400000 -4.205000 -1.230000 -4.035000 ;
      RECT -1.400000 -3.835000 -1.230000 -3.665000 ;
      RECT -1.400000 -3.465000 -1.230000 -3.295000 ;
      RECT -1.330000 -5.790000 -1.160000 -5.620000 ;
      RECT -1.330000 35.620000 -1.160000 35.790000 ;
      RECT -1.030000 -4.205000 -0.860000 -4.035000 ;
      RECT -1.030000 -3.835000 -0.860000 -3.665000 ;
      RECT -1.030000 -3.465000 -0.860000 -3.295000 ;
      RECT -0.970000 -5.790000 -0.800000 -5.620000 ;
      RECT -0.970000 35.620000 -0.800000 35.790000 ;
      RECT -0.660000 -4.205000 -0.490000 -4.035000 ;
      RECT -0.660000 -3.835000 -0.490000 -3.665000 ;
      RECT -0.660000 -3.465000 -0.490000 -3.295000 ;
      RECT -0.610000 -5.790000 -0.440000 -5.620000 ;
      RECT -0.610000 35.620000 -0.440000 35.790000 ;
      RECT -0.290000 -4.205000 -0.120000 -4.035000 ;
      RECT -0.290000 -3.835000 -0.120000 -3.665000 ;
      RECT -0.290000 -3.465000 -0.120000 -3.295000 ;
      RECT -0.250000 -5.790000 -0.080000 -5.620000 ;
      RECT -0.250000 35.620000 -0.080000 35.790000 ;
      RECT  0.080000 -4.205000  0.250000 -4.035000 ;
      RECT  0.080000 -3.835000  0.250000 -3.665000 ;
      RECT  0.080000 -3.465000  0.250000 -3.295000 ;
      RECT  0.110000 -5.790000  0.280000 -5.620000 ;
      RECT  0.110000  0.335000  0.640000 29.665000 ;
      RECT  0.110000 35.620000  0.280000 35.790000 ;
      RECT  0.450000 -4.205000  0.620000 -4.035000 ;
      RECT  0.450000 -3.835000  0.620000 -3.665000 ;
      RECT  0.450000 -3.465000  0.620000 -3.295000 ;
      RECT  0.470000 -5.790000  0.640000 -5.620000 ;
      RECT  0.470000 35.620000  0.640000 35.790000 ;
      RECT  0.820000 -4.205000  0.990000 -4.035000 ;
      RECT  0.820000 -3.835000  0.990000 -3.665000 ;
      RECT  0.820000 -3.465000  0.990000 -3.295000 ;
      RECT  0.830000 -5.790000  1.000000 -5.620000 ;
      RECT  0.830000 35.620000  1.000000 35.790000 ;
      RECT  1.190000 -5.790000  1.360000 -5.620000 ;
      RECT  1.190000 -4.205000  1.360000 -4.035000 ;
      RECT  1.190000 -3.835000  1.360000 -3.665000 ;
      RECT  1.190000 -3.465000  1.360000 -3.295000 ;
      RECT  1.190000 35.620000  1.360000 35.790000 ;
      RECT  1.550000 -5.790000  1.720000 -5.620000 ;
      RECT  1.550000 35.620000  1.720000 35.790000 ;
      RECT  1.560000 -4.205000  1.730000 -4.035000 ;
      RECT  1.560000 -3.835000  1.730000 -3.665000 ;
      RECT  1.560000 -3.465000  1.730000 -3.295000 ;
      RECT  1.910000 -5.790000  2.080000 -5.620000 ;
      RECT  1.910000 35.620000  2.080000 35.790000 ;
      RECT  1.930000 -4.205000  2.100000 -4.035000 ;
      RECT  1.930000 -3.835000  2.100000 -3.665000 ;
      RECT  1.930000 -3.465000  2.100000 -3.295000 ;
      RECT  2.270000 -5.790000  2.440000 -5.620000 ;
      RECT  2.270000 35.620000  2.440000 35.790000 ;
      RECT  2.630000 -5.790000  2.800000 -5.620000 ;
      RECT  2.630000 35.620000  2.800000 35.790000 ;
      RECT  2.990000 -5.790000  3.160000 -5.620000 ;
      RECT  2.990000 35.620000  3.160000 35.790000 ;
      RECT  3.350000 -5.790000  3.520000 -5.620000 ;
      RECT  3.350000 35.620000  3.520000 35.790000 ;
      RECT  3.710000 -5.790000  3.880000 -5.620000 ;
      RECT  3.710000 35.620000  3.880000 35.790000 ;
      RECT  4.070000 -5.790000  4.240000 -5.620000 ;
      RECT  4.070000 35.620000  4.240000 35.790000 ;
      RECT  4.430000 -5.790000  4.600000 -5.620000 ;
      RECT  4.430000 35.620000  4.600000 35.790000 ;
      RECT  4.790000 -5.790000  4.960000 -5.620000 ;
      RECT  4.790000 35.620000  4.960000 35.790000 ;
      RECT  5.150000 -5.790000  5.320000 -5.620000 ;
      RECT  5.150000 35.620000  5.320000 35.790000 ;
      RECT  5.310000  0.155000  5.480000  0.325000 ;
      RECT  5.310000  0.515000  5.480000  0.685000 ;
      RECT  5.310000  0.875000  5.480000  1.045000 ;
      RECT  5.310000  1.235000  5.480000  1.405000 ;
      RECT  5.310000  1.595000  5.480000  1.765000 ;
      RECT  5.310000  1.955000  5.480000  2.125000 ;
      RECT  5.310000  2.315000  5.480000  2.485000 ;
      RECT  5.310000  2.675000  5.480000  2.845000 ;
      RECT  5.310000  3.035000  5.480000  3.205000 ;
      RECT  5.310000  3.395000  5.480000  3.565000 ;
      RECT  5.310000  3.755000  5.480000  3.925000 ;
      RECT  5.310000  4.115000  5.480000  4.285000 ;
      RECT  5.310000  4.475000  5.480000  4.645000 ;
      RECT  5.310000  4.835000  5.480000  5.005000 ;
      RECT  5.310000  5.195000  5.480000  5.365000 ;
      RECT  5.310000  5.555000  5.480000  5.725000 ;
      RECT  5.310000  5.915000  5.480000  6.085000 ;
      RECT  5.310000  6.275000  5.480000  6.445000 ;
      RECT  5.310000  6.635000  5.480000  6.805000 ;
      RECT  5.310000  6.995000  5.480000  7.165000 ;
      RECT  5.310000  7.355000  5.480000  7.525000 ;
      RECT  5.310000  7.715000  5.480000  7.885000 ;
      RECT  5.310000  8.075000  5.480000  8.245000 ;
      RECT  5.310000  8.435000  5.480000  8.605000 ;
      RECT  5.310000  8.795000  5.480000  8.965000 ;
      RECT  5.310000  9.155000  5.480000  9.325000 ;
      RECT  5.310000  9.515000  5.480000  9.685000 ;
      RECT  5.310000  9.875000  5.480000 10.045000 ;
      RECT  5.310000 10.235000  5.480000 10.405000 ;
      RECT  5.310000 10.595000  5.480000 10.765000 ;
      RECT  5.310000 10.955000  5.480000 11.125000 ;
      RECT  5.310000 11.315000  5.480000 11.485000 ;
      RECT  5.310000 11.675000  5.480000 11.845000 ;
      RECT  5.310000 12.035000  5.480000 12.205000 ;
      RECT  5.310000 12.395000  5.480000 12.565000 ;
      RECT  5.310000 12.755000  5.480000 12.925000 ;
      RECT  5.310000 13.115000  5.480000 13.285000 ;
      RECT  5.310000 13.475000  5.480000 13.645000 ;
      RECT  5.310000 13.835000  5.480000 14.005000 ;
      RECT  5.310000 14.195000  5.480000 14.365000 ;
      RECT  5.310000 14.555000  5.480000 14.725000 ;
      RECT  5.310000 14.915000  5.480000 15.085000 ;
      RECT  5.310000 15.275000  5.480000 15.445000 ;
      RECT  5.310000 15.635000  5.480000 15.805000 ;
      RECT  5.310000 15.995000  5.480000 16.165000 ;
      RECT  5.310000 16.355000  5.480000 16.525000 ;
      RECT  5.310000 16.715000  5.480000 16.885000 ;
      RECT  5.310000 17.075000  5.480000 17.245000 ;
      RECT  5.310000 17.435000  5.480000 17.605000 ;
      RECT  5.310000 17.795000  5.480000 17.965000 ;
      RECT  5.310000 18.155000  5.480000 18.325000 ;
      RECT  5.310000 18.515000  5.480000 18.685000 ;
      RECT  5.310000 18.875000  5.480000 19.045000 ;
      RECT  5.310000 19.235000  5.480000 19.405000 ;
      RECT  5.310000 19.595000  5.480000 19.765000 ;
      RECT  5.310000 19.955000  5.480000 20.125000 ;
      RECT  5.310000 20.315000  5.480000 20.485000 ;
      RECT  5.310000 20.675000  5.480000 20.845000 ;
      RECT  5.310000 21.035000  5.480000 21.205000 ;
      RECT  5.310000 21.395000  5.480000 21.565000 ;
      RECT  5.310000 21.755000  5.480000 21.925000 ;
      RECT  5.310000 22.115000  5.480000 22.285000 ;
      RECT  5.310000 22.475000  5.480000 22.645000 ;
      RECT  5.310000 22.835000  5.480000 23.005000 ;
      RECT  5.310000 23.195000  5.480000 23.365000 ;
      RECT  5.310000 23.555000  5.480000 23.725000 ;
      RECT  5.310000 23.915000  5.480000 24.085000 ;
      RECT  5.310000 24.275000  5.480000 24.445000 ;
      RECT  5.310000 24.635000  5.480000 24.805000 ;
      RECT  5.310000 24.995000  5.480000 25.165000 ;
      RECT  5.310000 25.355000  5.480000 25.525000 ;
      RECT  5.310000 25.715000  5.480000 25.885000 ;
      RECT  5.310000 26.075000  5.480000 26.245000 ;
      RECT  5.310000 26.435000  5.480000 26.605000 ;
      RECT  5.310000 26.795000  5.480000 26.965000 ;
      RECT  5.310000 27.155000  5.480000 27.325000 ;
      RECT  5.310000 27.515000  5.480000 27.685000 ;
      RECT  5.310000 27.875000  5.480000 28.045000 ;
      RECT  5.310000 28.235000  5.480000 28.405000 ;
      RECT  5.310000 28.595000  5.480000 28.765000 ;
      RECT  5.310000 28.955000  5.480000 29.125000 ;
      RECT  5.310000 29.315000  5.480000 29.485000 ;
      RECT  5.310000 29.675000  5.480000 29.845000 ;
      RECT  5.510000 -5.790000  5.680000 -5.620000 ;
      RECT  5.510000 35.620000  5.680000 35.790000 ;
      RECT  6.160000 -5.425000  6.330000 -5.255000 ;
      RECT  6.160000 -5.065000  6.330000 -4.895000 ;
      RECT  6.160000 -4.705000  6.330000 -4.535000 ;
      RECT  6.160000 -4.345000  6.330000 -4.175000 ;
      RECT  6.160000 -3.985000  6.330000 -3.815000 ;
      RECT  6.160000 -3.625000  6.330000 -3.455000 ;
      RECT  6.160000 -3.265000  6.330000 -3.095000 ;
      RECT  6.160000 -2.905000  6.330000 -2.735000 ;
      RECT  6.160000 -2.545000  6.330000 -2.375000 ;
      RECT  6.160000 -2.185000  6.330000 -2.015000 ;
      RECT  6.160000 -1.825000  6.330000 -1.655000 ;
      RECT  6.160000 -1.465000  6.330000 -1.295000 ;
      RECT  6.160000 -1.105000  6.330000 -0.935000 ;
      RECT  6.160000 -0.745000  6.330000 -0.575000 ;
      RECT  6.160000 -0.385000  6.330000 -0.215000 ;
      RECT  6.160000 -0.025000  6.330000  0.145000 ;
      RECT  6.160000  0.335000  6.330000  0.505000 ;
      RECT  6.160000  0.695000  6.330000  0.865000 ;
      RECT  6.160000  1.055000  6.330000  1.225000 ;
      RECT  6.160000  1.415000  6.330000  1.585000 ;
      RECT  6.160000  1.775000  6.330000  1.945000 ;
      RECT  6.160000  2.135000  6.330000  2.305000 ;
      RECT  6.160000  2.495000  6.330000  2.665000 ;
      RECT  6.160000  2.855000  6.330000  3.025000 ;
      RECT  6.160000  3.215000  6.330000  3.385000 ;
      RECT  6.160000  3.575000  6.330000  3.745000 ;
      RECT  6.160000  3.935000  6.330000  4.105000 ;
      RECT  6.160000  4.295000  6.330000  4.465000 ;
      RECT  6.160000  4.655000  6.330000  4.825000 ;
      RECT  6.160000  5.015000  6.330000  5.185000 ;
      RECT  6.160000  5.375000  6.330000  5.545000 ;
      RECT  6.160000  5.735000  6.330000  5.905000 ;
      RECT  6.160000  6.095000  6.330000  6.265000 ;
      RECT  6.160000  6.455000  6.330000  6.625000 ;
      RECT  6.160000  6.815000  6.330000  6.985000 ;
      RECT  6.160000  7.175000  6.330000  7.345000 ;
      RECT  6.160000  7.535000  6.330000  7.705000 ;
      RECT  6.160000  7.895000  6.330000  8.065000 ;
      RECT  6.160000  8.255000  6.330000  8.425000 ;
      RECT  6.160000  8.615000  6.330000  8.785000 ;
      RECT  6.160000  8.975000  6.330000  9.145000 ;
      RECT  6.160000  9.335000  6.330000  9.505000 ;
      RECT  6.160000  9.695000  6.330000  9.865000 ;
      RECT  6.160000 10.055000  6.330000 10.225000 ;
      RECT  6.160000 10.415000  6.330000 10.585000 ;
      RECT  6.160000 10.775000  6.330000 10.945000 ;
      RECT  6.160000 11.135000  6.330000 11.305000 ;
      RECT  6.160000 11.495000  6.330000 11.665000 ;
      RECT  6.160000 11.855000  6.330000 12.025000 ;
      RECT  6.160000 12.215000  6.330000 12.385000 ;
      RECT  6.160000 12.575000  6.330000 12.745000 ;
      RECT  6.160000 12.935000  6.330000 13.105000 ;
      RECT  6.160000 13.295000  6.330000 13.465000 ;
      RECT  6.160000 13.655000  6.330000 13.825000 ;
      RECT  6.160000 14.015000  6.330000 14.185000 ;
      RECT  6.160000 14.375000  6.330000 14.545000 ;
      RECT  6.160000 14.735000  6.330000 14.905000 ;
      RECT  6.160000 15.095000  6.330000 15.265000 ;
      RECT  6.160000 15.455000  6.330000 15.625000 ;
      RECT  6.160000 15.815000  6.330000 15.985000 ;
      RECT  6.160000 16.175000  6.330000 16.345000 ;
      RECT  6.160000 16.535000  6.330000 16.705000 ;
      RECT  6.160000 16.895000  6.330000 17.065000 ;
      RECT  6.160000 17.255000  6.330000 17.425000 ;
      RECT  6.160000 17.615000  6.330000 17.785000 ;
      RECT  6.160000 17.975000  6.330000 18.145000 ;
      RECT  6.160000 18.335000  6.330000 18.505000 ;
      RECT  6.160000 18.695000  6.330000 18.865000 ;
      RECT  6.160000 19.055000  6.330000 19.225000 ;
      RECT  6.160000 19.415000  6.330000 19.585000 ;
      RECT  6.160000 19.775000  6.330000 19.945000 ;
      RECT  6.160000 20.135000  6.330000 20.305000 ;
      RECT  6.160000 20.495000  6.330000 20.665000 ;
      RECT  6.160000 20.855000  6.330000 21.025000 ;
      RECT  6.160000 21.215000  6.330000 21.385000 ;
      RECT  6.160000 21.575000  6.330000 21.745000 ;
      RECT  6.160000 21.935000  6.330000 22.105000 ;
      RECT  6.160000 22.295000  6.330000 22.465000 ;
      RECT  6.160000 22.655000  6.330000 22.825000 ;
      RECT  6.160000 23.015000  6.330000 23.185000 ;
      RECT  6.160000 23.375000  6.330000 23.545000 ;
      RECT  6.160000 23.735000  6.330000 23.905000 ;
      RECT  6.160000 24.095000  6.330000 24.265000 ;
      RECT  6.160000 24.455000  6.330000 24.625000 ;
      RECT  6.160000 24.815000  6.330000 24.985000 ;
      RECT  6.160000 25.175000  6.330000 25.345000 ;
      RECT  6.160000 25.535000  6.330000 25.705000 ;
      RECT  6.160000 25.895000  6.330000 26.065000 ;
      RECT  6.160000 26.255000  6.330000 26.425000 ;
      RECT  6.160000 26.615000  6.330000 26.785000 ;
      RECT  6.160000 26.975000  6.330000 27.145000 ;
      RECT  6.160000 27.335000  6.330000 27.505000 ;
      RECT  6.160000 27.695000  6.330000 27.865000 ;
      RECT  6.160000 28.055000  6.330000 28.225000 ;
      RECT  6.160000 28.415000  6.330000 28.585000 ;
      RECT  6.160000 28.775000  6.330000 28.945000 ;
      RECT  6.160000 29.135000  6.330000 29.305000 ;
      RECT  6.160000 29.495000  6.330000 29.665000 ;
      RECT  6.160000 29.855000  6.330000 30.025000 ;
      RECT  6.160000 30.215000  6.330000 30.385000 ;
      RECT  6.160000 30.575000  6.330000 30.745000 ;
      RECT  6.160000 30.935000  6.330000 31.105000 ;
      RECT  6.160000 31.295000  6.330000 31.465000 ;
      RECT  6.160000 31.655000  6.330000 31.825000 ;
      RECT  6.160000 32.015000  6.330000 32.185000 ;
      RECT  6.160000 32.375000  6.330000 32.545000 ;
      RECT  6.160000 32.735000  6.330000 32.905000 ;
      RECT  6.160000 33.095000  6.330000 33.265000 ;
      RECT  6.160000 33.455000  6.330000 33.625000 ;
      RECT  6.160000 33.815000  6.330000 33.985000 ;
      RECT  6.160000 34.175000  6.330000 34.345000 ;
      RECT  6.160000 34.535000  6.330000 34.705000 ;
      RECT  6.160000 34.895000  6.330000 35.065000 ;
      RECT  6.160000 35.255000  6.330000 35.425000 ;
    LAYER met1 ;
      RECT -5.700000 -5.910000  6.450000 -5.500000 ;
      RECT -5.700000 -5.500000 -5.290000 35.500000 ;
      RECT -5.700000 35.500000  6.450000 35.910000 ;
      RECT -4.790000  0.095000 -4.500000 29.905000 ;
      RECT -1.480000 -4.285000  2.300000 -3.215000 ;
      RECT  0.050000  0.275000  0.700000 29.725000 ;
      RECT  5.250000  0.095000  5.540000 29.905000 ;
      RECT  6.040000 -5.500000  6.450000 35.500000 ;
    LAYER met2 ;
      RECT -1.480000 -4.285000 2.300000 -3.215000 ;
      RECT  0.055000  0.285000 0.695000 29.725000 ;
    LAYER via ;
      RECT -1.445000 -4.250000 -1.185000 -3.990000 ;
      RECT -1.445000 -3.880000 -1.185000 -3.620000 ;
      RECT -1.445000 -3.510000 -1.185000 -3.250000 ;
      RECT -1.075000 -4.250000 -0.815000 -3.990000 ;
      RECT -1.075000 -3.880000 -0.815000 -3.620000 ;
      RECT -1.075000 -3.510000 -0.815000 -3.250000 ;
      RECT -0.705000 -4.250000 -0.445000 -3.990000 ;
      RECT -0.705000 -3.880000 -0.445000 -3.620000 ;
      RECT -0.705000 -3.510000 -0.445000 -3.250000 ;
      RECT -0.335000 -4.250000 -0.075000 -3.990000 ;
      RECT -0.335000 -3.880000 -0.075000 -3.620000 ;
      RECT -0.335000 -3.510000 -0.075000 -3.250000 ;
      RECT  0.035000 -4.250000  0.295000 -3.990000 ;
      RECT  0.035000 -3.880000  0.295000 -3.620000 ;
      RECT  0.035000 -3.510000  0.295000 -3.250000 ;
      RECT  0.085000  0.315000  0.665000 29.695000 ;
      RECT  0.405000 -4.250000  0.665000 -3.990000 ;
      RECT  0.405000 -3.880000  0.665000 -3.620000 ;
      RECT  0.405000 -3.510000  0.665000 -3.250000 ;
      RECT  0.775000 -4.250000  1.035000 -3.990000 ;
      RECT  0.775000 -3.880000  1.035000 -3.620000 ;
      RECT  0.775000 -3.510000  1.035000 -3.250000 ;
      RECT  1.145000 -4.250000  1.405000 -3.990000 ;
      RECT  1.145000 -3.880000  1.405000 -3.620000 ;
      RECT  1.145000 -3.510000  1.405000 -3.250000 ;
      RECT  1.515000 -4.250000  1.775000 -3.990000 ;
      RECT  1.515000 -3.880000  1.775000 -3.620000 ;
      RECT  1.515000 -3.510000  1.775000 -3.250000 ;
      RECT  1.885000 -4.250000  2.145000 -3.990000 ;
      RECT  1.885000 -3.880000  2.145000 -3.620000 ;
      RECT  1.885000 -3.510000  2.145000 -3.250000 ;
  END
END sky130_fd_pr__rf_nfet_20v0_withptap
END LIBRARY
