* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
*
* model corner
* , Bin 000, W = 30.0, L = 1.0
* ----------------------------
.param
+ sky130_fd_pr__nfet_20v0_nvt_iso__rdrift_mult = 1.8311e+0
+ sky130_fd_pr__nfet_20v0_nvt_iso__hvvsat_mult = 1.2679e+0
+ sky130_fd_pr__nfet_20v0_nvt_iso__vth0_diff = 1.4649e-1
+ sky130_fd_pr__nfet_20v0_nvt_iso__k2_diff = -1.1937e-1
.include "sky130_fd_pr__nfet_20v0_nvt_iso__subcircuit.pm3.spice"
