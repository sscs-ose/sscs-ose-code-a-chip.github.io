* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__res_generic_pd t1 t2 b
+ w=1 l=1
r0 t1 t2 sky130_fd_pr__res_generic_pd w = {w} l = {l}
d0 t1 b sky130_fd_pr__model__parasitic__diode_ps2nw area = 'w*l*0.5' pj = 'w+l'
d1 t2 b sky130_fd_pr__model__parasitic__diode_ps2nw area = 'w*l*0.5' pj = 'w+l'
.ends sky130_fd_pr__res_generic_pd
