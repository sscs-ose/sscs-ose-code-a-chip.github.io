# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p15 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  3.010000 BY  6.940000 ;
  PIN DRAIN
    ANTENNADIFFAREA  1.414000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 3.595000 3.080000 5.955000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.515000 ;
    PORT
      LAYER li1 ;
        RECT 1.240000 0.000000 1.910000 0.695000 ;
        RECT 1.240000 6.245000 1.910000 6.940000 ;
      LAYER mcon ;
        RECT 1.310000 0.095000 1.840000 0.625000 ;
        RECT 1.310000 6.315000 1.840000 6.845000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.250000 0.000000 1.900000 0.685000 ;
        RECT 1.250000 6.255000 1.900000 6.940000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 0.985000 3.080000 3.345000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  3.282500 ;
    ANTENNAGATEAREA  0.757500 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 0.985000 0.500000 5.955000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.650000 0.985000 2.945000 5.955000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 0.800000 6.015000 ;
      RECT 0.600000 0.485000 0.930000 0.815000 ;
      RECT 0.600000 0.815000 0.800000 0.925000 ;
      RECT 0.600000 6.015000 0.800000 6.125000 ;
      RECT 0.600000 6.125000 0.930000 6.455000 ;
      RECT 1.060000 0.925000 1.230000 6.015000 ;
      RECT 1.490000 0.925000 1.660000 6.015000 ;
      RECT 1.920000 0.925000 2.090000 6.015000 ;
      RECT 2.220000 0.485000 2.550000 0.815000 ;
      RECT 2.220000 6.125000 2.550000 6.455000 ;
      RECT 2.350000 0.815000 2.550000 0.925000 ;
      RECT 2.350000 0.925000 2.945000 6.015000 ;
      RECT 2.350000 6.015000 2.550000 6.125000 ;
    LAYER mcon ;
      RECT 0.300000 1.045000 0.470000 1.215000 ;
      RECT 0.300000 1.405000 0.470000 1.575000 ;
      RECT 0.300000 1.765000 0.470000 1.935000 ;
      RECT 0.300000 2.125000 0.470000 2.295000 ;
      RECT 0.300000 2.485000 0.470000 2.655000 ;
      RECT 0.300000 2.845000 0.470000 3.015000 ;
      RECT 0.300000 3.205000 0.470000 3.375000 ;
      RECT 0.300000 3.565000 0.470000 3.735000 ;
      RECT 0.300000 3.925000 0.470000 4.095000 ;
      RECT 0.300000 4.285000 0.470000 4.455000 ;
      RECT 0.300000 4.645000 0.470000 4.815000 ;
      RECT 0.300000 5.005000 0.470000 5.175000 ;
      RECT 0.300000 5.365000 0.470000 5.535000 ;
      RECT 0.300000 5.725000 0.470000 5.895000 ;
      RECT 1.060000 1.045000 1.230000 1.215000 ;
      RECT 1.060000 1.405000 1.230000 1.575000 ;
      RECT 1.060000 1.765000 1.230000 1.935000 ;
      RECT 1.060000 2.125000 1.230000 2.295000 ;
      RECT 1.060000 2.485000 1.230000 2.655000 ;
      RECT 1.060000 2.845000 1.230000 3.015000 ;
      RECT 1.060000 3.205000 1.230000 3.375000 ;
      RECT 1.060000 3.565000 1.230000 3.735000 ;
      RECT 1.060000 3.925000 1.230000 4.095000 ;
      RECT 1.060000 4.285000 1.230000 4.455000 ;
      RECT 1.060000 4.645000 1.230000 4.815000 ;
      RECT 1.060000 5.005000 1.230000 5.175000 ;
      RECT 1.060000 5.365000 1.230000 5.535000 ;
      RECT 1.060000 5.725000 1.230000 5.895000 ;
      RECT 1.490000 1.045000 1.660000 1.215000 ;
      RECT 1.490000 1.405000 1.660000 1.575000 ;
      RECT 1.490000 1.765000 1.660000 1.935000 ;
      RECT 1.490000 2.125000 1.660000 2.295000 ;
      RECT 1.490000 2.485000 1.660000 2.655000 ;
      RECT 1.490000 2.845000 1.660000 3.015000 ;
      RECT 1.490000 3.205000 1.660000 3.375000 ;
      RECT 1.490000 3.565000 1.660000 3.735000 ;
      RECT 1.490000 3.925000 1.660000 4.095000 ;
      RECT 1.490000 4.285000 1.660000 4.455000 ;
      RECT 1.490000 4.645000 1.660000 4.815000 ;
      RECT 1.490000 5.005000 1.660000 5.175000 ;
      RECT 1.490000 5.365000 1.660000 5.535000 ;
      RECT 1.490000 5.725000 1.660000 5.895000 ;
      RECT 1.920000 1.045000 2.090000 1.215000 ;
      RECT 1.920000 1.405000 2.090000 1.575000 ;
      RECT 1.920000 1.765000 2.090000 1.935000 ;
      RECT 1.920000 2.125000 2.090000 2.295000 ;
      RECT 1.920000 2.485000 2.090000 2.655000 ;
      RECT 1.920000 2.845000 2.090000 3.015000 ;
      RECT 1.920000 3.205000 2.090000 3.375000 ;
      RECT 1.920000 3.565000 2.090000 3.735000 ;
      RECT 1.920000 3.925000 2.090000 4.095000 ;
      RECT 1.920000 4.285000 2.090000 4.455000 ;
      RECT 1.920000 4.645000 2.090000 4.815000 ;
      RECT 1.920000 5.005000 2.090000 5.175000 ;
      RECT 1.920000 5.365000 2.090000 5.535000 ;
      RECT 1.920000 5.725000 2.090000 5.895000 ;
      RECT 2.680000 1.045000 2.850000 1.215000 ;
      RECT 2.680000 1.405000 2.850000 1.575000 ;
      RECT 2.680000 1.765000 2.850000 1.935000 ;
      RECT 2.680000 2.125000 2.850000 2.295000 ;
      RECT 2.680000 2.485000 2.850000 2.655000 ;
      RECT 2.680000 2.845000 2.850000 3.015000 ;
      RECT 2.680000 3.205000 2.850000 3.375000 ;
      RECT 2.680000 3.565000 2.850000 3.735000 ;
      RECT 2.680000 3.925000 2.850000 4.095000 ;
      RECT 2.680000 4.285000 2.850000 4.455000 ;
      RECT 2.680000 4.645000 2.850000 4.815000 ;
      RECT 2.680000 5.005000 2.850000 5.175000 ;
      RECT 2.680000 5.365000 2.850000 5.535000 ;
      RECT 2.680000 5.725000 2.850000 5.895000 ;
    LAYER met1 ;
      RECT 1.015000 0.985000 1.275000 5.955000 ;
      RECT 1.445000 0.985000 1.705000 5.955000 ;
      RECT 1.875000 0.985000 2.135000 5.955000 ;
    LAYER via ;
      RECT 1.015000 1.015000 1.275000 1.275000 ;
      RECT 1.015000 1.335000 1.275000 1.595000 ;
      RECT 1.015000 1.655000 1.275000 1.915000 ;
      RECT 1.015000 1.975000 1.275000 2.235000 ;
      RECT 1.015000 2.295000 1.275000 2.555000 ;
      RECT 1.015000 2.615000 1.275000 2.875000 ;
      RECT 1.015000 2.935000 1.275000 3.195000 ;
      RECT 1.445000 3.745000 1.705000 4.005000 ;
      RECT 1.445000 4.065000 1.705000 4.325000 ;
      RECT 1.445000 4.385000 1.705000 4.645000 ;
      RECT 1.445000 4.705000 1.705000 4.965000 ;
      RECT 1.445000 5.025000 1.705000 5.285000 ;
      RECT 1.445000 5.345000 1.705000 5.605000 ;
      RECT 1.445000 5.665000 1.705000 5.925000 ;
      RECT 1.875000 1.015000 2.135000 1.275000 ;
      RECT 1.875000 1.335000 2.135000 1.595000 ;
      RECT 1.875000 1.655000 2.135000 1.915000 ;
      RECT 1.875000 1.975000 2.135000 2.235000 ;
      RECT 1.875000 2.295000 2.135000 2.555000 ;
      RECT 1.875000 2.615000 2.135000 2.875000 ;
      RECT 1.875000 2.935000 2.135000 3.195000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p15
END LIBRARY
