MACRO DCL_NMOS_S_55663590_X148_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_55663590_X148_Y1 0 0 ;
  SIZE 129000 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64360 260 64640 4780 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64790 680 65070 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 7225 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 7225 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 7225 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 7225 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 7225 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 7225 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 7225 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 7225 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 7225 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 7225 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 7225 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 7225 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 7225 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 7225 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 7225 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 7225 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 7225 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 7225 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 7225 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 20085 335 20335 3865 ;
    LAYER M1 ;
      RECT 20085 4115 20335 5125 ;
    LAYER M1 ;
      RECT 20085 6215 20335 7225 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20945 335 21195 3865 ;
    LAYER M1 ;
      RECT 20945 4115 21195 5125 ;
    LAYER M1 ;
      RECT 20945 6215 21195 7225 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 21805 335 22055 3865 ;
    LAYER M1 ;
      RECT 21805 4115 22055 5125 ;
    LAYER M1 ;
      RECT 21805 6215 22055 7225 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22665 335 22915 3865 ;
    LAYER M1 ;
      RECT 22665 4115 22915 5125 ;
    LAYER M1 ;
      RECT 22665 6215 22915 7225 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23525 335 23775 3865 ;
    LAYER M1 ;
      RECT 23525 4115 23775 5125 ;
    LAYER M1 ;
      RECT 23525 6215 23775 7225 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 24385 335 24635 3865 ;
    LAYER M1 ;
      RECT 24385 4115 24635 5125 ;
    LAYER M1 ;
      RECT 24385 6215 24635 7225 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M1 ;
      RECT 25245 335 25495 3865 ;
    LAYER M1 ;
      RECT 25245 4115 25495 5125 ;
    LAYER M1 ;
      RECT 25245 6215 25495 7225 ;
    LAYER M1 ;
      RECT 25675 335 25925 3865 ;
    LAYER M1 ;
      RECT 26105 335 26355 3865 ;
    LAYER M1 ;
      RECT 26105 4115 26355 5125 ;
    LAYER M1 ;
      RECT 26105 6215 26355 7225 ;
    LAYER M1 ;
      RECT 26535 335 26785 3865 ;
    LAYER M1 ;
      RECT 26965 335 27215 3865 ;
    LAYER M1 ;
      RECT 26965 4115 27215 5125 ;
    LAYER M1 ;
      RECT 26965 6215 27215 7225 ;
    LAYER M1 ;
      RECT 27395 335 27645 3865 ;
    LAYER M1 ;
      RECT 27825 335 28075 3865 ;
    LAYER M1 ;
      RECT 27825 4115 28075 5125 ;
    LAYER M1 ;
      RECT 27825 6215 28075 7225 ;
    LAYER M1 ;
      RECT 28255 335 28505 3865 ;
    LAYER M1 ;
      RECT 28685 335 28935 3865 ;
    LAYER M1 ;
      RECT 28685 4115 28935 5125 ;
    LAYER M1 ;
      RECT 28685 6215 28935 7225 ;
    LAYER M1 ;
      RECT 29115 335 29365 3865 ;
    LAYER M1 ;
      RECT 29545 335 29795 3865 ;
    LAYER M1 ;
      RECT 29545 4115 29795 5125 ;
    LAYER M1 ;
      RECT 29545 6215 29795 7225 ;
    LAYER M1 ;
      RECT 29975 335 30225 3865 ;
    LAYER M1 ;
      RECT 30405 335 30655 3865 ;
    LAYER M1 ;
      RECT 30405 4115 30655 5125 ;
    LAYER M1 ;
      RECT 30405 6215 30655 7225 ;
    LAYER M1 ;
      RECT 30835 335 31085 3865 ;
    LAYER M1 ;
      RECT 31265 335 31515 3865 ;
    LAYER M1 ;
      RECT 31265 4115 31515 5125 ;
    LAYER M1 ;
      RECT 31265 6215 31515 7225 ;
    LAYER M1 ;
      RECT 31695 335 31945 3865 ;
    LAYER M1 ;
      RECT 32125 335 32375 3865 ;
    LAYER M1 ;
      RECT 32125 4115 32375 5125 ;
    LAYER M1 ;
      RECT 32125 6215 32375 7225 ;
    LAYER M1 ;
      RECT 32555 335 32805 3865 ;
    LAYER M1 ;
      RECT 32985 335 33235 3865 ;
    LAYER M1 ;
      RECT 32985 4115 33235 5125 ;
    LAYER M1 ;
      RECT 32985 6215 33235 7225 ;
    LAYER M1 ;
      RECT 33415 335 33665 3865 ;
    LAYER M1 ;
      RECT 33845 335 34095 3865 ;
    LAYER M1 ;
      RECT 33845 4115 34095 5125 ;
    LAYER M1 ;
      RECT 33845 6215 34095 7225 ;
    LAYER M1 ;
      RECT 34275 335 34525 3865 ;
    LAYER M1 ;
      RECT 34705 335 34955 3865 ;
    LAYER M1 ;
      RECT 34705 4115 34955 5125 ;
    LAYER M1 ;
      RECT 34705 6215 34955 7225 ;
    LAYER M1 ;
      RECT 35135 335 35385 3865 ;
    LAYER M1 ;
      RECT 35565 335 35815 3865 ;
    LAYER M1 ;
      RECT 35565 4115 35815 5125 ;
    LAYER M1 ;
      RECT 35565 6215 35815 7225 ;
    LAYER M1 ;
      RECT 35995 335 36245 3865 ;
    LAYER M1 ;
      RECT 36425 335 36675 3865 ;
    LAYER M1 ;
      RECT 36425 4115 36675 5125 ;
    LAYER M1 ;
      RECT 36425 6215 36675 7225 ;
    LAYER M1 ;
      RECT 36855 335 37105 3865 ;
    LAYER M1 ;
      RECT 37285 335 37535 3865 ;
    LAYER M1 ;
      RECT 37285 4115 37535 5125 ;
    LAYER M1 ;
      RECT 37285 6215 37535 7225 ;
    LAYER M1 ;
      RECT 37715 335 37965 3865 ;
    LAYER M1 ;
      RECT 38145 335 38395 3865 ;
    LAYER M1 ;
      RECT 38145 4115 38395 5125 ;
    LAYER M1 ;
      RECT 38145 6215 38395 7225 ;
    LAYER M1 ;
      RECT 38575 335 38825 3865 ;
    LAYER M1 ;
      RECT 39005 335 39255 3865 ;
    LAYER M1 ;
      RECT 39005 4115 39255 5125 ;
    LAYER M1 ;
      RECT 39005 6215 39255 7225 ;
    LAYER M1 ;
      RECT 39435 335 39685 3865 ;
    LAYER M1 ;
      RECT 39865 335 40115 3865 ;
    LAYER M1 ;
      RECT 39865 4115 40115 5125 ;
    LAYER M1 ;
      RECT 39865 6215 40115 7225 ;
    LAYER M1 ;
      RECT 40295 335 40545 3865 ;
    LAYER M1 ;
      RECT 40725 335 40975 3865 ;
    LAYER M1 ;
      RECT 40725 4115 40975 5125 ;
    LAYER M1 ;
      RECT 40725 6215 40975 7225 ;
    LAYER M1 ;
      RECT 41155 335 41405 3865 ;
    LAYER M1 ;
      RECT 41585 335 41835 3865 ;
    LAYER M1 ;
      RECT 41585 4115 41835 5125 ;
    LAYER M1 ;
      RECT 41585 6215 41835 7225 ;
    LAYER M1 ;
      RECT 42015 335 42265 3865 ;
    LAYER M1 ;
      RECT 42445 335 42695 3865 ;
    LAYER M1 ;
      RECT 42445 4115 42695 5125 ;
    LAYER M1 ;
      RECT 42445 6215 42695 7225 ;
    LAYER M1 ;
      RECT 42875 335 43125 3865 ;
    LAYER M1 ;
      RECT 43305 335 43555 3865 ;
    LAYER M1 ;
      RECT 43305 4115 43555 5125 ;
    LAYER M1 ;
      RECT 43305 6215 43555 7225 ;
    LAYER M1 ;
      RECT 43735 335 43985 3865 ;
    LAYER M1 ;
      RECT 44165 335 44415 3865 ;
    LAYER M1 ;
      RECT 44165 4115 44415 5125 ;
    LAYER M1 ;
      RECT 44165 6215 44415 7225 ;
    LAYER M1 ;
      RECT 44595 335 44845 3865 ;
    LAYER M1 ;
      RECT 45025 335 45275 3865 ;
    LAYER M1 ;
      RECT 45025 4115 45275 5125 ;
    LAYER M1 ;
      RECT 45025 6215 45275 7225 ;
    LAYER M1 ;
      RECT 45455 335 45705 3865 ;
    LAYER M1 ;
      RECT 45885 335 46135 3865 ;
    LAYER M1 ;
      RECT 45885 4115 46135 5125 ;
    LAYER M1 ;
      RECT 45885 6215 46135 7225 ;
    LAYER M1 ;
      RECT 46315 335 46565 3865 ;
    LAYER M1 ;
      RECT 46745 335 46995 3865 ;
    LAYER M1 ;
      RECT 46745 4115 46995 5125 ;
    LAYER M1 ;
      RECT 46745 6215 46995 7225 ;
    LAYER M1 ;
      RECT 47175 335 47425 3865 ;
    LAYER M1 ;
      RECT 47605 335 47855 3865 ;
    LAYER M1 ;
      RECT 47605 4115 47855 5125 ;
    LAYER M1 ;
      RECT 47605 6215 47855 7225 ;
    LAYER M1 ;
      RECT 48035 335 48285 3865 ;
    LAYER M1 ;
      RECT 48465 335 48715 3865 ;
    LAYER M1 ;
      RECT 48465 4115 48715 5125 ;
    LAYER M1 ;
      RECT 48465 6215 48715 7225 ;
    LAYER M1 ;
      RECT 48895 335 49145 3865 ;
    LAYER M1 ;
      RECT 49325 335 49575 3865 ;
    LAYER M1 ;
      RECT 49325 4115 49575 5125 ;
    LAYER M1 ;
      RECT 49325 6215 49575 7225 ;
    LAYER M1 ;
      RECT 49755 335 50005 3865 ;
    LAYER M1 ;
      RECT 50185 335 50435 3865 ;
    LAYER M1 ;
      RECT 50185 4115 50435 5125 ;
    LAYER M1 ;
      RECT 50185 6215 50435 7225 ;
    LAYER M1 ;
      RECT 50615 335 50865 3865 ;
    LAYER M1 ;
      RECT 51045 335 51295 3865 ;
    LAYER M1 ;
      RECT 51045 4115 51295 5125 ;
    LAYER M1 ;
      RECT 51045 6215 51295 7225 ;
    LAYER M1 ;
      RECT 51475 335 51725 3865 ;
    LAYER M1 ;
      RECT 51905 335 52155 3865 ;
    LAYER M1 ;
      RECT 51905 4115 52155 5125 ;
    LAYER M1 ;
      RECT 51905 6215 52155 7225 ;
    LAYER M1 ;
      RECT 52335 335 52585 3865 ;
    LAYER M1 ;
      RECT 52765 335 53015 3865 ;
    LAYER M1 ;
      RECT 52765 4115 53015 5125 ;
    LAYER M1 ;
      RECT 52765 6215 53015 7225 ;
    LAYER M1 ;
      RECT 53195 335 53445 3865 ;
    LAYER M1 ;
      RECT 53625 335 53875 3865 ;
    LAYER M1 ;
      RECT 53625 4115 53875 5125 ;
    LAYER M1 ;
      RECT 53625 6215 53875 7225 ;
    LAYER M1 ;
      RECT 54055 335 54305 3865 ;
    LAYER M1 ;
      RECT 54485 335 54735 3865 ;
    LAYER M1 ;
      RECT 54485 4115 54735 5125 ;
    LAYER M1 ;
      RECT 54485 6215 54735 7225 ;
    LAYER M1 ;
      RECT 54915 335 55165 3865 ;
    LAYER M1 ;
      RECT 55345 335 55595 3865 ;
    LAYER M1 ;
      RECT 55345 4115 55595 5125 ;
    LAYER M1 ;
      RECT 55345 6215 55595 7225 ;
    LAYER M1 ;
      RECT 55775 335 56025 3865 ;
    LAYER M1 ;
      RECT 56205 335 56455 3865 ;
    LAYER M1 ;
      RECT 56205 4115 56455 5125 ;
    LAYER M1 ;
      RECT 56205 6215 56455 7225 ;
    LAYER M1 ;
      RECT 56635 335 56885 3865 ;
    LAYER M1 ;
      RECT 57065 335 57315 3865 ;
    LAYER M1 ;
      RECT 57065 4115 57315 5125 ;
    LAYER M1 ;
      RECT 57065 6215 57315 7225 ;
    LAYER M1 ;
      RECT 57495 335 57745 3865 ;
    LAYER M1 ;
      RECT 57925 335 58175 3865 ;
    LAYER M1 ;
      RECT 57925 4115 58175 5125 ;
    LAYER M1 ;
      RECT 57925 6215 58175 7225 ;
    LAYER M1 ;
      RECT 58355 335 58605 3865 ;
    LAYER M1 ;
      RECT 58785 335 59035 3865 ;
    LAYER M1 ;
      RECT 58785 4115 59035 5125 ;
    LAYER M1 ;
      RECT 58785 6215 59035 7225 ;
    LAYER M1 ;
      RECT 59215 335 59465 3865 ;
    LAYER M1 ;
      RECT 59645 335 59895 3865 ;
    LAYER M1 ;
      RECT 59645 4115 59895 5125 ;
    LAYER M1 ;
      RECT 59645 6215 59895 7225 ;
    LAYER M1 ;
      RECT 60075 335 60325 3865 ;
    LAYER M1 ;
      RECT 60505 335 60755 3865 ;
    LAYER M1 ;
      RECT 60505 4115 60755 5125 ;
    LAYER M1 ;
      RECT 60505 6215 60755 7225 ;
    LAYER M1 ;
      RECT 60935 335 61185 3865 ;
    LAYER M1 ;
      RECT 61365 335 61615 3865 ;
    LAYER M1 ;
      RECT 61365 4115 61615 5125 ;
    LAYER M1 ;
      RECT 61365 6215 61615 7225 ;
    LAYER M1 ;
      RECT 61795 335 62045 3865 ;
    LAYER M1 ;
      RECT 62225 335 62475 3865 ;
    LAYER M1 ;
      RECT 62225 4115 62475 5125 ;
    LAYER M1 ;
      RECT 62225 6215 62475 7225 ;
    LAYER M1 ;
      RECT 62655 335 62905 3865 ;
    LAYER M1 ;
      RECT 63085 335 63335 3865 ;
    LAYER M1 ;
      RECT 63085 4115 63335 5125 ;
    LAYER M1 ;
      RECT 63085 6215 63335 7225 ;
    LAYER M1 ;
      RECT 63515 335 63765 3865 ;
    LAYER M1 ;
      RECT 63945 335 64195 3865 ;
    LAYER M1 ;
      RECT 63945 4115 64195 5125 ;
    LAYER M1 ;
      RECT 63945 6215 64195 7225 ;
    LAYER M1 ;
      RECT 64375 335 64625 3865 ;
    LAYER M1 ;
      RECT 64805 335 65055 3865 ;
    LAYER M1 ;
      RECT 64805 4115 65055 5125 ;
    LAYER M1 ;
      RECT 64805 6215 65055 7225 ;
    LAYER M1 ;
      RECT 65235 335 65485 3865 ;
    LAYER M1 ;
      RECT 65665 335 65915 3865 ;
    LAYER M1 ;
      RECT 65665 4115 65915 5125 ;
    LAYER M1 ;
      RECT 65665 6215 65915 7225 ;
    LAYER M1 ;
      RECT 66095 335 66345 3865 ;
    LAYER M1 ;
      RECT 66525 335 66775 3865 ;
    LAYER M1 ;
      RECT 66525 4115 66775 5125 ;
    LAYER M1 ;
      RECT 66525 6215 66775 7225 ;
    LAYER M1 ;
      RECT 66955 335 67205 3865 ;
    LAYER M1 ;
      RECT 67385 335 67635 3865 ;
    LAYER M1 ;
      RECT 67385 4115 67635 5125 ;
    LAYER M1 ;
      RECT 67385 6215 67635 7225 ;
    LAYER M1 ;
      RECT 67815 335 68065 3865 ;
    LAYER M1 ;
      RECT 68245 335 68495 3865 ;
    LAYER M1 ;
      RECT 68245 4115 68495 5125 ;
    LAYER M1 ;
      RECT 68245 6215 68495 7225 ;
    LAYER M1 ;
      RECT 68675 335 68925 3865 ;
    LAYER M1 ;
      RECT 69105 335 69355 3865 ;
    LAYER M1 ;
      RECT 69105 4115 69355 5125 ;
    LAYER M1 ;
      RECT 69105 6215 69355 7225 ;
    LAYER M1 ;
      RECT 69535 335 69785 3865 ;
    LAYER M1 ;
      RECT 69965 335 70215 3865 ;
    LAYER M1 ;
      RECT 69965 4115 70215 5125 ;
    LAYER M1 ;
      RECT 69965 6215 70215 7225 ;
    LAYER M1 ;
      RECT 70395 335 70645 3865 ;
    LAYER M1 ;
      RECT 70825 335 71075 3865 ;
    LAYER M1 ;
      RECT 70825 4115 71075 5125 ;
    LAYER M1 ;
      RECT 70825 6215 71075 7225 ;
    LAYER M1 ;
      RECT 71255 335 71505 3865 ;
    LAYER M1 ;
      RECT 71685 335 71935 3865 ;
    LAYER M1 ;
      RECT 71685 4115 71935 5125 ;
    LAYER M1 ;
      RECT 71685 6215 71935 7225 ;
    LAYER M1 ;
      RECT 72115 335 72365 3865 ;
    LAYER M1 ;
      RECT 72545 335 72795 3865 ;
    LAYER M1 ;
      RECT 72545 4115 72795 5125 ;
    LAYER M1 ;
      RECT 72545 6215 72795 7225 ;
    LAYER M1 ;
      RECT 72975 335 73225 3865 ;
    LAYER M1 ;
      RECT 73405 335 73655 3865 ;
    LAYER M1 ;
      RECT 73405 4115 73655 5125 ;
    LAYER M1 ;
      RECT 73405 6215 73655 7225 ;
    LAYER M1 ;
      RECT 73835 335 74085 3865 ;
    LAYER M1 ;
      RECT 74265 335 74515 3865 ;
    LAYER M1 ;
      RECT 74265 4115 74515 5125 ;
    LAYER M1 ;
      RECT 74265 6215 74515 7225 ;
    LAYER M1 ;
      RECT 74695 335 74945 3865 ;
    LAYER M1 ;
      RECT 75125 335 75375 3865 ;
    LAYER M1 ;
      RECT 75125 4115 75375 5125 ;
    LAYER M1 ;
      RECT 75125 6215 75375 7225 ;
    LAYER M1 ;
      RECT 75555 335 75805 3865 ;
    LAYER M1 ;
      RECT 75985 335 76235 3865 ;
    LAYER M1 ;
      RECT 75985 4115 76235 5125 ;
    LAYER M1 ;
      RECT 75985 6215 76235 7225 ;
    LAYER M1 ;
      RECT 76415 335 76665 3865 ;
    LAYER M1 ;
      RECT 76845 335 77095 3865 ;
    LAYER M1 ;
      RECT 76845 4115 77095 5125 ;
    LAYER M1 ;
      RECT 76845 6215 77095 7225 ;
    LAYER M1 ;
      RECT 77275 335 77525 3865 ;
    LAYER M1 ;
      RECT 77705 335 77955 3865 ;
    LAYER M1 ;
      RECT 77705 4115 77955 5125 ;
    LAYER M1 ;
      RECT 77705 6215 77955 7225 ;
    LAYER M1 ;
      RECT 78135 335 78385 3865 ;
    LAYER M1 ;
      RECT 78565 335 78815 3865 ;
    LAYER M1 ;
      RECT 78565 4115 78815 5125 ;
    LAYER M1 ;
      RECT 78565 6215 78815 7225 ;
    LAYER M1 ;
      RECT 78995 335 79245 3865 ;
    LAYER M1 ;
      RECT 79425 335 79675 3865 ;
    LAYER M1 ;
      RECT 79425 4115 79675 5125 ;
    LAYER M1 ;
      RECT 79425 6215 79675 7225 ;
    LAYER M1 ;
      RECT 79855 335 80105 3865 ;
    LAYER M1 ;
      RECT 80285 335 80535 3865 ;
    LAYER M1 ;
      RECT 80285 4115 80535 5125 ;
    LAYER M1 ;
      RECT 80285 6215 80535 7225 ;
    LAYER M1 ;
      RECT 80715 335 80965 3865 ;
    LAYER M1 ;
      RECT 81145 335 81395 3865 ;
    LAYER M1 ;
      RECT 81145 4115 81395 5125 ;
    LAYER M1 ;
      RECT 81145 6215 81395 7225 ;
    LAYER M1 ;
      RECT 81575 335 81825 3865 ;
    LAYER M1 ;
      RECT 82005 335 82255 3865 ;
    LAYER M1 ;
      RECT 82005 4115 82255 5125 ;
    LAYER M1 ;
      RECT 82005 6215 82255 7225 ;
    LAYER M1 ;
      RECT 82435 335 82685 3865 ;
    LAYER M1 ;
      RECT 82865 335 83115 3865 ;
    LAYER M1 ;
      RECT 82865 4115 83115 5125 ;
    LAYER M1 ;
      RECT 82865 6215 83115 7225 ;
    LAYER M1 ;
      RECT 83295 335 83545 3865 ;
    LAYER M1 ;
      RECT 83725 335 83975 3865 ;
    LAYER M1 ;
      RECT 83725 4115 83975 5125 ;
    LAYER M1 ;
      RECT 83725 6215 83975 7225 ;
    LAYER M1 ;
      RECT 84155 335 84405 3865 ;
    LAYER M1 ;
      RECT 84585 335 84835 3865 ;
    LAYER M1 ;
      RECT 84585 4115 84835 5125 ;
    LAYER M1 ;
      RECT 84585 6215 84835 7225 ;
    LAYER M1 ;
      RECT 85015 335 85265 3865 ;
    LAYER M1 ;
      RECT 85445 335 85695 3865 ;
    LAYER M1 ;
      RECT 85445 4115 85695 5125 ;
    LAYER M1 ;
      RECT 85445 6215 85695 7225 ;
    LAYER M1 ;
      RECT 85875 335 86125 3865 ;
    LAYER M1 ;
      RECT 86305 335 86555 3865 ;
    LAYER M1 ;
      RECT 86305 4115 86555 5125 ;
    LAYER M1 ;
      RECT 86305 6215 86555 7225 ;
    LAYER M1 ;
      RECT 86735 335 86985 3865 ;
    LAYER M1 ;
      RECT 87165 335 87415 3865 ;
    LAYER M1 ;
      RECT 87165 4115 87415 5125 ;
    LAYER M1 ;
      RECT 87165 6215 87415 7225 ;
    LAYER M1 ;
      RECT 87595 335 87845 3865 ;
    LAYER M1 ;
      RECT 88025 335 88275 3865 ;
    LAYER M1 ;
      RECT 88025 4115 88275 5125 ;
    LAYER M1 ;
      RECT 88025 6215 88275 7225 ;
    LAYER M1 ;
      RECT 88455 335 88705 3865 ;
    LAYER M1 ;
      RECT 88885 335 89135 3865 ;
    LAYER M1 ;
      RECT 88885 4115 89135 5125 ;
    LAYER M1 ;
      RECT 88885 6215 89135 7225 ;
    LAYER M1 ;
      RECT 89315 335 89565 3865 ;
    LAYER M1 ;
      RECT 89745 335 89995 3865 ;
    LAYER M1 ;
      RECT 89745 4115 89995 5125 ;
    LAYER M1 ;
      RECT 89745 6215 89995 7225 ;
    LAYER M1 ;
      RECT 90175 335 90425 3865 ;
    LAYER M1 ;
      RECT 90605 335 90855 3865 ;
    LAYER M1 ;
      RECT 90605 4115 90855 5125 ;
    LAYER M1 ;
      RECT 90605 6215 90855 7225 ;
    LAYER M1 ;
      RECT 91035 335 91285 3865 ;
    LAYER M1 ;
      RECT 91465 335 91715 3865 ;
    LAYER M1 ;
      RECT 91465 4115 91715 5125 ;
    LAYER M1 ;
      RECT 91465 6215 91715 7225 ;
    LAYER M1 ;
      RECT 91895 335 92145 3865 ;
    LAYER M1 ;
      RECT 92325 335 92575 3865 ;
    LAYER M1 ;
      RECT 92325 4115 92575 5125 ;
    LAYER M1 ;
      RECT 92325 6215 92575 7225 ;
    LAYER M1 ;
      RECT 92755 335 93005 3865 ;
    LAYER M1 ;
      RECT 93185 335 93435 3865 ;
    LAYER M1 ;
      RECT 93185 4115 93435 5125 ;
    LAYER M1 ;
      RECT 93185 6215 93435 7225 ;
    LAYER M1 ;
      RECT 93615 335 93865 3865 ;
    LAYER M1 ;
      RECT 94045 335 94295 3865 ;
    LAYER M1 ;
      RECT 94045 4115 94295 5125 ;
    LAYER M1 ;
      RECT 94045 6215 94295 7225 ;
    LAYER M1 ;
      RECT 94475 335 94725 3865 ;
    LAYER M1 ;
      RECT 94905 335 95155 3865 ;
    LAYER M1 ;
      RECT 94905 4115 95155 5125 ;
    LAYER M1 ;
      RECT 94905 6215 95155 7225 ;
    LAYER M1 ;
      RECT 95335 335 95585 3865 ;
    LAYER M1 ;
      RECT 95765 335 96015 3865 ;
    LAYER M1 ;
      RECT 95765 4115 96015 5125 ;
    LAYER M1 ;
      RECT 95765 6215 96015 7225 ;
    LAYER M1 ;
      RECT 96195 335 96445 3865 ;
    LAYER M1 ;
      RECT 96625 335 96875 3865 ;
    LAYER M1 ;
      RECT 96625 4115 96875 5125 ;
    LAYER M1 ;
      RECT 96625 6215 96875 7225 ;
    LAYER M1 ;
      RECT 97055 335 97305 3865 ;
    LAYER M1 ;
      RECT 97485 335 97735 3865 ;
    LAYER M1 ;
      RECT 97485 4115 97735 5125 ;
    LAYER M1 ;
      RECT 97485 6215 97735 7225 ;
    LAYER M1 ;
      RECT 97915 335 98165 3865 ;
    LAYER M1 ;
      RECT 98345 335 98595 3865 ;
    LAYER M1 ;
      RECT 98345 4115 98595 5125 ;
    LAYER M1 ;
      RECT 98345 6215 98595 7225 ;
    LAYER M1 ;
      RECT 98775 335 99025 3865 ;
    LAYER M1 ;
      RECT 99205 335 99455 3865 ;
    LAYER M1 ;
      RECT 99205 4115 99455 5125 ;
    LAYER M1 ;
      RECT 99205 6215 99455 7225 ;
    LAYER M1 ;
      RECT 99635 335 99885 3865 ;
    LAYER M1 ;
      RECT 100065 335 100315 3865 ;
    LAYER M1 ;
      RECT 100065 4115 100315 5125 ;
    LAYER M1 ;
      RECT 100065 6215 100315 7225 ;
    LAYER M1 ;
      RECT 100495 335 100745 3865 ;
    LAYER M1 ;
      RECT 100925 335 101175 3865 ;
    LAYER M1 ;
      RECT 100925 4115 101175 5125 ;
    LAYER M1 ;
      RECT 100925 6215 101175 7225 ;
    LAYER M1 ;
      RECT 101355 335 101605 3865 ;
    LAYER M1 ;
      RECT 101785 335 102035 3865 ;
    LAYER M1 ;
      RECT 101785 4115 102035 5125 ;
    LAYER M1 ;
      RECT 101785 6215 102035 7225 ;
    LAYER M1 ;
      RECT 102215 335 102465 3865 ;
    LAYER M1 ;
      RECT 102645 335 102895 3865 ;
    LAYER M1 ;
      RECT 102645 4115 102895 5125 ;
    LAYER M1 ;
      RECT 102645 6215 102895 7225 ;
    LAYER M1 ;
      RECT 103075 335 103325 3865 ;
    LAYER M1 ;
      RECT 103505 335 103755 3865 ;
    LAYER M1 ;
      RECT 103505 4115 103755 5125 ;
    LAYER M1 ;
      RECT 103505 6215 103755 7225 ;
    LAYER M1 ;
      RECT 103935 335 104185 3865 ;
    LAYER M1 ;
      RECT 104365 335 104615 3865 ;
    LAYER M1 ;
      RECT 104365 4115 104615 5125 ;
    LAYER M1 ;
      RECT 104365 6215 104615 7225 ;
    LAYER M1 ;
      RECT 104795 335 105045 3865 ;
    LAYER M1 ;
      RECT 105225 335 105475 3865 ;
    LAYER M1 ;
      RECT 105225 4115 105475 5125 ;
    LAYER M1 ;
      RECT 105225 6215 105475 7225 ;
    LAYER M1 ;
      RECT 105655 335 105905 3865 ;
    LAYER M1 ;
      RECT 106085 335 106335 3865 ;
    LAYER M1 ;
      RECT 106085 4115 106335 5125 ;
    LAYER M1 ;
      RECT 106085 6215 106335 7225 ;
    LAYER M1 ;
      RECT 106515 335 106765 3865 ;
    LAYER M1 ;
      RECT 106945 335 107195 3865 ;
    LAYER M1 ;
      RECT 106945 4115 107195 5125 ;
    LAYER M1 ;
      RECT 106945 6215 107195 7225 ;
    LAYER M1 ;
      RECT 107375 335 107625 3865 ;
    LAYER M1 ;
      RECT 107805 335 108055 3865 ;
    LAYER M1 ;
      RECT 107805 4115 108055 5125 ;
    LAYER M1 ;
      RECT 107805 6215 108055 7225 ;
    LAYER M1 ;
      RECT 108235 335 108485 3865 ;
    LAYER M1 ;
      RECT 108665 335 108915 3865 ;
    LAYER M1 ;
      RECT 108665 4115 108915 5125 ;
    LAYER M1 ;
      RECT 108665 6215 108915 7225 ;
    LAYER M1 ;
      RECT 109095 335 109345 3865 ;
    LAYER M1 ;
      RECT 109525 335 109775 3865 ;
    LAYER M1 ;
      RECT 109525 4115 109775 5125 ;
    LAYER M1 ;
      RECT 109525 6215 109775 7225 ;
    LAYER M1 ;
      RECT 109955 335 110205 3865 ;
    LAYER M1 ;
      RECT 110385 335 110635 3865 ;
    LAYER M1 ;
      RECT 110385 4115 110635 5125 ;
    LAYER M1 ;
      RECT 110385 6215 110635 7225 ;
    LAYER M1 ;
      RECT 110815 335 111065 3865 ;
    LAYER M1 ;
      RECT 111245 335 111495 3865 ;
    LAYER M1 ;
      RECT 111245 4115 111495 5125 ;
    LAYER M1 ;
      RECT 111245 6215 111495 7225 ;
    LAYER M1 ;
      RECT 111675 335 111925 3865 ;
    LAYER M1 ;
      RECT 112105 335 112355 3865 ;
    LAYER M1 ;
      RECT 112105 4115 112355 5125 ;
    LAYER M1 ;
      RECT 112105 6215 112355 7225 ;
    LAYER M1 ;
      RECT 112535 335 112785 3865 ;
    LAYER M1 ;
      RECT 112965 335 113215 3865 ;
    LAYER M1 ;
      RECT 112965 4115 113215 5125 ;
    LAYER M1 ;
      RECT 112965 6215 113215 7225 ;
    LAYER M1 ;
      RECT 113395 335 113645 3865 ;
    LAYER M1 ;
      RECT 113825 335 114075 3865 ;
    LAYER M1 ;
      RECT 113825 4115 114075 5125 ;
    LAYER M1 ;
      RECT 113825 6215 114075 7225 ;
    LAYER M1 ;
      RECT 114255 335 114505 3865 ;
    LAYER M1 ;
      RECT 114685 335 114935 3865 ;
    LAYER M1 ;
      RECT 114685 4115 114935 5125 ;
    LAYER M1 ;
      RECT 114685 6215 114935 7225 ;
    LAYER M1 ;
      RECT 115115 335 115365 3865 ;
    LAYER M1 ;
      RECT 115545 335 115795 3865 ;
    LAYER M1 ;
      RECT 115545 4115 115795 5125 ;
    LAYER M1 ;
      RECT 115545 6215 115795 7225 ;
    LAYER M1 ;
      RECT 115975 335 116225 3865 ;
    LAYER M1 ;
      RECT 116405 335 116655 3865 ;
    LAYER M1 ;
      RECT 116405 4115 116655 5125 ;
    LAYER M1 ;
      RECT 116405 6215 116655 7225 ;
    LAYER M1 ;
      RECT 116835 335 117085 3865 ;
    LAYER M1 ;
      RECT 117265 335 117515 3865 ;
    LAYER M1 ;
      RECT 117265 4115 117515 5125 ;
    LAYER M1 ;
      RECT 117265 6215 117515 7225 ;
    LAYER M1 ;
      RECT 117695 335 117945 3865 ;
    LAYER M1 ;
      RECT 118125 335 118375 3865 ;
    LAYER M1 ;
      RECT 118125 4115 118375 5125 ;
    LAYER M1 ;
      RECT 118125 6215 118375 7225 ;
    LAYER M1 ;
      RECT 118555 335 118805 3865 ;
    LAYER M1 ;
      RECT 118985 335 119235 3865 ;
    LAYER M1 ;
      RECT 118985 4115 119235 5125 ;
    LAYER M1 ;
      RECT 118985 6215 119235 7225 ;
    LAYER M1 ;
      RECT 119415 335 119665 3865 ;
    LAYER M1 ;
      RECT 119845 335 120095 3865 ;
    LAYER M1 ;
      RECT 119845 4115 120095 5125 ;
    LAYER M1 ;
      RECT 119845 6215 120095 7225 ;
    LAYER M1 ;
      RECT 120275 335 120525 3865 ;
    LAYER M1 ;
      RECT 120705 335 120955 3865 ;
    LAYER M1 ;
      RECT 120705 4115 120955 5125 ;
    LAYER M1 ;
      RECT 120705 6215 120955 7225 ;
    LAYER M1 ;
      RECT 121135 335 121385 3865 ;
    LAYER M1 ;
      RECT 121565 335 121815 3865 ;
    LAYER M1 ;
      RECT 121565 4115 121815 5125 ;
    LAYER M1 ;
      RECT 121565 6215 121815 7225 ;
    LAYER M1 ;
      RECT 121995 335 122245 3865 ;
    LAYER M1 ;
      RECT 122425 335 122675 3865 ;
    LAYER M1 ;
      RECT 122425 4115 122675 5125 ;
    LAYER M1 ;
      RECT 122425 6215 122675 7225 ;
    LAYER M1 ;
      RECT 122855 335 123105 3865 ;
    LAYER M1 ;
      RECT 123285 335 123535 3865 ;
    LAYER M1 ;
      RECT 123285 4115 123535 5125 ;
    LAYER M1 ;
      RECT 123285 6215 123535 7225 ;
    LAYER M1 ;
      RECT 123715 335 123965 3865 ;
    LAYER M1 ;
      RECT 124145 335 124395 3865 ;
    LAYER M1 ;
      RECT 124145 4115 124395 5125 ;
    LAYER M1 ;
      RECT 124145 6215 124395 7225 ;
    LAYER M1 ;
      RECT 124575 335 124825 3865 ;
    LAYER M1 ;
      RECT 125005 335 125255 3865 ;
    LAYER M1 ;
      RECT 125005 4115 125255 5125 ;
    LAYER M1 ;
      RECT 125005 6215 125255 7225 ;
    LAYER M1 ;
      RECT 125435 335 125685 3865 ;
    LAYER M1 ;
      RECT 125865 335 126115 3865 ;
    LAYER M1 ;
      RECT 125865 4115 126115 5125 ;
    LAYER M1 ;
      RECT 125865 6215 126115 7225 ;
    LAYER M1 ;
      RECT 126295 335 126545 3865 ;
    LAYER M1 ;
      RECT 126725 335 126975 3865 ;
    LAYER M1 ;
      RECT 126725 4115 126975 5125 ;
    LAYER M1 ;
      RECT 126725 6215 126975 7225 ;
    LAYER M1 ;
      RECT 127155 335 127405 3865 ;
    LAYER M1 ;
      RECT 127585 335 127835 3865 ;
    LAYER M1 ;
      RECT 127585 4115 127835 5125 ;
    LAYER M1 ;
      RECT 127585 6215 127835 7225 ;
    LAYER M1 ;
      RECT 128015 335 128265 3865 ;
    LAYER M2 ;
      RECT 1120 4480 127880 4760 ;
    LAYER M2 ;
      RECT 1120 280 127880 560 ;
    LAYER M2 ;
      RECT 1120 6580 127880 6860 ;
    LAYER M2 ;
      RECT 690 700 128310 980 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6635 3955 6805 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6635 5675 6805 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6635 6535 6805 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6635 7395 6805 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6635 8255 6805 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6635 9115 6805 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6635 9975 6805 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6635 10835 6805 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6635 11695 6805 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6635 12555 6805 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6635 13415 6805 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6635 14275 6805 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6635 15135 6805 ;
    LAYER V1 ;
      RECT 15825 335 15995 505 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6635 15995 6805 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6635 16855 6805 ;
    LAYER V1 ;
      RECT 17545 335 17715 505 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6635 17715 6805 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6635 18575 6805 ;
    LAYER V1 ;
      RECT 19265 335 19435 505 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6635 19435 6805 ;
    LAYER V1 ;
      RECT 20125 335 20295 505 ;
    LAYER V1 ;
      RECT 20125 4535 20295 4705 ;
    LAYER V1 ;
      RECT 20125 6635 20295 6805 ;
    LAYER V1 ;
      RECT 20985 335 21155 505 ;
    LAYER V1 ;
      RECT 20985 4535 21155 4705 ;
    LAYER V1 ;
      RECT 20985 6635 21155 6805 ;
    LAYER V1 ;
      RECT 21845 335 22015 505 ;
    LAYER V1 ;
      RECT 21845 4535 22015 4705 ;
    LAYER V1 ;
      RECT 21845 6635 22015 6805 ;
    LAYER V1 ;
      RECT 22705 335 22875 505 ;
    LAYER V1 ;
      RECT 22705 4535 22875 4705 ;
    LAYER V1 ;
      RECT 22705 6635 22875 6805 ;
    LAYER V1 ;
      RECT 23565 335 23735 505 ;
    LAYER V1 ;
      RECT 23565 4535 23735 4705 ;
    LAYER V1 ;
      RECT 23565 6635 23735 6805 ;
    LAYER V1 ;
      RECT 24425 335 24595 505 ;
    LAYER V1 ;
      RECT 24425 4535 24595 4705 ;
    LAYER V1 ;
      RECT 24425 6635 24595 6805 ;
    LAYER V1 ;
      RECT 25285 335 25455 505 ;
    LAYER V1 ;
      RECT 25285 4535 25455 4705 ;
    LAYER V1 ;
      RECT 25285 6635 25455 6805 ;
    LAYER V1 ;
      RECT 26145 335 26315 505 ;
    LAYER V1 ;
      RECT 26145 4535 26315 4705 ;
    LAYER V1 ;
      RECT 26145 6635 26315 6805 ;
    LAYER V1 ;
      RECT 27005 335 27175 505 ;
    LAYER V1 ;
      RECT 27005 4535 27175 4705 ;
    LAYER V1 ;
      RECT 27005 6635 27175 6805 ;
    LAYER V1 ;
      RECT 27865 335 28035 505 ;
    LAYER V1 ;
      RECT 27865 4535 28035 4705 ;
    LAYER V1 ;
      RECT 27865 6635 28035 6805 ;
    LAYER V1 ;
      RECT 28725 335 28895 505 ;
    LAYER V1 ;
      RECT 28725 4535 28895 4705 ;
    LAYER V1 ;
      RECT 28725 6635 28895 6805 ;
    LAYER V1 ;
      RECT 29585 335 29755 505 ;
    LAYER V1 ;
      RECT 29585 4535 29755 4705 ;
    LAYER V1 ;
      RECT 29585 6635 29755 6805 ;
    LAYER V1 ;
      RECT 30445 335 30615 505 ;
    LAYER V1 ;
      RECT 30445 4535 30615 4705 ;
    LAYER V1 ;
      RECT 30445 6635 30615 6805 ;
    LAYER V1 ;
      RECT 31305 335 31475 505 ;
    LAYER V1 ;
      RECT 31305 4535 31475 4705 ;
    LAYER V1 ;
      RECT 31305 6635 31475 6805 ;
    LAYER V1 ;
      RECT 32165 335 32335 505 ;
    LAYER V1 ;
      RECT 32165 4535 32335 4705 ;
    LAYER V1 ;
      RECT 32165 6635 32335 6805 ;
    LAYER V1 ;
      RECT 33025 335 33195 505 ;
    LAYER V1 ;
      RECT 33025 4535 33195 4705 ;
    LAYER V1 ;
      RECT 33025 6635 33195 6805 ;
    LAYER V1 ;
      RECT 33885 335 34055 505 ;
    LAYER V1 ;
      RECT 33885 4535 34055 4705 ;
    LAYER V1 ;
      RECT 33885 6635 34055 6805 ;
    LAYER V1 ;
      RECT 34745 335 34915 505 ;
    LAYER V1 ;
      RECT 34745 4535 34915 4705 ;
    LAYER V1 ;
      RECT 34745 6635 34915 6805 ;
    LAYER V1 ;
      RECT 35605 335 35775 505 ;
    LAYER V1 ;
      RECT 35605 4535 35775 4705 ;
    LAYER V1 ;
      RECT 35605 6635 35775 6805 ;
    LAYER V1 ;
      RECT 36465 335 36635 505 ;
    LAYER V1 ;
      RECT 36465 4535 36635 4705 ;
    LAYER V1 ;
      RECT 36465 6635 36635 6805 ;
    LAYER V1 ;
      RECT 37325 335 37495 505 ;
    LAYER V1 ;
      RECT 37325 4535 37495 4705 ;
    LAYER V1 ;
      RECT 37325 6635 37495 6805 ;
    LAYER V1 ;
      RECT 38185 335 38355 505 ;
    LAYER V1 ;
      RECT 38185 4535 38355 4705 ;
    LAYER V1 ;
      RECT 38185 6635 38355 6805 ;
    LAYER V1 ;
      RECT 39045 335 39215 505 ;
    LAYER V1 ;
      RECT 39045 4535 39215 4705 ;
    LAYER V1 ;
      RECT 39045 6635 39215 6805 ;
    LAYER V1 ;
      RECT 39905 335 40075 505 ;
    LAYER V1 ;
      RECT 39905 4535 40075 4705 ;
    LAYER V1 ;
      RECT 39905 6635 40075 6805 ;
    LAYER V1 ;
      RECT 40765 335 40935 505 ;
    LAYER V1 ;
      RECT 40765 4535 40935 4705 ;
    LAYER V1 ;
      RECT 40765 6635 40935 6805 ;
    LAYER V1 ;
      RECT 41625 335 41795 505 ;
    LAYER V1 ;
      RECT 41625 4535 41795 4705 ;
    LAYER V1 ;
      RECT 41625 6635 41795 6805 ;
    LAYER V1 ;
      RECT 42485 335 42655 505 ;
    LAYER V1 ;
      RECT 42485 4535 42655 4705 ;
    LAYER V1 ;
      RECT 42485 6635 42655 6805 ;
    LAYER V1 ;
      RECT 43345 335 43515 505 ;
    LAYER V1 ;
      RECT 43345 4535 43515 4705 ;
    LAYER V1 ;
      RECT 43345 6635 43515 6805 ;
    LAYER V1 ;
      RECT 44205 335 44375 505 ;
    LAYER V1 ;
      RECT 44205 4535 44375 4705 ;
    LAYER V1 ;
      RECT 44205 6635 44375 6805 ;
    LAYER V1 ;
      RECT 45065 335 45235 505 ;
    LAYER V1 ;
      RECT 45065 4535 45235 4705 ;
    LAYER V1 ;
      RECT 45065 6635 45235 6805 ;
    LAYER V1 ;
      RECT 45925 335 46095 505 ;
    LAYER V1 ;
      RECT 45925 4535 46095 4705 ;
    LAYER V1 ;
      RECT 45925 6635 46095 6805 ;
    LAYER V1 ;
      RECT 46785 335 46955 505 ;
    LAYER V1 ;
      RECT 46785 4535 46955 4705 ;
    LAYER V1 ;
      RECT 46785 6635 46955 6805 ;
    LAYER V1 ;
      RECT 47645 335 47815 505 ;
    LAYER V1 ;
      RECT 47645 4535 47815 4705 ;
    LAYER V1 ;
      RECT 47645 6635 47815 6805 ;
    LAYER V1 ;
      RECT 48505 335 48675 505 ;
    LAYER V1 ;
      RECT 48505 4535 48675 4705 ;
    LAYER V1 ;
      RECT 48505 6635 48675 6805 ;
    LAYER V1 ;
      RECT 49365 335 49535 505 ;
    LAYER V1 ;
      RECT 49365 4535 49535 4705 ;
    LAYER V1 ;
      RECT 49365 6635 49535 6805 ;
    LAYER V1 ;
      RECT 50225 335 50395 505 ;
    LAYER V1 ;
      RECT 50225 4535 50395 4705 ;
    LAYER V1 ;
      RECT 50225 6635 50395 6805 ;
    LAYER V1 ;
      RECT 51085 335 51255 505 ;
    LAYER V1 ;
      RECT 51085 4535 51255 4705 ;
    LAYER V1 ;
      RECT 51085 6635 51255 6805 ;
    LAYER V1 ;
      RECT 51945 335 52115 505 ;
    LAYER V1 ;
      RECT 51945 4535 52115 4705 ;
    LAYER V1 ;
      RECT 51945 6635 52115 6805 ;
    LAYER V1 ;
      RECT 52805 335 52975 505 ;
    LAYER V1 ;
      RECT 52805 4535 52975 4705 ;
    LAYER V1 ;
      RECT 52805 6635 52975 6805 ;
    LAYER V1 ;
      RECT 53665 335 53835 505 ;
    LAYER V1 ;
      RECT 53665 4535 53835 4705 ;
    LAYER V1 ;
      RECT 53665 6635 53835 6805 ;
    LAYER V1 ;
      RECT 54525 335 54695 505 ;
    LAYER V1 ;
      RECT 54525 4535 54695 4705 ;
    LAYER V1 ;
      RECT 54525 6635 54695 6805 ;
    LAYER V1 ;
      RECT 55385 335 55555 505 ;
    LAYER V1 ;
      RECT 55385 4535 55555 4705 ;
    LAYER V1 ;
      RECT 55385 6635 55555 6805 ;
    LAYER V1 ;
      RECT 56245 335 56415 505 ;
    LAYER V1 ;
      RECT 56245 4535 56415 4705 ;
    LAYER V1 ;
      RECT 56245 6635 56415 6805 ;
    LAYER V1 ;
      RECT 57105 335 57275 505 ;
    LAYER V1 ;
      RECT 57105 4535 57275 4705 ;
    LAYER V1 ;
      RECT 57105 6635 57275 6805 ;
    LAYER V1 ;
      RECT 57965 335 58135 505 ;
    LAYER V1 ;
      RECT 57965 4535 58135 4705 ;
    LAYER V1 ;
      RECT 57965 6635 58135 6805 ;
    LAYER V1 ;
      RECT 58825 335 58995 505 ;
    LAYER V1 ;
      RECT 58825 4535 58995 4705 ;
    LAYER V1 ;
      RECT 58825 6635 58995 6805 ;
    LAYER V1 ;
      RECT 59685 335 59855 505 ;
    LAYER V1 ;
      RECT 59685 4535 59855 4705 ;
    LAYER V1 ;
      RECT 59685 6635 59855 6805 ;
    LAYER V1 ;
      RECT 60545 335 60715 505 ;
    LAYER V1 ;
      RECT 60545 4535 60715 4705 ;
    LAYER V1 ;
      RECT 60545 6635 60715 6805 ;
    LAYER V1 ;
      RECT 61405 335 61575 505 ;
    LAYER V1 ;
      RECT 61405 4535 61575 4705 ;
    LAYER V1 ;
      RECT 61405 6635 61575 6805 ;
    LAYER V1 ;
      RECT 62265 335 62435 505 ;
    LAYER V1 ;
      RECT 62265 4535 62435 4705 ;
    LAYER V1 ;
      RECT 62265 6635 62435 6805 ;
    LAYER V1 ;
      RECT 63125 335 63295 505 ;
    LAYER V1 ;
      RECT 63125 4535 63295 4705 ;
    LAYER V1 ;
      RECT 63125 6635 63295 6805 ;
    LAYER V1 ;
      RECT 63985 335 64155 505 ;
    LAYER V1 ;
      RECT 63985 4535 64155 4705 ;
    LAYER V1 ;
      RECT 63985 6635 64155 6805 ;
    LAYER V1 ;
      RECT 64845 335 65015 505 ;
    LAYER V1 ;
      RECT 64845 4535 65015 4705 ;
    LAYER V1 ;
      RECT 64845 6635 65015 6805 ;
    LAYER V1 ;
      RECT 65705 335 65875 505 ;
    LAYER V1 ;
      RECT 65705 4535 65875 4705 ;
    LAYER V1 ;
      RECT 65705 6635 65875 6805 ;
    LAYER V1 ;
      RECT 66565 335 66735 505 ;
    LAYER V1 ;
      RECT 66565 4535 66735 4705 ;
    LAYER V1 ;
      RECT 66565 6635 66735 6805 ;
    LAYER V1 ;
      RECT 67425 335 67595 505 ;
    LAYER V1 ;
      RECT 67425 4535 67595 4705 ;
    LAYER V1 ;
      RECT 67425 6635 67595 6805 ;
    LAYER V1 ;
      RECT 68285 335 68455 505 ;
    LAYER V1 ;
      RECT 68285 4535 68455 4705 ;
    LAYER V1 ;
      RECT 68285 6635 68455 6805 ;
    LAYER V1 ;
      RECT 69145 335 69315 505 ;
    LAYER V1 ;
      RECT 69145 4535 69315 4705 ;
    LAYER V1 ;
      RECT 69145 6635 69315 6805 ;
    LAYER V1 ;
      RECT 70005 335 70175 505 ;
    LAYER V1 ;
      RECT 70005 4535 70175 4705 ;
    LAYER V1 ;
      RECT 70005 6635 70175 6805 ;
    LAYER V1 ;
      RECT 70865 335 71035 505 ;
    LAYER V1 ;
      RECT 70865 4535 71035 4705 ;
    LAYER V1 ;
      RECT 70865 6635 71035 6805 ;
    LAYER V1 ;
      RECT 71725 335 71895 505 ;
    LAYER V1 ;
      RECT 71725 4535 71895 4705 ;
    LAYER V1 ;
      RECT 71725 6635 71895 6805 ;
    LAYER V1 ;
      RECT 72585 335 72755 505 ;
    LAYER V1 ;
      RECT 72585 4535 72755 4705 ;
    LAYER V1 ;
      RECT 72585 6635 72755 6805 ;
    LAYER V1 ;
      RECT 73445 335 73615 505 ;
    LAYER V1 ;
      RECT 73445 4535 73615 4705 ;
    LAYER V1 ;
      RECT 73445 6635 73615 6805 ;
    LAYER V1 ;
      RECT 74305 335 74475 505 ;
    LAYER V1 ;
      RECT 74305 4535 74475 4705 ;
    LAYER V1 ;
      RECT 74305 6635 74475 6805 ;
    LAYER V1 ;
      RECT 75165 335 75335 505 ;
    LAYER V1 ;
      RECT 75165 4535 75335 4705 ;
    LAYER V1 ;
      RECT 75165 6635 75335 6805 ;
    LAYER V1 ;
      RECT 76025 335 76195 505 ;
    LAYER V1 ;
      RECT 76025 4535 76195 4705 ;
    LAYER V1 ;
      RECT 76025 6635 76195 6805 ;
    LAYER V1 ;
      RECT 76885 335 77055 505 ;
    LAYER V1 ;
      RECT 76885 4535 77055 4705 ;
    LAYER V1 ;
      RECT 76885 6635 77055 6805 ;
    LAYER V1 ;
      RECT 77745 335 77915 505 ;
    LAYER V1 ;
      RECT 77745 4535 77915 4705 ;
    LAYER V1 ;
      RECT 77745 6635 77915 6805 ;
    LAYER V1 ;
      RECT 78605 335 78775 505 ;
    LAYER V1 ;
      RECT 78605 4535 78775 4705 ;
    LAYER V1 ;
      RECT 78605 6635 78775 6805 ;
    LAYER V1 ;
      RECT 79465 335 79635 505 ;
    LAYER V1 ;
      RECT 79465 4535 79635 4705 ;
    LAYER V1 ;
      RECT 79465 6635 79635 6805 ;
    LAYER V1 ;
      RECT 80325 335 80495 505 ;
    LAYER V1 ;
      RECT 80325 4535 80495 4705 ;
    LAYER V1 ;
      RECT 80325 6635 80495 6805 ;
    LAYER V1 ;
      RECT 81185 335 81355 505 ;
    LAYER V1 ;
      RECT 81185 4535 81355 4705 ;
    LAYER V1 ;
      RECT 81185 6635 81355 6805 ;
    LAYER V1 ;
      RECT 82045 335 82215 505 ;
    LAYER V1 ;
      RECT 82045 4535 82215 4705 ;
    LAYER V1 ;
      RECT 82045 6635 82215 6805 ;
    LAYER V1 ;
      RECT 82905 335 83075 505 ;
    LAYER V1 ;
      RECT 82905 4535 83075 4705 ;
    LAYER V1 ;
      RECT 82905 6635 83075 6805 ;
    LAYER V1 ;
      RECT 83765 335 83935 505 ;
    LAYER V1 ;
      RECT 83765 4535 83935 4705 ;
    LAYER V1 ;
      RECT 83765 6635 83935 6805 ;
    LAYER V1 ;
      RECT 84625 335 84795 505 ;
    LAYER V1 ;
      RECT 84625 4535 84795 4705 ;
    LAYER V1 ;
      RECT 84625 6635 84795 6805 ;
    LAYER V1 ;
      RECT 85485 335 85655 505 ;
    LAYER V1 ;
      RECT 85485 4535 85655 4705 ;
    LAYER V1 ;
      RECT 85485 6635 85655 6805 ;
    LAYER V1 ;
      RECT 86345 335 86515 505 ;
    LAYER V1 ;
      RECT 86345 4535 86515 4705 ;
    LAYER V1 ;
      RECT 86345 6635 86515 6805 ;
    LAYER V1 ;
      RECT 87205 335 87375 505 ;
    LAYER V1 ;
      RECT 87205 4535 87375 4705 ;
    LAYER V1 ;
      RECT 87205 6635 87375 6805 ;
    LAYER V1 ;
      RECT 88065 335 88235 505 ;
    LAYER V1 ;
      RECT 88065 4535 88235 4705 ;
    LAYER V1 ;
      RECT 88065 6635 88235 6805 ;
    LAYER V1 ;
      RECT 88925 335 89095 505 ;
    LAYER V1 ;
      RECT 88925 4535 89095 4705 ;
    LAYER V1 ;
      RECT 88925 6635 89095 6805 ;
    LAYER V1 ;
      RECT 89785 335 89955 505 ;
    LAYER V1 ;
      RECT 89785 4535 89955 4705 ;
    LAYER V1 ;
      RECT 89785 6635 89955 6805 ;
    LAYER V1 ;
      RECT 90645 335 90815 505 ;
    LAYER V1 ;
      RECT 90645 4535 90815 4705 ;
    LAYER V1 ;
      RECT 90645 6635 90815 6805 ;
    LAYER V1 ;
      RECT 91505 335 91675 505 ;
    LAYER V1 ;
      RECT 91505 4535 91675 4705 ;
    LAYER V1 ;
      RECT 91505 6635 91675 6805 ;
    LAYER V1 ;
      RECT 92365 335 92535 505 ;
    LAYER V1 ;
      RECT 92365 4535 92535 4705 ;
    LAYER V1 ;
      RECT 92365 6635 92535 6805 ;
    LAYER V1 ;
      RECT 93225 335 93395 505 ;
    LAYER V1 ;
      RECT 93225 4535 93395 4705 ;
    LAYER V1 ;
      RECT 93225 6635 93395 6805 ;
    LAYER V1 ;
      RECT 94085 335 94255 505 ;
    LAYER V1 ;
      RECT 94085 4535 94255 4705 ;
    LAYER V1 ;
      RECT 94085 6635 94255 6805 ;
    LAYER V1 ;
      RECT 94945 335 95115 505 ;
    LAYER V1 ;
      RECT 94945 4535 95115 4705 ;
    LAYER V1 ;
      RECT 94945 6635 95115 6805 ;
    LAYER V1 ;
      RECT 95805 335 95975 505 ;
    LAYER V1 ;
      RECT 95805 4535 95975 4705 ;
    LAYER V1 ;
      RECT 95805 6635 95975 6805 ;
    LAYER V1 ;
      RECT 96665 335 96835 505 ;
    LAYER V1 ;
      RECT 96665 4535 96835 4705 ;
    LAYER V1 ;
      RECT 96665 6635 96835 6805 ;
    LAYER V1 ;
      RECT 97525 335 97695 505 ;
    LAYER V1 ;
      RECT 97525 4535 97695 4705 ;
    LAYER V1 ;
      RECT 97525 6635 97695 6805 ;
    LAYER V1 ;
      RECT 98385 335 98555 505 ;
    LAYER V1 ;
      RECT 98385 4535 98555 4705 ;
    LAYER V1 ;
      RECT 98385 6635 98555 6805 ;
    LAYER V1 ;
      RECT 99245 335 99415 505 ;
    LAYER V1 ;
      RECT 99245 4535 99415 4705 ;
    LAYER V1 ;
      RECT 99245 6635 99415 6805 ;
    LAYER V1 ;
      RECT 100105 335 100275 505 ;
    LAYER V1 ;
      RECT 100105 4535 100275 4705 ;
    LAYER V1 ;
      RECT 100105 6635 100275 6805 ;
    LAYER V1 ;
      RECT 100965 335 101135 505 ;
    LAYER V1 ;
      RECT 100965 4535 101135 4705 ;
    LAYER V1 ;
      RECT 100965 6635 101135 6805 ;
    LAYER V1 ;
      RECT 101825 335 101995 505 ;
    LAYER V1 ;
      RECT 101825 4535 101995 4705 ;
    LAYER V1 ;
      RECT 101825 6635 101995 6805 ;
    LAYER V1 ;
      RECT 102685 335 102855 505 ;
    LAYER V1 ;
      RECT 102685 4535 102855 4705 ;
    LAYER V1 ;
      RECT 102685 6635 102855 6805 ;
    LAYER V1 ;
      RECT 103545 335 103715 505 ;
    LAYER V1 ;
      RECT 103545 4535 103715 4705 ;
    LAYER V1 ;
      RECT 103545 6635 103715 6805 ;
    LAYER V1 ;
      RECT 104405 335 104575 505 ;
    LAYER V1 ;
      RECT 104405 4535 104575 4705 ;
    LAYER V1 ;
      RECT 104405 6635 104575 6805 ;
    LAYER V1 ;
      RECT 105265 335 105435 505 ;
    LAYER V1 ;
      RECT 105265 4535 105435 4705 ;
    LAYER V1 ;
      RECT 105265 6635 105435 6805 ;
    LAYER V1 ;
      RECT 106125 335 106295 505 ;
    LAYER V1 ;
      RECT 106125 4535 106295 4705 ;
    LAYER V1 ;
      RECT 106125 6635 106295 6805 ;
    LAYER V1 ;
      RECT 106985 335 107155 505 ;
    LAYER V1 ;
      RECT 106985 4535 107155 4705 ;
    LAYER V1 ;
      RECT 106985 6635 107155 6805 ;
    LAYER V1 ;
      RECT 107845 335 108015 505 ;
    LAYER V1 ;
      RECT 107845 4535 108015 4705 ;
    LAYER V1 ;
      RECT 107845 6635 108015 6805 ;
    LAYER V1 ;
      RECT 108705 335 108875 505 ;
    LAYER V1 ;
      RECT 108705 4535 108875 4705 ;
    LAYER V1 ;
      RECT 108705 6635 108875 6805 ;
    LAYER V1 ;
      RECT 109565 335 109735 505 ;
    LAYER V1 ;
      RECT 109565 4535 109735 4705 ;
    LAYER V1 ;
      RECT 109565 6635 109735 6805 ;
    LAYER V1 ;
      RECT 110425 335 110595 505 ;
    LAYER V1 ;
      RECT 110425 4535 110595 4705 ;
    LAYER V1 ;
      RECT 110425 6635 110595 6805 ;
    LAYER V1 ;
      RECT 111285 335 111455 505 ;
    LAYER V1 ;
      RECT 111285 4535 111455 4705 ;
    LAYER V1 ;
      RECT 111285 6635 111455 6805 ;
    LAYER V1 ;
      RECT 112145 335 112315 505 ;
    LAYER V1 ;
      RECT 112145 4535 112315 4705 ;
    LAYER V1 ;
      RECT 112145 6635 112315 6805 ;
    LAYER V1 ;
      RECT 113005 335 113175 505 ;
    LAYER V1 ;
      RECT 113005 4535 113175 4705 ;
    LAYER V1 ;
      RECT 113005 6635 113175 6805 ;
    LAYER V1 ;
      RECT 113865 335 114035 505 ;
    LAYER V1 ;
      RECT 113865 4535 114035 4705 ;
    LAYER V1 ;
      RECT 113865 6635 114035 6805 ;
    LAYER V1 ;
      RECT 114725 335 114895 505 ;
    LAYER V1 ;
      RECT 114725 4535 114895 4705 ;
    LAYER V1 ;
      RECT 114725 6635 114895 6805 ;
    LAYER V1 ;
      RECT 115585 335 115755 505 ;
    LAYER V1 ;
      RECT 115585 4535 115755 4705 ;
    LAYER V1 ;
      RECT 115585 6635 115755 6805 ;
    LAYER V1 ;
      RECT 116445 335 116615 505 ;
    LAYER V1 ;
      RECT 116445 4535 116615 4705 ;
    LAYER V1 ;
      RECT 116445 6635 116615 6805 ;
    LAYER V1 ;
      RECT 117305 335 117475 505 ;
    LAYER V1 ;
      RECT 117305 4535 117475 4705 ;
    LAYER V1 ;
      RECT 117305 6635 117475 6805 ;
    LAYER V1 ;
      RECT 118165 335 118335 505 ;
    LAYER V1 ;
      RECT 118165 4535 118335 4705 ;
    LAYER V1 ;
      RECT 118165 6635 118335 6805 ;
    LAYER V1 ;
      RECT 119025 335 119195 505 ;
    LAYER V1 ;
      RECT 119025 4535 119195 4705 ;
    LAYER V1 ;
      RECT 119025 6635 119195 6805 ;
    LAYER V1 ;
      RECT 119885 335 120055 505 ;
    LAYER V1 ;
      RECT 119885 4535 120055 4705 ;
    LAYER V1 ;
      RECT 119885 6635 120055 6805 ;
    LAYER V1 ;
      RECT 120745 335 120915 505 ;
    LAYER V1 ;
      RECT 120745 4535 120915 4705 ;
    LAYER V1 ;
      RECT 120745 6635 120915 6805 ;
    LAYER V1 ;
      RECT 121605 335 121775 505 ;
    LAYER V1 ;
      RECT 121605 4535 121775 4705 ;
    LAYER V1 ;
      RECT 121605 6635 121775 6805 ;
    LAYER V1 ;
      RECT 122465 335 122635 505 ;
    LAYER V1 ;
      RECT 122465 4535 122635 4705 ;
    LAYER V1 ;
      RECT 122465 6635 122635 6805 ;
    LAYER V1 ;
      RECT 123325 335 123495 505 ;
    LAYER V1 ;
      RECT 123325 4535 123495 4705 ;
    LAYER V1 ;
      RECT 123325 6635 123495 6805 ;
    LAYER V1 ;
      RECT 124185 335 124355 505 ;
    LAYER V1 ;
      RECT 124185 4535 124355 4705 ;
    LAYER V1 ;
      RECT 124185 6635 124355 6805 ;
    LAYER V1 ;
      RECT 125045 335 125215 505 ;
    LAYER V1 ;
      RECT 125045 4535 125215 4705 ;
    LAYER V1 ;
      RECT 125045 6635 125215 6805 ;
    LAYER V1 ;
      RECT 125905 335 126075 505 ;
    LAYER V1 ;
      RECT 125905 4535 126075 4705 ;
    LAYER V1 ;
      RECT 125905 6635 126075 6805 ;
    LAYER V1 ;
      RECT 126765 335 126935 505 ;
    LAYER V1 ;
      RECT 126765 4535 126935 4705 ;
    LAYER V1 ;
      RECT 126765 6635 126935 6805 ;
    LAYER V1 ;
      RECT 127625 335 127795 505 ;
    LAYER V1 ;
      RECT 127625 4535 127795 4705 ;
    LAYER V1 ;
      RECT 127625 6635 127795 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 15395 755 15565 925 ;
    LAYER V1 ;
      RECT 16255 755 16425 925 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17975 755 18145 925 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 19695 755 19865 925 ;
    LAYER V1 ;
      RECT 20555 755 20725 925 ;
    LAYER V1 ;
      RECT 21415 755 21585 925 ;
    LAYER V1 ;
      RECT 22275 755 22445 925 ;
    LAYER V1 ;
      RECT 23135 755 23305 925 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 24855 755 25025 925 ;
    LAYER V1 ;
      RECT 25715 755 25885 925 ;
    LAYER V1 ;
      RECT 26575 755 26745 925 ;
    LAYER V1 ;
      RECT 27435 755 27605 925 ;
    LAYER V1 ;
      RECT 28295 755 28465 925 ;
    LAYER V1 ;
      RECT 29155 755 29325 925 ;
    LAYER V1 ;
      RECT 30015 755 30185 925 ;
    LAYER V1 ;
      RECT 30875 755 31045 925 ;
    LAYER V1 ;
      RECT 31735 755 31905 925 ;
    LAYER V1 ;
      RECT 32595 755 32765 925 ;
    LAYER V1 ;
      RECT 33455 755 33625 925 ;
    LAYER V1 ;
      RECT 34315 755 34485 925 ;
    LAYER V1 ;
      RECT 35175 755 35345 925 ;
    LAYER V1 ;
      RECT 36035 755 36205 925 ;
    LAYER V1 ;
      RECT 36895 755 37065 925 ;
    LAYER V1 ;
      RECT 37755 755 37925 925 ;
    LAYER V1 ;
      RECT 38615 755 38785 925 ;
    LAYER V1 ;
      RECT 39475 755 39645 925 ;
    LAYER V1 ;
      RECT 40335 755 40505 925 ;
    LAYER V1 ;
      RECT 41195 755 41365 925 ;
    LAYER V1 ;
      RECT 42055 755 42225 925 ;
    LAYER V1 ;
      RECT 42915 755 43085 925 ;
    LAYER V1 ;
      RECT 43775 755 43945 925 ;
    LAYER V1 ;
      RECT 44635 755 44805 925 ;
    LAYER V1 ;
      RECT 45495 755 45665 925 ;
    LAYER V1 ;
      RECT 46355 755 46525 925 ;
    LAYER V1 ;
      RECT 47215 755 47385 925 ;
    LAYER V1 ;
      RECT 48075 755 48245 925 ;
    LAYER V1 ;
      RECT 48935 755 49105 925 ;
    LAYER V1 ;
      RECT 49795 755 49965 925 ;
    LAYER V1 ;
      RECT 50655 755 50825 925 ;
    LAYER V1 ;
      RECT 51515 755 51685 925 ;
    LAYER V1 ;
      RECT 52375 755 52545 925 ;
    LAYER V1 ;
      RECT 53235 755 53405 925 ;
    LAYER V1 ;
      RECT 54095 755 54265 925 ;
    LAYER V1 ;
      RECT 54955 755 55125 925 ;
    LAYER V1 ;
      RECT 55815 755 55985 925 ;
    LAYER V1 ;
      RECT 56675 755 56845 925 ;
    LAYER V1 ;
      RECT 57535 755 57705 925 ;
    LAYER V1 ;
      RECT 58395 755 58565 925 ;
    LAYER V1 ;
      RECT 59255 755 59425 925 ;
    LAYER V1 ;
      RECT 60115 755 60285 925 ;
    LAYER V1 ;
      RECT 60975 755 61145 925 ;
    LAYER V1 ;
      RECT 61835 755 62005 925 ;
    LAYER V1 ;
      RECT 62695 755 62865 925 ;
    LAYER V1 ;
      RECT 63555 755 63725 925 ;
    LAYER V1 ;
      RECT 64415 755 64585 925 ;
    LAYER V1 ;
      RECT 65275 755 65445 925 ;
    LAYER V1 ;
      RECT 66135 755 66305 925 ;
    LAYER V1 ;
      RECT 66995 755 67165 925 ;
    LAYER V1 ;
      RECT 67855 755 68025 925 ;
    LAYER V1 ;
      RECT 68715 755 68885 925 ;
    LAYER V1 ;
      RECT 69575 755 69745 925 ;
    LAYER V1 ;
      RECT 70435 755 70605 925 ;
    LAYER V1 ;
      RECT 71295 755 71465 925 ;
    LAYER V1 ;
      RECT 72155 755 72325 925 ;
    LAYER V1 ;
      RECT 73015 755 73185 925 ;
    LAYER V1 ;
      RECT 73875 755 74045 925 ;
    LAYER V1 ;
      RECT 74735 755 74905 925 ;
    LAYER V1 ;
      RECT 75595 755 75765 925 ;
    LAYER V1 ;
      RECT 76455 755 76625 925 ;
    LAYER V1 ;
      RECT 77315 755 77485 925 ;
    LAYER V1 ;
      RECT 78175 755 78345 925 ;
    LAYER V1 ;
      RECT 79035 755 79205 925 ;
    LAYER V1 ;
      RECT 79895 755 80065 925 ;
    LAYER V1 ;
      RECT 80755 755 80925 925 ;
    LAYER V1 ;
      RECT 81615 755 81785 925 ;
    LAYER V1 ;
      RECT 82475 755 82645 925 ;
    LAYER V1 ;
      RECT 83335 755 83505 925 ;
    LAYER V1 ;
      RECT 84195 755 84365 925 ;
    LAYER V1 ;
      RECT 85055 755 85225 925 ;
    LAYER V1 ;
      RECT 85915 755 86085 925 ;
    LAYER V1 ;
      RECT 86775 755 86945 925 ;
    LAYER V1 ;
      RECT 87635 755 87805 925 ;
    LAYER V1 ;
      RECT 88495 755 88665 925 ;
    LAYER V1 ;
      RECT 89355 755 89525 925 ;
    LAYER V1 ;
      RECT 90215 755 90385 925 ;
    LAYER V1 ;
      RECT 91075 755 91245 925 ;
    LAYER V1 ;
      RECT 91935 755 92105 925 ;
    LAYER V1 ;
      RECT 92795 755 92965 925 ;
    LAYER V1 ;
      RECT 93655 755 93825 925 ;
    LAYER V1 ;
      RECT 94515 755 94685 925 ;
    LAYER V1 ;
      RECT 95375 755 95545 925 ;
    LAYER V1 ;
      RECT 96235 755 96405 925 ;
    LAYER V1 ;
      RECT 97095 755 97265 925 ;
    LAYER V1 ;
      RECT 97955 755 98125 925 ;
    LAYER V1 ;
      RECT 98815 755 98985 925 ;
    LAYER V1 ;
      RECT 99675 755 99845 925 ;
    LAYER V1 ;
      RECT 100535 755 100705 925 ;
    LAYER V1 ;
      RECT 101395 755 101565 925 ;
    LAYER V1 ;
      RECT 102255 755 102425 925 ;
    LAYER V1 ;
      RECT 103115 755 103285 925 ;
    LAYER V1 ;
      RECT 103975 755 104145 925 ;
    LAYER V1 ;
      RECT 104835 755 105005 925 ;
    LAYER V1 ;
      RECT 105695 755 105865 925 ;
    LAYER V1 ;
      RECT 106555 755 106725 925 ;
    LAYER V1 ;
      RECT 107415 755 107585 925 ;
    LAYER V1 ;
      RECT 108275 755 108445 925 ;
    LAYER V1 ;
      RECT 109135 755 109305 925 ;
    LAYER V1 ;
      RECT 109995 755 110165 925 ;
    LAYER V1 ;
      RECT 110855 755 111025 925 ;
    LAYER V1 ;
      RECT 111715 755 111885 925 ;
    LAYER V1 ;
      RECT 112575 755 112745 925 ;
    LAYER V1 ;
      RECT 113435 755 113605 925 ;
    LAYER V1 ;
      RECT 114295 755 114465 925 ;
    LAYER V1 ;
      RECT 115155 755 115325 925 ;
    LAYER V1 ;
      RECT 116015 755 116185 925 ;
    LAYER V1 ;
      RECT 116875 755 117045 925 ;
    LAYER V1 ;
      RECT 117735 755 117905 925 ;
    LAYER V1 ;
      RECT 118595 755 118765 925 ;
    LAYER V1 ;
      RECT 119455 755 119625 925 ;
    LAYER V1 ;
      RECT 120315 755 120485 925 ;
    LAYER V1 ;
      RECT 121175 755 121345 925 ;
    LAYER V1 ;
      RECT 122035 755 122205 925 ;
    LAYER V1 ;
      RECT 122895 755 123065 925 ;
    LAYER V1 ;
      RECT 123755 755 123925 925 ;
    LAYER V1 ;
      RECT 124615 755 124785 925 ;
    LAYER V1 ;
      RECT 125475 755 125645 925 ;
    LAYER V1 ;
      RECT 126335 755 126505 925 ;
    LAYER V1 ;
      RECT 127195 755 127365 925 ;
    LAYER V1 ;
      RECT 128055 755 128225 925 ;
    LAYER V2 ;
      RECT 64425 345 64575 495 ;
    LAYER V2 ;
      RECT 64425 4545 64575 4695 ;
    LAYER V2 ;
      RECT 64855 765 65005 915 ;
    LAYER V2 ;
      RECT 64855 6645 65005 6795 ;
  END
END DCL_NMOS_S_55663590_X148_Y1
