MACRO SCM_NMOS_B_8106910_X9_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_8106910_X9_Y2 0 0 ;
  SIZE 17200 BY 13440 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 12460 16080 12740 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8030 260 8310 10660 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8460 680 8740 6880 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8890 1100 9170 7300 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 13105 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 13105 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 13105 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 13105 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 13105 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 13105 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 13105 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 13105 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 13105 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 13105 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 9745 ;
    LAYER M1 ;
      RECT 9765 9995 10015 11005 ;
    LAYER M1 ;
      RECT 9765 12095 10015 13105 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 6215 10445 9745 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 9745 ;
    LAYER M1 ;
      RECT 10625 9995 10875 11005 ;
    LAYER M1 ;
      RECT 10625 12095 10875 13105 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11055 6215 11305 9745 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 9745 ;
    LAYER M1 ;
      RECT 11485 9995 11735 11005 ;
    LAYER M1 ;
      RECT 11485 12095 11735 13105 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 11915 6215 12165 9745 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 9745 ;
    LAYER M1 ;
      RECT 12345 9995 12595 11005 ;
    LAYER M1 ;
      RECT 12345 12095 12595 13105 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 12775 6215 13025 9745 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 9745 ;
    LAYER M1 ;
      RECT 13205 9995 13455 11005 ;
    LAYER M1 ;
      RECT 13205 12095 13455 13105 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 13635 6215 13885 9745 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 9745 ;
    LAYER M1 ;
      RECT 14065 9995 14315 11005 ;
    LAYER M1 ;
      RECT 14065 12095 14315 13105 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14495 6215 14745 9745 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 9745 ;
    LAYER M1 ;
      RECT 14925 9995 15175 11005 ;
    LAYER M1 ;
      RECT 14925 12095 15175 13105 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15355 6215 15605 9745 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 9745 ;
    LAYER M1 ;
      RECT 15785 9995 16035 11005 ;
    LAYER M1 ;
      RECT 15785 12095 16035 13105 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16215 6215 16465 9745 ;
    LAYER M2 ;
      RECT 1120 4480 16080 4760 ;
    LAYER M2 ;
      RECT 1120 280 15220 560 ;
    LAYER M2 ;
      RECT 1980 700 16080 980 ;
    LAYER M2 ;
      RECT 690 1120 16510 1400 ;
    LAYER M2 ;
      RECT 1980 6160 16080 6440 ;
    LAYER M2 ;
      RECT 1120 10360 16080 10640 ;
    LAYER M2 ;
      RECT 1120 6580 15220 6860 ;
    LAYER M2 ;
      RECT 690 7000 16510 7280 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6635 13415 6805 ;
    LAYER V1 ;
      RECT 13245 10415 13415 10585 ;
    LAYER V1 ;
      RECT 13245 12515 13415 12685 ;
    LAYER V1 ;
      RECT 14105 755 14275 925 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6215 14275 6385 ;
    LAYER V1 ;
      RECT 14105 10415 14275 10585 ;
    LAYER V1 ;
      RECT 14105 12515 14275 12685 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12515 1375 12685 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6635 15135 6805 ;
    LAYER V1 ;
      RECT 14965 10415 15135 10585 ;
    LAYER V1 ;
      RECT 14965 12515 15135 12685 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12515 2235 12685 ;
    LAYER V1 ;
      RECT 15825 755 15995 925 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6215 15995 6385 ;
    LAYER V1 ;
      RECT 15825 10415 15995 10585 ;
    LAYER V1 ;
      RECT 15825 12515 15995 12685 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12515 3095 12685 ;
    LAYER V1 ;
      RECT 3785 755 3955 925 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12515 3955 12685 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12515 4815 12685 ;
    LAYER V1 ;
      RECT 5505 755 5675 925 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12515 5675 12685 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6635 6535 6805 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12515 6535 12685 ;
    LAYER V1 ;
      RECT 7225 755 7395 925 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12515 7395 12685 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6635 8255 6805 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12515 8255 12685 ;
    LAYER V1 ;
      RECT 8945 755 9115 925 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12515 9115 12685 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6635 9975 6805 ;
    LAYER V1 ;
      RECT 9805 10415 9975 10585 ;
    LAYER V1 ;
      RECT 9805 12515 9975 12685 ;
    LAYER V1 ;
      RECT 10665 755 10835 925 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6215 10835 6385 ;
    LAYER V1 ;
      RECT 10665 10415 10835 10585 ;
    LAYER V1 ;
      RECT 10665 12515 10835 12685 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6635 11695 6805 ;
    LAYER V1 ;
      RECT 11525 10415 11695 10585 ;
    LAYER V1 ;
      RECT 11525 12515 11695 12685 ;
    LAYER V1 ;
      RECT 12385 755 12555 925 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6215 12555 6385 ;
    LAYER V1 ;
      RECT 12385 10415 12555 10585 ;
    LAYER V1 ;
      RECT 12385 12515 12555 12685 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 775 7055 945 7225 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 1635 7055 1805 7225 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 2495 7055 2665 7225 ;
    LAYER V1 ;
      RECT 3355 1175 3525 1345 ;
    LAYER V1 ;
      RECT 3355 7055 3525 7225 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 4215 7055 4385 7225 ;
    LAYER V1 ;
      RECT 5075 1175 5245 1345 ;
    LAYER V1 ;
      RECT 5075 7055 5245 7225 ;
    LAYER V1 ;
      RECT 5935 1175 6105 1345 ;
    LAYER V1 ;
      RECT 5935 7055 6105 7225 ;
    LAYER V1 ;
      RECT 6795 1175 6965 1345 ;
    LAYER V1 ;
      RECT 6795 7055 6965 7225 ;
    LAYER V1 ;
      RECT 7655 1175 7825 1345 ;
    LAYER V1 ;
      RECT 7655 7055 7825 7225 ;
    LAYER V1 ;
      RECT 8515 1175 8685 1345 ;
    LAYER V1 ;
      RECT 8515 7055 8685 7225 ;
    LAYER V1 ;
      RECT 9375 1175 9545 1345 ;
    LAYER V1 ;
      RECT 9375 7055 9545 7225 ;
    LAYER V1 ;
      RECT 10235 1175 10405 1345 ;
    LAYER V1 ;
      RECT 10235 7055 10405 7225 ;
    LAYER V1 ;
      RECT 11095 1175 11265 1345 ;
    LAYER V1 ;
      RECT 11095 7055 11265 7225 ;
    LAYER V1 ;
      RECT 11955 1175 12125 1345 ;
    LAYER V1 ;
      RECT 11955 7055 12125 7225 ;
    LAYER V1 ;
      RECT 12815 1175 12985 1345 ;
    LAYER V1 ;
      RECT 12815 7055 12985 7225 ;
    LAYER V1 ;
      RECT 13675 1175 13845 1345 ;
    LAYER V1 ;
      RECT 13675 7055 13845 7225 ;
    LAYER V1 ;
      RECT 14535 1175 14705 1345 ;
    LAYER V1 ;
      RECT 14535 7055 14705 7225 ;
    LAYER V1 ;
      RECT 15395 1175 15565 1345 ;
    LAYER V1 ;
      RECT 15395 7055 15565 7225 ;
    LAYER V1 ;
      RECT 16255 1175 16425 1345 ;
    LAYER V1 ;
      RECT 16255 7055 16425 7225 ;
    LAYER V2 ;
      RECT 8095 345 8245 495 ;
    LAYER V2 ;
      RECT 8095 4545 8245 4695 ;
    LAYER V2 ;
      RECT 8095 6225 8245 6375 ;
    LAYER V2 ;
      RECT 8095 10425 8245 10575 ;
    LAYER V2 ;
      RECT 8525 765 8675 915 ;
    LAYER V2 ;
      RECT 8525 6645 8675 6795 ;
    LAYER V2 ;
      RECT 8955 1185 9105 1335 ;
    LAYER V2 ;
      RECT 8955 7065 9105 7215 ;
  END
END SCM_NMOS_B_8106910_X9_Y2
