# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18 ;
  ORIGIN -0.050000 -0.050000 ;
  SIZE  2.580000 BY  2.570000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.462000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 1.460000 2.630000 2.100000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.594000 ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.150000 1.845000 0.320000 ;
        RECT 0.835000 2.350000 1.845000 2.520000 ;
      LAYER mcon ;
        RECT 0.895000 0.150000 1.065000 0.320000 ;
        RECT 0.895000 2.350000 1.065000 2.520000 ;
        RECT 1.255000 0.150000 1.425000 0.320000 ;
        RECT 1.255000 2.350000 1.425000 2.520000 ;
        RECT 1.615000 0.150000 1.785000 0.320000 ;
        RECT 1.615000 2.350000 1.785000 2.520000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.835000 0.050000 1.845000 0.380000 ;
        RECT 0.835000 2.290000 1.845000 2.620000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.924000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.570000 2.630000 1.210000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  0.478500 ;
    PORT
      LAYER met1 ;
        RECT 0.180000 0.570000 0.470000 2.100000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.210000 0.570000 2.500000 2.100000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.660000 0.410000 2.010000 ;
      RECT 0.795000 0.490000 0.965000 2.180000 ;
      RECT 1.255000 0.490000 1.425000 2.180000 ;
      RECT 1.715000 0.490000 1.885000 2.180000 ;
      RECT 2.270000 0.660000 2.440000 2.010000 ;
    LAYER mcon ;
      RECT 0.240000 0.710000 0.410000 0.880000 ;
      RECT 0.240000 1.070000 0.410000 1.240000 ;
      RECT 0.240000 1.430000 0.410000 1.600000 ;
      RECT 0.240000 1.790000 0.410000 1.960000 ;
      RECT 0.795000 0.710000 0.965000 0.880000 ;
      RECT 0.795000 1.070000 0.965000 1.240000 ;
      RECT 0.795000 1.430000 0.965000 1.600000 ;
      RECT 0.795000 1.790000 0.965000 1.960000 ;
      RECT 1.255000 0.710000 1.425000 0.880000 ;
      RECT 1.255000 1.070000 1.425000 1.240000 ;
      RECT 1.255000 1.430000 1.425000 1.600000 ;
      RECT 1.255000 1.790000 1.425000 1.960000 ;
      RECT 1.715000 0.710000 1.885000 0.880000 ;
      RECT 1.715000 1.070000 1.885000 1.240000 ;
      RECT 1.715000 1.430000 1.885000 1.600000 ;
      RECT 1.715000 1.790000 1.885000 1.960000 ;
      RECT 2.270000 0.710000 2.440000 0.880000 ;
      RECT 2.270000 1.070000 2.440000 1.240000 ;
      RECT 2.270000 1.430000 2.440000 1.600000 ;
      RECT 2.270000 1.790000 2.440000 1.960000 ;
    LAYER met1 ;
      RECT 0.750000 0.570000 1.010000 2.100000 ;
      RECT 1.210000 0.570000 1.470000 2.100000 ;
      RECT 1.670000 0.570000 1.930000 2.100000 ;
    LAYER via ;
      RECT 0.750000 0.600000 1.010000 0.860000 ;
      RECT 0.750000 0.920000 1.010000 1.180000 ;
      RECT 1.210000 1.490000 1.470000 1.750000 ;
      RECT 1.210000 1.810000 1.470000 2.070000 ;
      RECT 1.670000 0.600000 1.930000 0.860000 ;
      RECT 1.670000 0.920000 1.930000 1.180000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18
END LIBRARY
