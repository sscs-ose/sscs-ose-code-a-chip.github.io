magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< error_p >>
rect -29 26143 29 26149
rect -29 26109 -17 26143
rect -29 26103 29 26109
rect -29 23633 29 23639
rect -29 23599 -17 23633
rect -29 23593 29 23599
rect -29 23525 29 23531
rect -29 23491 -17 23525
rect -29 23485 29 23491
rect -29 21015 29 21021
rect -29 20981 -17 21015
rect -29 20975 29 20981
rect -29 20907 29 20913
rect -29 20873 -17 20907
rect -29 20867 29 20873
rect -29 18397 29 18403
rect -29 18363 -17 18397
rect -29 18357 29 18363
rect -29 18289 29 18295
rect -29 18255 -17 18289
rect -29 18249 29 18255
rect -29 15779 29 15785
rect -29 15745 -17 15779
rect -29 15739 29 15745
rect -29 15671 29 15677
rect -29 15637 -17 15671
rect -29 15631 29 15637
rect -29 13161 29 13167
rect -29 13127 -17 13161
rect -29 13121 29 13127
rect -29 13053 29 13059
rect -29 13019 -17 13053
rect -29 13013 29 13019
rect -29 10543 29 10549
rect -29 10509 -17 10543
rect -29 10503 29 10509
rect -29 10435 29 10441
rect -29 10401 -17 10435
rect -29 10395 29 10401
rect -29 7925 29 7931
rect -29 7891 -17 7925
rect -29 7885 29 7891
rect -29 7817 29 7823
rect -29 7783 -17 7817
rect -29 7777 29 7783
rect -29 5307 29 5313
rect -29 5273 -17 5307
rect -29 5267 29 5273
rect -29 5199 29 5205
rect -29 5165 -17 5199
rect -29 5159 29 5165
rect -29 2689 29 2695
rect -29 2655 -17 2689
rect -29 2649 29 2655
rect -29 2581 29 2587
rect -29 2547 -17 2581
rect -29 2541 29 2547
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -2547 29 -2541
rect -29 -2581 -17 -2547
rect -29 -2587 29 -2581
rect -29 -2655 29 -2649
rect -29 -2689 -17 -2655
rect -29 -2695 29 -2689
rect -29 -5165 29 -5159
rect -29 -5199 -17 -5165
rect -29 -5205 29 -5199
rect -29 -5273 29 -5267
rect -29 -5307 -17 -5273
rect -29 -5313 29 -5307
rect -29 -7783 29 -7777
rect -29 -7817 -17 -7783
rect -29 -7823 29 -7817
rect -29 -7891 29 -7885
rect -29 -7925 -17 -7891
rect -29 -7931 29 -7925
rect -29 -10401 29 -10395
rect -29 -10435 -17 -10401
rect -29 -10441 29 -10435
rect -29 -10509 29 -10503
rect -29 -10543 -17 -10509
rect -29 -10549 29 -10543
rect -29 -13019 29 -13013
rect -29 -13053 -17 -13019
rect -29 -13059 29 -13053
rect -29 -13127 29 -13121
rect -29 -13161 -17 -13127
rect -29 -13167 29 -13161
rect -29 -15637 29 -15631
rect -29 -15671 -17 -15637
rect -29 -15677 29 -15671
rect -29 -15745 29 -15739
rect -29 -15779 -17 -15745
rect -29 -15785 29 -15779
rect -29 -18255 29 -18249
rect -29 -18289 -17 -18255
rect -29 -18295 29 -18289
rect -29 -18363 29 -18357
rect -29 -18397 -17 -18363
rect -29 -18403 29 -18397
rect -29 -20873 29 -20867
rect -29 -20907 -17 -20873
rect -29 -20913 29 -20907
rect -29 -20981 29 -20975
rect -29 -21015 -17 -20981
rect -29 -21021 29 -21015
rect -29 -23491 29 -23485
rect -29 -23525 -17 -23491
rect -29 -23531 29 -23525
rect -29 -23599 29 -23593
rect -29 -23633 -17 -23599
rect -29 -23639 29 -23633
rect -29 -26109 29 -26103
rect -29 -26143 -17 -26109
rect -29 -26149 29 -26143
<< pwell >>
rect -211 -26281 211 26281
<< nmos >>
rect -15 23671 15 26071
rect -15 21053 15 23453
rect -15 18435 15 20835
rect -15 15817 15 18217
rect -15 13199 15 15599
rect -15 10581 15 12981
rect -15 7963 15 10363
rect -15 5345 15 7745
rect -15 2727 15 5127
rect -15 109 15 2509
rect -15 -2509 15 -109
rect -15 -5127 15 -2727
rect -15 -7745 15 -5345
rect -15 -10363 15 -7963
rect -15 -12981 15 -10581
rect -15 -15599 15 -13199
rect -15 -18217 15 -15817
rect -15 -20835 15 -18435
rect -15 -23453 15 -21053
rect -15 -26071 15 -23671
<< ndiff >>
rect -73 26059 -15 26071
rect -73 23683 -61 26059
rect -27 23683 -15 26059
rect -73 23671 -15 23683
rect 15 26059 73 26071
rect 15 23683 27 26059
rect 61 23683 73 26059
rect 15 23671 73 23683
rect -73 23441 -15 23453
rect -73 21065 -61 23441
rect -27 21065 -15 23441
rect -73 21053 -15 21065
rect 15 23441 73 23453
rect 15 21065 27 23441
rect 61 21065 73 23441
rect 15 21053 73 21065
rect -73 20823 -15 20835
rect -73 18447 -61 20823
rect -27 18447 -15 20823
rect -73 18435 -15 18447
rect 15 20823 73 20835
rect 15 18447 27 20823
rect 61 18447 73 20823
rect 15 18435 73 18447
rect -73 18205 -15 18217
rect -73 15829 -61 18205
rect -27 15829 -15 18205
rect -73 15817 -15 15829
rect 15 18205 73 18217
rect 15 15829 27 18205
rect 61 15829 73 18205
rect 15 15817 73 15829
rect -73 15587 -15 15599
rect -73 13211 -61 15587
rect -27 13211 -15 15587
rect -73 13199 -15 13211
rect 15 15587 73 15599
rect 15 13211 27 15587
rect 61 13211 73 15587
rect 15 13199 73 13211
rect -73 12969 -15 12981
rect -73 10593 -61 12969
rect -27 10593 -15 12969
rect -73 10581 -15 10593
rect 15 12969 73 12981
rect 15 10593 27 12969
rect 61 10593 73 12969
rect 15 10581 73 10593
rect -73 10351 -15 10363
rect -73 7975 -61 10351
rect -27 7975 -15 10351
rect -73 7963 -15 7975
rect 15 10351 73 10363
rect 15 7975 27 10351
rect 61 7975 73 10351
rect 15 7963 73 7975
rect -73 7733 -15 7745
rect -73 5357 -61 7733
rect -27 5357 -15 7733
rect -73 5345 -15 5357
rect 15 7733 73 7745
rect 15 5357 27 7733
rect 61 5357 73 7733
rect 15 5345 73 5357
rect -73 5115 -15 5127
rect -73 2739 -61 5115
rect -27 2739 -15 5115
rect -73 2727 -15 2739
rect 15 5115 73 5127
rect 15 2739 27 5115
rect 61 2739 73 5115
rect 15 2727 73 2739
rect -73 2497 -15 2509
rect -73 121 -61 2497
rect -27 121 -15 2497
rect -73 109 -15 121
rect 15 2497 73 2509
rect 15 121 27 2497
rect 61 121 73 2497
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -2497 -61 -121
rect -27 -2497 -15 -121
rect -73 -2509 -15 -2497
rect 15 -121 73 -109
rect 15 -2497 27 -121
rect 61 -2497 73 -121
rect 15 -2509 73 -2497
rect -73 -2739 -15 -2727
rect -73 -5115 -61 -2739
rect -27 -5115 -15 -2739
rect -73 -5127 -15 -5115
rect 15 -2739 73 -2727
rect 15 -5115 27 -2739
rect 61 -5115 73 -2739
rect 15 -5127 73 -5115
rect -73 -5357 -15 -5345
rect -73 -7733 -61 -5357
rect -27 -7733 -15 -5357
rect -73 -7745 -15 -7733
rect 15 -5357 73 -5345
rect 15 -7733 27 -5357
rect 61 -7733 73 -5357
rect 15 -7745 73 -7733
rect -73 -7975 -15 -7963
rect -73 -10351 -61 -7975
rect -27 -10351 -15 -7975
rect -73 -10363 -15 -10351
rect 15 -7975 73 -7963
rect 15 -10351 27 -7975
rect 61 -10351 73 -7975
rect 15 -10363 73 -10351
rect -73 -10593 -15 -10581
rect -73 -12969 -61 -10593
rect -27 -12969 -15 -10593
rect -73 -12981 -15 -12969
rect 15 -10593 73 -10581
rect 15 -12969 27 -10593
rect 61 -12969 73 -10593
rect 15 -12981 73 -12969
rect -73 -13211 -15 -13199
rect -73 -15587 -61 -13211
rect -27 -15587 -15 -13211
rect -73 -15599 -15 -15587
rect 15 -13211 73 -13199
rect 15 -15587 27 -13211
rect 61 -15587 73 -13211
rect 15 -15599 73 -15587
rect -73 -15829 -15 -15817
rect -73 -18205 -61 -15829
rect -27 -18205 -15 -15829
rect -73 -18217 -15 -18205
rect 15 -15829 73 -15817
rect 15 -18205 27 -15829
rect 61 -18205 73 -15829
rect 15 -18217 73 -18205
rect -73 -18447 -15 -18435
rect -73 -20823 -61 -18447
rect -27 -20823 -15 -18447
rect -73 -20835 -15 -20823
rect 15 -18447 73 -18435
rect 15 -20823 27 -18447
rect 61 -20823 73 -18447
rect 15 -20835 73 -20823
rect -73 -21065 -15 -21053
rect -73 -23441 -61 -21065
rect -27 -23441 -15 -21065
rect -73 -23453 -15 -23441
rect 15 -21065 73 -21053
rect 15 -23441 27 -21065
rect 61 -23441 73 -21065
rect 15 -23453 73 -23441
rect -73 -23683 -15 -23671
rect -73 -26059 -61 -23683
rect -27 -26059 -15 -23683
rect -73 -26071 -15 -26059
rect 15 -23683 73 -23671
rect 15 -26059 27 -23683
rect 61 -26059 73 -23683
rect 15 -26071 73 -26059
<< ndiffc >>
rect -61 23683 -27 26059
rect 27 23683 61 26059
rect -61 21065 -27 23441
rect 27 21065 61 23441
rect -61 18447 -27 20823
rect 27 18447 61 20823
rect -61 15829 -27 18205
rect 27 15829 61 18205
rect -61 13211 -27 15587
rect 27 13211 61 15587
rect -61 10593 -27 12969
rect 27 10593 61 12969
rect -61 7975 -27 10351
rect 27 7975 61 10351
rect -61 5357 -27 7733
rect 27 5357 61 7733
rect -61 2739 -27 5115
rect 27 2739 61 5115
rect -61 121 -27 2497
rect 27 121 61 2497
rect -61 -2497 -27 -121
rect 27 -2497 61 -121
rect -61 -5115 -27 -2739
rect 27 -5115 61 -2739
rect -61 -7733 -27 -5357
rect 27 -7733 61 -5357
rect -61 -10351 -27 -7975
rect 27 -10351 61 -7975
rect -61 -12969 -27 -10593
rect 27 -12969 61 -10593
rect -61 -15587 -27 -13211
rect 27 -15587 61 -13211
rect -61 -18205 -27 -15829
rect 27 -18205 61 -15829
rect -61 -20823 -27 -18447
rect 27 -20823 61 -18447
rect -61 -23441 -27 -21065
rect 27 -23441 61 -21065
rect -61 -26059 -27 -23683
rect 27 -26059 61 -23683
<< psubdiff >>
rect -175 26211 -79 26245
rect 79 26211 175 26245
rect -175 26149 -141 26211
rect 141 26149 175 26211
rect -175 -26211 -141 -26149
rect 141 -26211 175 -26149
rect -175 -26245 -79 -26211
rect 79 -26245 175 -26211
<< psubdiffcont >>
rect -79 26211 79 26245
rect -175 -26149 -141 26149
rect 141 -26149 175 26149
rect -79 -26245 79 -26211
<< poly >>
rect -33 26143 33 26159
rect -33 26109 -17 26143
rect 17 26109 33 26143
rect -33 26093 33 26109
rect -15 26071 15 26093
rect -15 23649 15 23671
rect -33 23633 33 23649
rect -33 23599 -17 23633
rect 17 23599 33 23633
rect -33 23583 33 23599
rect -33 23525 33 23541
rect -33 23491 -17 23525
rect 17 23491 33 23525
rect -33 23475 33 23491
rect -15 23453 15 23475
rect -15 21031 15 21053
rect -33 21015 33 21031
rect -33 20981 -17 21015
rect 17 20981 33 21015
rect -33 20965 33 20981
rect -33 20907 33 20923
rect -33 20873 -17 20907
rect 17 20873 33 20907
rect -33 20857 33 20873
rect -15 20835 15 20857
rect -15 18413 15 18435
rect -33 18397 33 18413
rect -33 18363 -17 18397
rect 17 18363 33 18397
rect -33 18347 33 18363
rect -33 18289 33 18305
rect -33 18255 -17 18289
rect 17 18255 33 18289
rect -33 18239 33 18255
rect -15 18217 15 18239
rect -15 15795 15 15817
rect -33 15779 33 15795
rect -33 15745 -17 15779
rect 17 15745 33 15779
rect -33 15729 33 15745
rect -33 15671 33 15687
rect -33 15637 -17 15671
rect 17 15637 33 15671
rect -33 15621 33 15637
rect -15 15599 15 15621
rect -15 13177 15 13199
rect -33 13161 33 13177
rect -33 13127 -17 13161
rect 17 13127 33 13161
rect -33 13111 33 13127
rect -33 13053 33 13069
rect -33 13019 -17 13053
rect 17 13019 33 13053
rect -33 13003 33 13019
rect -15 12981 15 13003
rect -15 10559 15 10581
rect -33 10543 33 10559
rect -33 10509 -17 10543
rect 17 10509 33 10543
rect -33 10493 33 10509
rect -33 10435 33 10451
rect -33 10401 -17 10435
rect 17 10401 33 10435
rect -33 10385 33 10401
rect -15 10363 15 10385
rect -15 7941 15 7963
rect -33 7925 33 7941
rect -33 7891 -17 7925
rect 17 7891 33 7925
rect -33 7875 33 7891
rect -33 7817 33 7833
rect -33 7783 -17 7817
rect 17 7783 33 7817
rect -33 7767 33 7783
rect -15 7745 15 7767
rect -15 5323 15 5345
rect -33 5307 33 5323
rect -33 5273 -17 5307
rect 17 5273 33 5307
rect -33 5257 33 5273
rect -33 5199 33 5215
rect -33 5165 -17 5199
rect 17 5165 33 5199
rect -33 5149 33 5165
rect -15 5127 15 5149
rect -15 2705 15 2727
rect -33 2689 33 2705
rect -33 2655 -17 2689
rect 17 2655 33 2689
rect -33 2639 33 2655
rect -33 2581 33 2597
rect -33 2547 -17 2581
rect 17 2547 33 2581
rect -33 2531 33 2547
rect -15 2509 15 2531
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -2531 15 -2509
rect -33 -2547 33 -2531
rect -33 -2581 -17 -2547
rect 17 -2581 33 -2547
rect -33 -2597 33 -2581
rect -33 -2655 33 -2639
rect -33 -2689 -17 -2655
rect 17 -2689 33 -2655
rect -33 -2705 33 -2689
rect -15 -2727 15 -2705
rect -15 -5149 15 -5127
rect -33 -5165 33 -5149
rect -33 -5199 -17 -5165
rect 17 -5199 33 -5165
rect -33 -5215 33 -5199
rect -33 -5273 33 -5257
rect -33 -5307 -17 -5273
rect 17 -5307 33 -5273
rect -33 -5323 33 -5307
rect -15 -5345 15 -5323
rect -15 -7767 15 -7745
rect -33 -7783 33 -7767
rect -33 -7817 -17 -7783
rect 17 -7817 33 -7783
rect -33 -7833 33 -7817
rect -33 -7891 33 -7875
rect -33 -7925 -17 -7891
rect 17 -7925 33 -7891
rect -33 -7941 33 -7925
rect -15 -7963 15 -7941
rect -15 -10385 15 -10363
rect -33 -10401 33 -10385
rect -33 -10435 -17 -10401
rect 17 -10435 33 -10401
rect -33 -10451 33 -10435
rect -33 -10509 33 -10493
rect -33 -10543 -17 -10509
rect 17 -10543 33 -10509
rect -33 -10559 33 -10543
rect -15 -10581 15 -10559
rect -15 -13003 15 -12981
rect -33 -13019 33 -13003
rect -33 -13053 -17 -13019
rect 17 -13053 33 -13019
rect -33 -13069 33 -13053
rect -33 -13127 33 -13111
rect -33 -13161 -17 -13127
rect 17 -13161 33 -13127
rect -33 -13177 33 -13161
rect -15 -13199 15 -13177
rect -15 -15621 15 -15599
rect -33 -15637 33 -15621
rect -33 -15671 -17 -15637
rect 17 -15671 33 -15637
rect -33 -15687 33 -15671
rect -33 -15745 33 -15729
rect -33 -15779 -17 -15745
rect 17 -15779 33 -15745
rect -33 -15795 33 -15779
rect -15 -15817 15 -15795
rect -15 -18239 15 -18217
rect -33 -18255 33 -18239
rect -33 -18289 -17 -18255
rect 17 -18289 33 -18255
rect -33 -18305 33 -18289
rect -33 -18363 33 -18347
rect -33 -18397 -17 -18363
rect 17 -18397 33 -18363
rect -33 -18413 33 -18397
rect -15 -18435 15 -18413
rect -15 -20857 15 -20835
rect -33 -20873 33 -20857
rect -33 -20907 -17 -20873
rect 17 -20907 33 -20873
rect -33 -20923 33 -20907
rect -33 -20981 33 -20965
rect -33 -21015 -17 -20981
rect 17 -21015 33 -20981
rect -33 -21031 33 -21015
rect -15 -21053 15 -21031
rect -15 -23475 15 -23453
rect -33 -23491 33 -23475
rect -33 -23525 -17 -23491
rect 17 -23525 33 -23491
rect -33 -23541 33 -23525
rect -33 -23599 33 -23583
rect -33 -23633 -17 -23599
rect 17 -23633 33 -23599
rect -33 -23649 33 -23633
rect -15 -23671 15 -23649
rect -15 -26093 15 -26071
rect -33 -26109 33 -26093
rect -33 -26143 -17 -26109
rect 17 -26143 33 -26109
rect -33 -26159 33 -26143
<< polycont >>
rect -17 26109 17 26143
rect -17 23599 17 23633
rect -17 23491 17 23525
rect -17 20981 17 21015
rect -17 20873 17 20907
rect -17 18363 17 18397
rect -17 18255 17 18289
rect -17 15745 17 15779
rect -17 15637 17 15671
rect -17 13127 17 13161
rect -17 13019 17 13053
rect -17 10509 17 10543
rect -17 10401 17 10435
rect -17 7891 17 7925
rect -17 7783 17 7817
rect -17 5273 17 5307
rect -17 5165 17 5199
rect -17 2655 17 2689
rect -17 2547 17 2581
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -2581 17 -2547
rect -17 -2689 17 -2655
rect -17 -5199 17 -5165
rect -17 -5307 17 -5273
rect -17 -7817 17 -7783
rect -17 -7925 17 -7891
rect -17 -10435 17 -10401
rect -17 -10543 17 -10509
rect -17 -13053 17 -13019
rect -17 -13161 17 -13127
rect -17 -15671 17 -15637
rect -17 -15779 17 -15745
rect -17 -18289 17 -18255
rect -17 -18397 17 -18363
rect -17 -20907 17 -20873
rect -17 -21015 17 -20981
rect -17 -23525 17 -23491
rect -17 -23633 17 -23599
rect -17 -26143 17 -26109
<< locali >>
rect -175 26211 -79 26245
rect 79 26211 175 26245
rect -175 26149 -141 26211
rect 141 26149 175 26211
rect -33 26109 -17 26143
rect 17 26109 33 26143
rect -61 26059 -27 26075
rect -61 23667 -27 23683
rect 27 26059 61 26075
rect 27 23667 61 23683
rect -33 23599 -17 23633
rect 17 23599 33 23633
rect -33 23491 -17 23525
rect 17 23491 33 23525
rect -61 23441 -27 23457
rect -61 21049 -27 21065
rect 27 23441 61 23457
rect 27 21049 61 21065
rect -33 20981 -17 21015
rect 17 20981 33 21015
rect -33 20873 -17 20907
rect 17 20873 33 20907
rect -61 20823 -27 20839
rect -61 18431 -27 18447
rect 27 20823 61 20839
rect 27 18431 61 18447
rect -33 18363 -17 18397
rect 17 18363 33 18397
rect -33 18255 -17 18289
rect 17 18255 33 18289
rect -61 18205 -27 18221
rect -61 15813 -27 15829
rect 27 18205 61 18221
rect 27 15813 61 15829
rect -33 15745 -17 15779
rect 17 15745 33 15779
rect -33 15637 -17 15671
rect 17 15637 33 15671
rect -61 15587 -27 15603
rect -61 13195 -27 13211
rect 27 15587 61 15603
rect 27 13195 61 13211
rect -33 13127 -17 13161
rect 17 13127 33 13161
rect -33 13019 -17 13053
rect 17 13019 33 13053
rect -61 12969 -27 12985
rect -61 10577 -27 10593
rect 27 12969 61 12985
rect 27 10577 61 10593
rect -33 10509 -17 10543
rect 17 10509 33 10543
rect -33 10401 -17 10435
rect 17 10401 33 10435
rect -61 10351 -27 10367
rect -61 7959 -27 7975
rect 27 10351 61 10367
rect 27 7959 61 7975
rect -33 7891 -17 7925
rect 17 7891 33 7925
rect -33 7783 -17 7817
rect 17 7783 33 7817
rect -61 7733 -27 7749
rect -61 5341 -27 5357
rect 27 7733 61 7749
rect 27 5341 61 5357
rect -33 5273 -17 5307
rect 17 5273 33 5307
rect -33 5165 -17 5199
rect 17 5165 33 5199
rect -61 5115 -27 5131
rect -61 2723 -27 2739
rect 27 5115 61 5131
rect 27 2723 61 2739
rect -33 2655 -17 2689
rect 17 2655 33 2689
rect -33 2547 -17 2581
rect 17 2547 33 2581
rect -61 2497 -27 2513
rect -61 105 -27 121
rect 27 2497 61 2513
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -2513 -27 -2497
rect 27 -121 61 -105
rect 27 -2513 61 -2497
rect -33 -2581 -17 -2547
rect 17 -2581 33 -2547
rect -33 -2689 -17 -2655
rect 17 -2689 33 -2655
rect -61 -2739 -27 -2723
rect -61 -5131 -27 -5115
rect 27 -2739 61 -2723
rect 27 -5131 61 -5115
rect -33 -5199 -17 -5165
rect 17 -5199 33 -5165
rect -33 -5307 -17 -5273
rect 17 -5307 33 -5273
rect -61 -5357 -27 -5341
rect -61 -7749 -27 -7733
rect 27 -5357 61 -5341
rect 27 -7749 61 -7733
rect -33 -7817 -17 -7783
rect 17 -7817 33 -7783
rect -33 -7925 -17 -7891
rect 17 -7925 33 -7891
rect -61 -7975 -27 -7959
rect -61 -10367 -27 -10351
rect 27 -7975 61 -7959
rect 27 -10367 61 -10351
rect -33 -10435 -17 -10401
rect 17 -10435 33 -10401
rect -33 -10543 -17 -10509
rect 17 -10543 33 -10509
rect -61 -10593 -27 -10577
rect -61 -12985 -27 -12969
rect 27 -10593 61 -10577
rect 27 -12985 61 -12969
rect -33 -13053 -17 -13019
rect 17 -13053 33 -13019
rect -33 -13161 -17 -13127
rect 17 -13161 33 -13127
rect -61 -13211 -27 -13195
rect -61 -15603 -27 -15587
rect 27 -13211 61 -13195
rect 27 -15603 61 -15587
rect -33 -15671 -17 -15637
rect 17 -15671 33 -15637
rect -33 -15779 -17 -15745
rect 17 -15779 33 -15745
rect -61 -15829 -27 -15813
rect -61 -18221 -27 -18205
rect 27 -15829 61 -15813
rect 27 -18221 61 -18205
rect -33 -18289 -17 -18255
rect 17 -18289 33 -18255
rect -33 -18397 -17 -18363
rect 17 -18397 33 -18363
rect -61 -18447 -27 -18431
rect -61 -20839 -27 -20823
rect 27 -18447 61 -18431
rect 27 -20839 61 -20823
rect -33 -20907 -17 -20873
rect 17 -20907 33 -20873
rect -33 -21015 -17 -20981
rect 17 -21015 33 -20981
rect -61 -21065 -27 -21049
rect -61 -23457 -27 -23441
rect 27 -21065 61 -21049
rect 27 -23457 61 -23441
rect -33 -23525 -17 -23491
rect 17 -23525 33 -23491
rect -33 -23633 -17 -23599
rect 17 -23633 33 -23599
rect -61 -23683 -27 -23667
rect -61 -26075 -27 -26059
rect 27 -23683 61 -23667
rect 27 -26075 61 -26059
rect -33 -26143 -17 -26109
rect 17 -26143 33 -26109
rect -175 -26211 -141 -26149
rect 141 -26211 175 -26149
rect -175 -26245 -79 -26211
rect 79 -26245 175 -26211
<< viali >>
rect -17 26109 17 26143
rect -61 23683 -27 26059
rect 27 23683 61 26059
rect -17 23599 17 23633
rect -17 23491 17 23525
rect -61 21065 -27 23441
rect 27 21065 61 23441
rect -17 20981 17 21015
rect -17 20873 17 20907
rect -61 18447 -27 20823
rect 27 18447 61 20823
rect -17 18363 17 18397
rect -17 18255 17 18289
rect -61 15829 -27 18205
rect 27 15829 61 18205
rect -17 15745 17 15779
rect -17 15637 17 15671
rect -61 13211 -27 15587
rect 27 13211 61 15587
rect -17 13127 17 13161
rect -17 13019 17 13053
rect -61 10593 -27 12969
rect 27 10593 61 12969
rect -17 10509 17 10543
rect -17 10401 17 10435
rect -61 7975 -27 10351
rect 27 7975 61 10351
rect -17 7891 17 7925
rect -17 7783 17 7817
rect -61 5357 -27 7733
rect 27 5357 61 7733
rect -17 5273 17 5307
rect -17 5165 17 5199
rect -61 2739 -27 5115
rect 27 2739 61 5115
rect -17 2655 17 2689
rect -17 2547 17 2581
rect -61 121 -27 2497
rect 27 121 61 2497
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -2497 -27 -121
rect 27 -2497 61 -121
rect -17 -2581 17 -2547
rect -17 -2689 17 -2655
rect -61 -5115 -27 -2739
rect 27 -5115 61 -2739
rect -17 -5199 17 -5165
rect -17 -5307 17 -5273
rect -61 -7733 -27 -5357
rect 27 -7733 61 -5357
rect -17 -7817 17 -7783
rect -17 -7925 17 -7891
rect -61 -10351 -27 -7975
rect 27 -10351 61 -7975
rect -17 -10435 17 -10401
rect -17 -10543 17 -10509
rect -61 -12969 -27 -10593
rect 27 -12969 61 -10593
rect -17 -13053 17 -13019
rect -17 -13161 17 -13127
rect -61 -15587 -27 -13211
rect 27 -15587 61 -13211
rect -17 -15671 17 -15637
rect -17 -15779 17 -15745
rect -61 -18205 -27 -15829
rect 27 -18205 61 -15829
rect -17 -18289 17 -18255
rect -17 -18397 17 -18363
rect -61 -20823 -27 -18447
rect 27 -20823 61 -18447
rect -17 -20907 17 -20873
rect -17 -21015 17 -20981
rect -61 -23441 -27 -21065
rect 27 -23441 61 -21065
rect -17 -23525 17 -23491
rect -17 -23633 17 -23599
rect -61 -26059 -27 -23683
rect 27 -26059 61 -23683
rect -17 -26143 17 -26109
<< metal1 >>
rect -29 26143 29 26149
rect -29 26109 -17 26143
rect 17 26109 29 26143
rect -29 26103 29 26109
rect -67 26059 -21 26071
rect -67 23683 -61 26059
rect -27 23683 -21 26059
rect -67 23671 -21 23683
rect 21 26059 67 26071
rect 21 23683 27 26059
rect 61 23683 67 26059
rect 21 23671 67 23683
rect -29 23633 29 23639
rect -29 23599 -17 23633
rect 17 23599 29 23633
rect -29 23593 29 23599
rect -29 23525 29 23531
rect -29 23491 -17 23525
rect 17 23491 29 23525
rect -29 23485 29 23491
rect -67 23441 -21 23453
rect -67 21065 -61 23441
rect -27 21065 -21 23441
rect -67 21053 -21 21065
rect 21 23441 67 23453
rect 21 21065 27 23441
rect 61 21065 67 23441
rect 21 21053 67 21065
rect -29 21015 29 21021
rect -29 20981 -17 21015
rect 17 20981 29 21015
rect -29 20975 29 20981
rect -29 20907 29 20913
rect -29 20873 -17 20907
rect 17 20873 29 20907
rect -29 20867 29 20873
rect -67 20823 -21 20835
rect -67 18447 -61 20823
rect -27 18447 -21 20823
rect -67 18435 -21 18447
rect 21 20823 67 20835
rect 21 18447 27 20823
rect 61 18447 67 20823
rect 21 18435 67 18447
rect -29 18397 29 18403
rect -29 18363 -17 18397
rect 17 18363 29 18397
rect -29 18357 29 18363
rect -29 18289 29 18295
rect -29 18255 -17 18289
rect 17 18255 29 18289
rect -29 18249 29 18255
rect -67 18205 -21 18217
rect -67 15829 -61 18205
rect -27 15829 -21 18205
rect -67 15817 -21 15829
rect 21 18205 67 18217
rect 21 15829 27 18205
rect 61 15829 67 18205
rect 21 15817 67 15829
rect -29 15779 29 15785
rect -29 15745 -17 15779
rect 17 15745 29 15779
rect -29 15739 29 15745
rect -29 15671 29 15677
rect -29 15637 -17 15671
rect 17 15637 29 15671
rect -29 15631 29 15637
rect -67 15587 -21 15599
rect -67 13211 -61 15587
rect -27 13211 -21 15587
rect -67 13199 -21 13211
rect 21 15587 67 15599
rect 21 13211 27 15587
rect 61 13211 67 15587
rect 21 13199 67 13211
rect -29 13161 29 13167
rect -29 13127 -17 13161
rect 17 13127 29 13161
rect -29 13121 29 13127
rect -29 13053 29 13059
rect -29 13019 -17 13053
rect 17 13019 29 13053
rect -29 13013 29 13019
rect -67 12969 -21 12981
rect -67 10593 -61 12969
rect -27 10593 -21 12969
rect -67 10581 -21 10593
rect 21 12969 67 12981
rect 21 10593 27 12969
rect 61 10593 67 12969
rect 21 10581 67 10593
rect -29 10543 29 10549
rect -29 10509 -17 10543
rect 17 10509 29 10543
rect -29 10503 29 10509
rect -29 10435 29 10441
rect -29 10401 -17 10435
rect 17 10401 29 10435
rect -29 10395 29 10401
rect -67 10351 -21 10363
rect -67 7975 -61 10351
rect -27 7975 -21 10351
rect -67 7963 -21 7975
rect 21 10351 67 10363
rect 21 7975 27 10351
rect 61 7975 67 10351
rect 21 7963 67 7975
rect -29 7925 29 7931
rect -29 7891 -17 7925
rect 17 7891 29 7925
rect -29 7885 29 7891
rect -29 7817 29 7823
rect -29 7783 -17 7817
rect 17 7783 29 7817
rect -29 7777 29 7783
rect -67 7733 -21 7745
rect -67 5357 -61 7733
rect -27 5357 -21 7733
rect -67 5345 -21 5357
rect 21 7733 67 7745
rect 21 5357 27 7733
rect 61 5357 67 7733
rect 21 5345 67 5357
rect -29 5307 29 5313
rect -29 5273 -17 5307
rect 17 5273 29 5307
rect -29 5267 29 5273
rect -29 5199 29 5205
rect -29 5165 -17 5199
rect 17 5165 29 5199
rect -29 5159 29 5165
rect -67 5115 -21 5127
rect -67 2739 -61 5115
rect -27 2739 -21 5115
rect -67 2727 -21 2739
rect 21 5115 67 5127
rect 21 2739 27 5115
rect 61 2739 67 5115
rect 21 2727 67 2739
rect -29 2689 29 2695
rect -29 2655 -17 2689
rect 17 2655 29 2689
rect -29 2649 29 2655
rect -29 2581 29 2587
rect -29 2547 -17 2581
rect 17 2547 29 2581
rect -29 2541 29 2547
rect -67 2497 -21 2509
rect -67 121 -61 2497
rect -27 121 -21 2497
rect -67 109 -21 121
rect 21 2497 67 2509
rect 21 121 27 2497
rect 61 121 67 2497
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -2497 -61 -121
rect -27 -2497 -21 -121
rect -67 -2509 -21 -2497
rect 21 -121 67 -109
rect 21 -2497 27 -121
rect 61 -2497 67 -121
rect 21 -2509 67 -2497
rect -29 -2547 29 -2541
rect -29 -2581 -17 -2547
rect 17 -2581 29 -2547
rect -29 -2587 29 -2581
rect -29 -2655 29 -2649
rect -29 -2689 -17 -2655
rect 17 -2689 29 -2655
rect -29 -2695 29 -2689
rect -67 -2739 -21 -2727
rect -67 -5115 -61 -2739
rect -27 -5115 -21 -2739
rect -67 -5127 -21 -5115
rect 21 -2739 67 -2727
rect 21 -5115 27 -2739
rect 61 -5115 67 -2739
rect 21 -5127 67 -5115
rect -29 -5165 29 -5159
rect -29 -5199 -17 -5165
rect 17 -5199 29 -5165
rect -29 -5205 29 -5199
rect -29 -5273 29 -5267
rect -29 -5307 -17 -5273
rect 17 -5307 29 -5273
rect -29 -5313 29 -5307
rect -67 -5357 -21 -5345
rect -67 -7733 -61 -5357
rect -27 -7733 -21 -5357
rect -67 -7745 -21 -7733
rect 21 -5357 67 -5345
rect 21 -7733 27 -5357
rect 61 -7733 67 -5357
rect 21 -7745 67 -7733
rect -29 -7783 29 -7777
rect -29 -7817 -17 -7783
rect 17 -7817 29 -7783
rect -29 -7823 29 -7817
rect -29 -7891 29 -7885
rect -29 -7925 -17 -7891
rect 17 -7925 29 -7891
rect -29 -7931 29 -7925
rect -67 -7975 -21 -7963
rect -67 -10351 -61 -7975
rect -27 -10351 -21 -7975
rect -67 -10363 -21 -10351
rect 21 -7975 67 -7963
rect 21 -10351 27 -7975
rect 61 -10351 67 -7975
rect 21 -10363 67 -10351
rect -29 -10401 29 -10395
rect -29 -10435 -17 -10401
rect 17 -10435 29 -10401
rect -29 -10441 29 -10435
rect -29 -10509 29 -10503
rect -29 -10543 -17 -10509
rect 17 -10543 29 -10509
rect -29 -10549 29 -10543
rect -67 -10593 -21 -10581
rect -67 -12969 -61 -10593
rect -27 -12969 -21 -10593
rect -67 -12981 -21 -12969
rect 21 -10593 67 -10581
rect 21 -12969 27 -10593
rect 61 -12969 67 -10593
rect 21 -12981 67 -12969
rect -29 -13019 29 -13013
rect -29 -13053 -17 -13019
rect 17 -13053 29 -13019
rect -29 -13059 29 -13053
rect -29 -13127 29 -13121
rect -29 -13161 -17 -13127
rect 17 -13161 29 -13127
rect -29 -13167 29 -13161
rect -67 -13211 -21 -13199
rect -67 -15587 -61 -13211
rect -27 -15587 -21 -13211
rect -67 -15599 -21 -15587
rect 21 -13211 67 -13199
rect 21 -15587 27 -13211
rect 61 -15587 67 -13211
rect 21 -15599 67 -15587
rect -29 -15637 29 -15631
rect -29 -15671 -17 -15637
rect 17 -15671 29 -15637
rect -29 -15677 29 -15671
rect -29 -15745 29 -15739
rect -29 -15779 -17 -15745
rect 17 -15779 29 -15745
rect -29 -15785 29 -15779
rect -67 -15829 -21 -15817
rect -67 -18205 -61 -15829
rect -27 -18205 -21 -15829
rect -67 -18217 -21 -18205
rect 21 -15829 67 -15817
rect 21 -18205 27 -15829
rect 61 -18205 67 -15829
rect 21 -18217 67 -18205
rect -29 -18255 29 -18249
rect -29 -18289 -17 -18255
rect 17 -18289 29 -18255
rect -29 -18295 29 -18289
rect -29 -18363 29 -18357
rect -29 -18397 -17 -18363
rect 17 -18397 29 -18363
rect -29 -18403 29 -18397
rect -67 -18447 -21 -18435
rect -67 -20823 -61 -18447
rect -27 -20823 -21 -18447
rect -67 -20835 -21 -20823
rect 21 -18447 67 -18435
rect 21 -20823 27 -18447
rect 61 -20823 67 -18447
rect 21 -20835 67 -20823
rect -29 -20873 29 -20867
rect -29 -20907 -17 -20873
rect 17 -20907 29 -20873
rect -29 -20913 29 -20907
rect -29 -20981 29 -20975
rect -29 -21015 -17 -20981
rect 17 -21015 29 -20981
rect -29 -21021 29 -21015
rect -67 -21065 -21 -21053
rect -67 -23441 -61 -21065
rect -27 -23441 -21 -21065
rect -67 -23453 -21 -23441
rect 21 -21065 67 -21053
rect 21 -23441 27 -21065
rect 61 -23441 67 -21065
rect 21 -23453 67 -23441
rect -29 -23491 29 -23485
rect -29 -23525 -17 -23491
rect 17 -23525 29 -23491
rect -29 -23531 29 -23525
rect -29 -23599 29 -23593
rect -29 -23633 -17 -23599
rect 17 -23633 29 -23599
rect -29 -23639 29 -23633
rect -67 -23683 -21 -23671
rect -67 -26059 -61 -23683
rect -27 -26059 -21 -23683
rect -67 -26071 -21 -26059
rect 21 -23683 67 -23671
rect 21 -26059 27 -23683
rect 61 -26059 67 -23683
rect 21 -26071 67 -26059
rect -29 -26109 29 -26103
rect -29 -26143 -17 -26109
rect 17 -26143 29 -26109
rect -29 -26149 29 -26143
<< labels >>
rlabel psubdiffcont 0 -26228 0 -26228 0 B
port 1 nsew
rlabel ndiffc -44 -24871 -44 -24871 0 D0
port 2 nsew
rlabel ndiffc 44 -24871 44 -24871 0 S0
port 3 nsew
rlabel polycont 0 -23616 0 -23616 0 G0
port 4 nsew
rlabel ndiffc -44 -22253 -44 -22253 0 D1
port 5 nsew
rlabel ndiffc 44 -22253 44 -22253 0 S1
port 6 nsew
rlabel polycont 0 -20998 0 -20998 0 G1
port 7 nsew
rlabel ndiffc -44 -19635 -44 -19635 0 D2
port 8 nsew
rlabel ndiffc 44 -19635 44 -19635 0 S2
port 9 nsew
rlabel polycont 0 -18380 0 -18380 0 G2
port 10 nsew
rlabel ndiffc -44 -17017 -44 -17017 0 D3
port 11 nsew
rlabel ndiffc 44 -17017 44 -17017 0 S3
port 12 nsew
rlabel polycont 0 -15762 0 -15762 0 G3
port 13 nsew
rlabel ndiffc -44 -14399 -44 -14399 0 D4
port 14 nsew
rlabel ndiffc 44 -14399 44 -14399 0 S4
port 15 nsew
rlabel polycont 0 -13144 0 -13144 0 G4
port 16 nsew
rlabel ndiffc -44 -11781 -44 -11781 0 D5
port 17 nsew
rlabel ndiffc 44 -11781 44 -11781 0 S5
port 18 nsew
rlabel polycont 0 -10526 0 -10526 0 G5
port 19 nsew
rlabel ndiffc -44 -9163 -44 -9163 0 D6
port 20 nsew
rlabel ndiffc 44 -9163 44 -9163 0 S6
port 21 nsew
rlabel polycont 0 -7908 0 -7908 0 G6
port 22 nsew
rlabel ndiffc -44 -6545 -44 -6545 0 D7
port 23 nsew
rlabel ndiffc 44 -6545 44 -6545 0 S7
port 24 nsew
rlabel polycont 0 -5290 0 -5290 0 G7
port 25 nsew
rlabel ndiffc -44 -3927 -44 -3927 0 D8
port 26 nsew
rlabel ndiffc 44 -3927 44 -3927 0 S8
port 27 nsew
rlabel polycont 0 -2672 0 -2672 0 G8
port 28 nsew
rlabel ndiffc -44 -1309 -44 -1309 0 D9
port 29 nsew
rlabel ndiffc 44 -1309 44 -1309 0 S9
port 30 nsew
rlabel polycont 0 -54 0 -54 0 G9
port 31 nsew
rlabel ndiffc -44 1309 -44 1309 0 D10
port 32 nsew
rlabel ndiffc 44 1309 44 1309 0 S10
port 33 nsew
rlabel polycont 0 2564 0 2564 0 G10
port 34 nsew
rlabel ndiffc -44 3927 -44 3927 0 D11
port 35 nsew
rlabel ndiffc 44 3927 44 3927 0 S11
port 36 nsew
rlabel polycont 0 5182 0 5182 0 G11
port 37 nsew
rlabel ndiffc -44 6545 -44 6545 0 D12
port 38 nsew
rlabel ndiffc 44 6545 44 6545 0 S12
port 39 nsew
rlabel polycont 0 7800 0 7800 0 G12
port 40 nsew
rlabel ndiffc -44 9163 -44 9163 0 D13
port 41 nsew
rlabel ndiffc 44 9163 44 9163 0 S13
port 42 nsew
rlabel polycont 0 10418 0 10418 0 G13
port 43 nsew
rlabel ndiffc -44 11781 -44 11781 0 D14
port 44 nsew
rlabel ndiffc 44 11781 44 11781 0 S14
port 45 nsew
rlabel polycont 0 13036 0 13036 0 G14
port 46 nsew
rlabel ndiffc -44 14399 -44 14399 0 D15
port 47 nsew
rlabel ndiffc 44 14399 44 14399 0 S15
port 48 nsew
rlabel polycont 0 15654 0 15654 0 G15
port 49 nsew
rlabel ndiffc -44 17017 -44 17017 0 D16
port 50 nsew
rlabel ndiffc 44 17017 44 17017 0 S16
port 51 nsew
rlabel polycont 0 18272 0 18272 0 G16
port 52 nsew
rlabel ndiffc -44 19635 -44 19635 0 D17
port 53 nsew
rlabel ndiffc 44 19635 44 19635 0 S17
port 54 nsew
rlabel polycont 0 20890 0 20890 0 G17
port 55 nsew
rlabel ndiffc -44 22253 -44 22253 0 D18
port 56 nsew
rlabel ndiffc 44 22253 44 22253 0 S18
port 57 nsew
rlabel polycont 0 23508 0 23508 0 G18
port 58 nsew
rlabel ndiffc -44 24871 -44 24871 0 D19
port 59 nsew
rlabel ndiffc 44 24871 44 24871 0 S19
port 60 nsew
rlabel polycont 0 26126 0 26126 0 G19
port 61 nsew
<< properties >>
string FIXED_BBOX -158 -26228 158 26228
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12.0 l 0.15 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1 ad 3.48 as 3.48 pd 24.58 ps 24.58 nrd 0.0241666666666667 nrs 0.0241666666666667 sa 0 sb 0 sd 0 mult 20
<< end >>
