# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhvtop
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhvtop ;
  ORIGIN  0.000000  0.025000 ;
  SIZE  21.75000 BY  23.32000 ;
  PIN C0
    ANTENNAGATEAREA  320.0000 ;
    PORT
      LAYER met4 ;
        RECT  0.300000  0.140000  0.630000 23.220000 ;
        RECT  1.595000  0.865000  1.895000  5.665000 ;
        RECT  1.595000  5.665000  9.745000  5.995000 ;
        RECT  1.595000  5.995000  1.895000 10.795000 ;
        RECT  1.595000 12.405000  1.895000 17.205000 ;
        RECT  1.595000 17.205000  9.745000 17.535000 ;
        RECT  1.595000 17.535000  1.895000 22.335000 ;
        RECT  2.795000  0.865000  3.095000  5.665000 ;
        RECT  2.795000  5.995000  3.095000 10.795000 ;
        RECT  2.795000 12.405000  3.095000 17.205000 ;
        RECT  2.795000 17.535000  3.095000 22.335000 ;
        RECT  3.995000  0.865000  4.295000  5.665000 ;
        RECT  3.995000  5.995000  4.295000 10.795000 ;
        RECT  3.995000 12.405000  4.295000 17.205000 ;
        RECT  3.995000 17.535000  4.295000 22.335000 ;
        RECT  5.310000  0.865000  5.835000  5.665000 ;
        RECT  5.310000  5.995000  5.835000 10.795000 ;
        RECT  5.310000 12.405000  5.835000 17.205000 ;
        RECT  5.310000 17.535000  5.835000 22.335000 ;
        RECT  7.045000  0.865000  7.345000  5.665000 ;
        RECT  7.045000  5.995000  7.345000 10.795000 ;
        RECT  7.045000 12.405000  7.345000 17.205000 ;
        RECT  7.045000 17.535000  7.345000 22.335000 ;
        RECT  8.245000  0.865000  8.545000  5.665000 ;
        RECT  8.245000  5.995000  8.545000 10.795000 ;
        RECT  8.245000 12.405000  8.545000 17.205000 ;
        RECT  8.245000 17.535000  8.545000 22.335000 ;
        RECT  9.445000  0.865000  9.745000  5.665000 ;
        RECT  9.445000  5.995000  9.745000 10.795000 ;
        RECT  9.445000 12.405000  9.745000 17.205000 ;
        RECT  9.445000 17.535000  9.745000 22.335000 ;
        RECT 10.710000  0.140000 11.040000 23.220000 ;
        RECT 12.005000  0.865000 12.305000  5.665000 ;
        RECT 12.005000  5.665000 20.155000  5.995000 ;
        RECT 12.005000  5.995000 12.305000 10.795000 ;
        RECT 12.005000 12.405000 12.305000 17.205000 ;
        RECT 12.005000 17.205000 20.155000 17.535000 ;
        RECT 12.005000 17.535000 12.305000 22.335000 ;
        RECT 13.205000  0.865000 13.505000  5.665000 ;
        RECT 13.205000  5.995000 13.505000 10.795000 ;
        RECT 13.205000 12.405000 13.505000 17.205000 ;
        RECT 13.205000 17.535000 13.505000 22.335000 ;
        RECT 14.405000  0.865000 14.705000  5.665000 ;
        RECT 14.405000  5.995000 14.705000 10.795000 ;
        RECT 14.405000 12.405000 14.705000 17.205000 ;
        RECT 14.405000 17.535000 14.705000 22.335000 ;
        RECT 15.720000  0.865000 16.245000  5.665000 ;
        RECT 15.720000  5.995000 16.245000 10.795000 ;
        RECT 15.720000 12.405000 16.245000 17.205000 ;
        RECT 15.720000 17.535000 16.245000 22.335000 ;
        RECT 17.455000  0.865000 17.755000  5.665000 ;
        RECT 17.455000  5.995000 17.755000 10.795000 ;
        RECT 17.455000 12.405000 17.755000 17.205000 ;
        RECT 17.455000 17.535000 17.755000 22.335000 ;
        RECT 18.655000  0.865000 18.955000  5.665000 ;
        RECT 18.655000  5.995000 18.955000 10.795000 ;
        RECT 18.655000 12.405000 18.955000 17.205000 ;
        RECT 18.655000 17.535000 18.955000 22.335000 ;
        RECT 19.855000  0.865000 20.155000  5.665000 ;
        RECT 19.855000  5.995000 20.155000 10.795000 ;
        RECT 19.855000 12.405000 20.155000 17.205000 ;
        RECT 19.855000 17.535000 20.155000 22.335000 ;
        RECT 21.120000  0.140000 21.450000 23.220000 ;
    END
  END C0
  PIN M5
    PORT
      LAYER met5 ;
        RECT 0.000000 0.065000 21.750000 23.295000 ;
    END
  END M5
  PIN SUB
    ANTENNADIFFAREA  107.799995 ;
    PORT
      LAYER met4 ;
        RECT  0.965000  0.235000 10.375000  0.565000 ;
        RECT  0.965000  0.565000  1.295000 11.095000 ;
        RECT  0.965000 11.095000 10.375000 11.395000 ;
        RECT  0.965000 11.395000 10.045000 11.425000 ;
        RECT  0.965000 11.775000 10.375000 12.105000 ;
        RECT  0.965000 12.105000  1.295000 22.635000 ;
        RECT  0.965000 22.635000 10.375000 22.935000 ;
        RECT  0.965000 22.935000 10.045000 22.965000 ;
        RECT  2.195000  0.565000  2.495000  5.365000 ;
        RECT  2.195000  6.295000  2.495000 11.095000 ;
        RECT  2.195000 12.105000  2.495000 16.905000 ;
        RECT  2.195000 17.835000  2.495000 22.635000 ;
        RECT  3.395000  0.565000  3.695000  5.365000 ;
        RECT  3.395000  6.295000  3.695000 11.095000 ;
        RECT  3.395000 12.105000  3.695000 16.905000 ;
        RECT  3.395000 17.835000  3.695000 22.635000 ;
        RECT  4.595000  0.565000  5.010000  5.365000 ;
        RECT  4.595000  6.295000  5.010000 11.095000 ;
        RECT  4.595000 12.105000  5.010000 16.905000 ;
        RECT  4.595000 17.835000  5.010000 22.635000 ;
        RECT  6.135000  0.565000  6.745000  5.365000 ;
        RECT  6.135000  6.295000  6.745000 11.095000 ;
        RECT  6.135000 12.105000  6.745000 16.905000 ;
        RECT  6.135000 17.835000  6.745000 22.635000 ;
        RECT  7.645000  0.565000  7.945000  5.365000 ;
        RECT  7.645000  6.295000  7.945000 11.095000 ;
        RECT  7.645000 12.105000  7.945000 16.905000 ;
        RECT  7.645000 17.835000  7.945000 22.635000 ;
        RECT  8.845000  0.565000  9.145000  5.365000 ;
        RECT  8.845000  6.295000  9.145000 11.095000 ;
        RECT  8.845000 12.105000  9.145000 16.905000 ;
        RECT  8.845000 17.835000  9.145000 22.635000 ;
        RECT 10.045000  0.565000 10.375000 11.095000 ;
        RECT 10.045000 12.105000 10.375000 22.635000 ;
        RECT 11.375000  0.235000 20.785000  0.565000 ;
        RECT 11.375000  0.565000 11.705000 11.095000 ;
        RECT 11.375000 11.095000 20.785000 11.395000 ;
        RECT 11.375000 11.395000 20.455000 11.425000 ;
        RECT 11.375000 11.775000 20.785000 12.105000 ;
        RECT 11.375000 12.105000 11.705000 22.635000 ;
        RECT 11.375000 22.635000 20.785000 22.935000 ;
        RECT 11.375000 22.935000 20.455000 22.965000 ;
        RECT 12.605000  0.565000 12.905000  5.365000 ;
        RECT 12.605000  6.295000 12.905000 11.095000 ;
        RECT 12.605000 12.105000 12.905000 16.905000 ;
        RECT 12.605000 17.835000 12.905000 22.635000 ;
        RECT 13.805000  0.565000 14.105000  5.365000 ;
        RECT 13.805000  6.295000 14.105000 11.095000 ;
        RECT 13.805000 12.105000 14.105000 16.905000 ;
        RECT 13.805000 17.835000 14.105000 22.635000 ;
        RECT 15.005000  0.565000 15.420000  5.365000 ;
        RECT 15.005000  6.295000 15.420000 11.095000 ;
        RECT 15.005000 12.105000 15.420000 16.905000 ;
        RECT 15.005000 17.835000 15.420000 22.635000 ;
        RECT 16.545000  0.565000 17.155000  5.365000 ;
        RECT 16.545000  6.295000 17.155000 11.095000 ;
        RECT 16.545000 12.105000 17.155000 16.905000 ;
        RECT 16.545000 17.835000 17.155000 22.635000 ;
        RECT 18.055000  0.565000 18.355000  5.365000 ;
        RECT 18.055000  6.295000 18.355000 11.095000 ;
        RECT 18.055000 12.105000 18.355000 16.905000 ;
        RECT 18.055000 17.835000 18.355000 22.635000 ;
        RECT 19.255000  0.565000 19.555000  5.365000 ;
        RECT 19.255000  6.295000 19.555000 11.095000 ;
        RECT 19.255000 12.105000 19.555000 16.905000 ;
        RECT 19.255000 17.835000 19.555000 22.635000 ;
        RECT 20.455000  0.565000 20.785000 11.095000 ;
        RECT 20.455000 12.105000 20.785000 22.635000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT  0.465000  0.890000 21.285000  1.690000 ;
      RECT  0.465000  1.690000  1.175000 10.000000 ;
      RECT  0.465000 10.000000 21.285000 10.800000 ;
      RECT  0.465000 12.430000 21.285000 13.230000 ;
      RECT  0.465000 13.230000  1.175000 21.540000 ;
      RECT  0.465000 21.540000 21.285000 22.340000 ;
      RECT  1.355000  0.355000  9.980000  0.400000 ;
      RECT  1.355000  0.400000  9.985000  0.570000 ;
      RECT  1.355000  0.570000  9.980000  0.615000 ;
      RECT  1.355000 11.205000  9.980000 11.250000 ;
      RECT  1.355000 11.250000  9.985000 11.420000 ;
      RECT  1.355000 11.420000  9.980000 11.465000 ;
      RECT  1.355000 11.895000  9.980000 11.940000 ;
      RECT  1.355000 11.940000  9.985000 12.110000 ;
      RECT  1.355000 12.110000  9.980000 12.155000 ;
      RECT  1.355000 22.745000  9.980000 22.790000 ;
      RECT  1.355000 22.790000  9.985000 22.960000 ;
      RECT  1.355000 22.960000  9.980000 23.005000 ;
      RECT  1.450000  1.860000  1.620000  5.530000 ;
      RECT  1.450000  5.530000  5.260000  6.160000 ;
      RECT  1.450000  6.160000  1.620000  9.830000 ;
      RECT  1.450000 13.400000  1.620000 17.070000 ;
      RECT  1.450000 17.070000  5.260000 17.700000 ;
      RECT  1.450000 17.700000  1.620000 21.370000 ;
      RECT  1.800000  1.690000  1.970000  5.360000 ;
      RECT  1.800000  6.330000  1.970000 10.000000 ;
      RECT  1.800000 13.230000  1.970000 16.900000 ;
      RECT  1.800000 17.870000  1.970000 21.540000 ;
      RECT  2.150000  1.860000  2.320000  5.530000 ;
      RECT  2.150000  6.160000  2.320000  9.830000 ;
      RECT  2.150000 13.400000  2.320000 17.070000 ;
      RECT  2.150000 17.700000  2.320000 21.370000 ;
      RECT  2.500000  1.690000  2.670000  5.360000 ;
      RECT  2.500000  6.330000  2.670000 10.000000 ;
      RECT  2.500000 13.230000  2.670000 16.900000 ;
      RECT  2.500000 17.870000  2.670000 21.540000 ;
      RECT  2.850000  1.860000  3.020000  5.530000 ;
      RECT  2.850000  6.160000  3.020000  9.830000 ;
      RECT  2.850000 13.400000  3.020000 17.070000 ;
      RECT  2.850000 17.700000  3.020000 21.370000 ;
      RECT  3.200000  1.690000  3.370000  5.360000 ;
      RECT  3.200000  6.330000  3.370000 10.000000 ;
      RECT  3.200000 13.230000  3.370000 16.900000 ;
      RECT  3.200000 17.870000  3.370000 21.540000 ;
      RECT  3.550000  1.860000  3.720000  5.530000 ;
      RECT  3.550000  6.160000  3.720000  9.830000 ;
      RECT  3.550000 13.400000  3.720000 17.070000 ;
      RECT  3.550000 17.700000  3.720000 21.370000 ;
      RECT  3.900000  1.690000  4.070000  5.360000 ;
      RECT  3.900000  6.330000  4.070000 10.000000 ;
      RECT  3.900000 13.230000  4.070000 16.900000 ;
      RECT  3.900000 17.870000  4.070000 21.540000 ;
      RECT  4.250000  1.860000  4.420000  5.530000 ;
      RECT  4.250000  6.160000  4.420000  9.830000 ;
      RECT  4.250000 13.400000  4.420000 17.070000 ;
      RECT  4.250000 17.700000  4.420000 21.370000 ;
      RECT  4.600000  1.690000  4.770000  5.360000 ;
      RECT  4.600000  6.330000  4.770000 10.000000 ;
      RECT  4.600000 13.230000  4.770000 16.900000 ;
      RECT  4.600000 17.870000  4.770000 21.540000 ;
      RECT  4.950000  1.860000  5.120000  5.530000 ;
      RECT  4.950000  6.160000  5.120000  9.830000 ;
      RECT  4.950000 13.400000  5.120000 17.070000 ;
      RECT  4.950000 17.700000  5.120000 21.370000 ;
      RECT  5.300000  1.690000  6.040000  5.350000 ;
      RECT  5.300000  6.340000  5.900000  6.345000 ;
      RECT  5.300000  6.345000  6.040000 10.000000 ;
      RECT  5.300000 13.230000  6.040000 16.890000 ;
      RECT  5.300000 17.880000  5.900000 17.885000 ;
      RECT  5.300000 17.885000  6.040000 21.540000 ;
      RECT  5.440000  5.350000  5.900000  6.340000 ;
      RECT  5.440000 16.890000  5.900000 17.880000 ;
      RECT  6.080000  5.530000  9.890000  6.160000 ;
      RECT  6.080000 17.070000  9.890000 17.700000 ;
      RECT  6.220000  1.860000  6.390000  5.530000 ;
      RECT  6.220000  6.160000  6.390000  9.830000 ;
      RECT  6.220000 13.400000  6.390000 17.070000 ;
      RECT  6.220000 17.700000  6.390000 21.370000 ;
      RECT  6.570000  1.690000  6.740000  5.360000 ;
      RECT  6.570000  6.330000  6.740000 10.000000 ;
      RECT  6.570000 13.230000  6.740000 16.900000 ;
      RECT  6.570000 17.870000  6.740000 21.540000 ;
      RECT  6.920000  1.860000  7.090000  5.530000 ;
      RECT  6.920000  6.160000  7.090000  9.830000 ;
      RECT  6.920000 13.400000  7.090000 17.070000 ;
      RECT  6.920000 17.700000  7.090000 21.370000 ;
      RECT  7.270000  1.690000  7.440000  5.360000 ;
      RECT  7.270000  6.330000  7.440000 10.000000 ;
      RECT  7.270000 13.230000  7.440000 16.900000 ;
      RECT  7.270000 17.870000  7.440000 21.540000 ;
      RECT  7.620000  1.860000  7.790000  5.530000 ;
      RECT  7.620000  6.160000  7.790000  9.830000 ;
      RECT  7.620000 13.400000  7.790000 17.070000 ;
      RECT  7.620000 17.700000  7.790000 21.370000 ;
      RECT  7.970000  1.690000  8.140000  5.360000 ;
      RECT  7.970000  6.330000  8.140000 10.000000 ;
      RECT  7.970000 13.230000  8.140000 16.900000 ;
      RECT  7.970000 17.870000  8.140000 21.540000 ;
      RECT  8.320000  1.860000  8.490000  5.530000 ;
      RECT  8.320000  6.160000  8.490000  9.830000 ;
      RECT  8.320000 13.400000  8.490000 17.070000 ;
      RECT  8.320000 17.700000  8.490000 21.370000 ;
      RECT  8.670000  1.690000  8.840000  5.360000 ;
      RECT  8.670000  6.330000  8.840000 10.000000 ;
      RECT  8.670000 13.230000  8.840000 16.900000 ;
      RECT  8.670000 17.870000  8.840000 21.540000 ;
      RECT  9.020000  1.860000  9.190000  5.530000 ;
      RECT  9.020000  6.160000  9.190000  9.830000 ;
      RECT  9.020000 13.400000  9.190000 17.070000 ;
      RECT  9.020000 17.700000  9.190000 21.370000 ;
      RECT  9.370000  1.690000  9.540000  5.360000 ;
      RECT  9.370000  6.330000  9.540000 10.000000 ;
      RECT  9.370000 13.230000  9.540000 16.900000 ;
      RECT  9.370000 17.870000  9.540000 21.540000 ;
      RECT  9.720000  1.860000  9.890000  5.530000 ;
      RECT  9.720000  6.160000  9.890000  9.830000 ;
      RECT  9.720000 13.400000  9.890000 17.070000 ;
      RECT  9.720000 17.700000  9.890000 21.370000 ;
      RECT 10.165000  1.690000 11.585000 10.000000 ;
      RECT 10.165000 13.230000 11.585000 21.540000 ;
      RECT 11.765000  0.355000 20.390000  0.400000 ;
      RECT 11.765000  0.400000 20.395000  0.570000 ;
      RECT 11.765000  0.570000 20.390000  0.615000 ;
      RECT 11.765000 11.205000 20.390000 11.250000 ;
      RECT 11.765000 11.250000 20.395000 11.420000 ;
      RECT 11.765000 11.420000 20.390000 11.465000 ;
      RECT 11.765000 11.895000 20.390000 11.940000 ;
      RECT 11.765000 11.940000 20.395000 12.110000 ;
      RECT 11.765000 12.110000 20.390000 12.155000 ;
      RECT 11.765000 22.745000 20.390000 22.790000 ;
      RECT 11.765000 22.790000 20.395000 22.960000 ;
      RECT 11.765000 22.960000 20.390000 23.005000 ;
      RECT 11.860000  1.860000 12.030000  5.530000 ;
      RECT 11.860000  5.530000 15.670000  6.160000 ;
      RECT 11.860000  6.160000 12.030000  9.830000 ;
      RECT 11.860000 13.400000 12.030000 17.070000 ;
      RECT 11.860000 17.070000 15.670000 17.700000 ;
      RECT 11.860000 17.700000 12.030000 21.370000 ;
      RECT 12.210000  1.690000 12.380000  5.360000 ;
      RECT 12.210000  6.330000 12.380000 10.000000 ;
      RECT 12.210000 13.230000 12.380000 16.900000 ;
      RECT 12.210000 17.870000 12.380000 21.540000 ;
      RECT 12.560000  1.860000 12.730000  5.530000 ;
      RECT 12.560000  6.160000 12.730000  9.830000 ;
      RECT 12.560000 13.400000 12.730000 17.070000 ;
      RECT 12.560000 17.700000 12.730000 21.370000 ;
      RECT 12.910000  1.690000 13.080000  5.360000 ;
      RECT 12.910000  6.330000 13.080000 10.000000 ;
      RECT 12.910000 13.230000 13.080000 16.900000 ;
      RECT 12.910000 17.870000 13.080000 21.540000 ;
      RECT 13.260000  1.860000 13.430000  5.530000 ;
      RECT 13.260000  6.160000 13.430000  9.830000 ;
      RECT 13.260000 13.400000 13.430000 17.070000 ;
      RECT 13.260000 17.700000 13.430000 21.370000 ;
      RECT 13.610000  1.690000 13.780000  5.360000 ;
      RECT 13.610000  6.330000 13.780000 10.000000 ;
      RECT 13.610000 13.230000 13.780000 16.900000 ;
      RECT 13.610000 17.870000 13.780000 21.540000 ;
      RECT 13.960000  1.860000 14.130000  5.530000 ;
      RECT 13.960000  6.160000 14.130000  9.830000 ;
      RECT 13.960000 13.400000 14.130000 17.070000 ;
      RECT 13.960000 17.700000 14.130000 21.370000 ;
      RECT 14.310000  1.690000 14.480000  5.360000 ;
      RECT 14.310000  6.330000 14.480000 10.000000 ;
      RECT 14.310000 13.230000 14.480000 16.900000 ;
      RECT 14.310000 17.870000 14.480000 21.540000 ;
      RECT 14.660000  1.860000 14.830000  5.530000 ;
      RECT 14.660000  6.160000 14.830000  9.830000 ;
      RECT 14.660000 13.400000 14.830000 17.070000 ;
      RECT 14.660000 17.700000 14.830000 21.370000 ;
      RECT 15.010000  1.690000 15.180000  5.360000 ;
      RECT 15.010000  6.330000 15.180000 10.000000 ;
      RECT 15.010000 13.230000 15.180000 16.900000 ;
      RECT 15.010000 17.870000 15.180000 21.540000 ;
      RECT 15.360000  1.860000 15.530000  5.530000 ;
      RECT 15.360000  6.160000 15.530000  9.830000 ;
      RECT 15.360000 13.400000 15.530000 17.070000 ;
      RECT 15.360000 17.700000 15.530000 21.370000 ;
      RECT 15.710000  1.690000 16.450000  5.350000 ;
      RECT 15.710000  6.340000 16.310000  6.345000 ;
      RECT 15.710000  6.345000 16.450000 10.000000 ;
      RECT 15.710000 13.230000 16.450000 16.890000 ;
      RECT 15.710000 17.880000 16.310000 17.885000 ;
      RECT 15.710000 17.885000 16.450000 21.540000 ;
      RECT 15.850000  5.350000 16.310000  6.340000 ;
      RECT 15.850000 16.890000 16.310000 17.880000 ;
      RECT 16.490000  5.530000 20.300000  6.160000 ;
      RECT 16.490000 17.070000 20.300000 17.700000 ;
      RECT 16.630000  1.860000 16.800000  5.530000 ;
      RECT 16.630000  6.160000 16.800000  9.830000 ;
      RECT 16.630000 13.400000 16.800000 17.070000 ;
      RECT 16.630000 17.700000 16.800000 21.370000 ;
      RECT 16.980000  1.690000 17.150000  5.360000 ;
      RECT 16.980000  6.330000 17.150000 10.000000 ;
      RECT 16.980000 13.230000 17.150000 16.900000 ;
      RECT 16.980000 17.870000 17.150000 21.540000 ;
      RECT 17.330000  1.860000 17.500000  5.530000 ;
      RECT 17.330000  6.160000 17.500000  9.830000 ;
      RECT 17.330000 13.400000 17.500000 17.070000 ;
      RECT 17.330000 17.700000 17.500000 21.370000 ;
      RECT 17.680000  1.690000 17.850000  5.360000 ;
      RECT 17.680000  6.330000 17.850000 10.000000 ;
      RECT 17.680000 13.230000 17.850000 16.900000 ;
      RECT 17.680000 17.870000 17.850000 21.540000 ;
      RECT 18.030000  1.860000 18.200000  5.530000 ;
      RECT 18.030000  6.160000 18.200000  9.830000 ;
      RECT 18.030000 13.400000 18.200000 17.070000 ;
      RECT 18.030000 17.700000 18.200000 21.370000 ;
      RECT 18.380000  1.690000 18.550000  5.360000 ;
      RECT 18.380000  6.330000 18.550000 10.000000 ;
      RECT 18.380000 13.230000 18.550000 16.900000 ;
      RECT 18.380000 17.870000 18.550000 21.540000 ;
      RECT 18.730000  1.860000 18.900000  5.530000 ;
      RECT 18.730000  6.160000 18.900000  9.830000 ;
      RECT 18.730000 13.400000 18.900000 17.070000 ;
      RECT 18.730000 17.700000 18.900000 21.370000 ;
      RECT 19.080000  1.690000 19.250000  5.360000 ;
      RECT 19.080000  6.330000 19.250000 10.000000 ;
      RECT 19.080000 13.230000 19.250000 16.900000 ;
      RECT 19.080000 17.870000 19.250000 21.540000 ;
      RECT 19.430000  1.860000 19.600000  5.530000 ;
      RECT 19.430000  6.160000 19.600000  9.830000 ;
      RECT 19.430000 13.400000 19.600000 17.070000 ;
      RECT 19.430000 17.700000 19.600000 21.370000 ;
      RECT 19.780000  1.690000 19.950000  5.360000 ;
      RECT 19.780000  6.330000 19.950000 10.000000 ;
      RECT 19.780000 13.230000 19.950000 16.900000 ;
      RECT 19.780000 17.870000 19.950000 21.540000 ;
      RECT 20.130000  1.860000 20.300000  5.530000 ;
      RECT 20.130000  6.160000 20.300000  9.830000 ;
      RECT 20.130000 13.400000 20.300000 17.070000 ;
      RECT 20.130000 17.700000 20.300000 21.370000 ;
      RECT 20.575000  1.690000 21.285000 10.000000 ;
      RECT 20.575000 13.230000 21.285000 21.540000 ;
    LAYER mcon ;
      RECT  0.645000  1.080000  1.175000 10.610000 ;
      RECT  0.645000 12.620000  1.175000 22.150000 ;
      RECT  1.415000  0.400000  1.585000  0.570000 ;
      RECT  1.415000 11.250000  1.585000 11.420000 ;
      RECT  1.415000 11.940000  1.585000 12.110000 ;
      RECT  1.415000 22.790000  1.585000 22.960000 ;
      RECT  1.595000  1.470000  1.765000  1.640000 ;
      RECT  1.595000 10.050000  1.765000 10.220000 ;
      RECT  1.595000 13.010000  1.765000 13.180000 ;
      RECT  1.595000 21.590000  1.765000 21.760000 ;
      RECT  1.720000  5.580000  5.130000  6.110000 ;
      RECT  1.720000 17.120000  5.130000 17.650000 ;
      RECT  1.775000  0.400000  1.945000  0.570000 ;
      RECT  1.775000 11.250000  1.945000 11.420000 ;
      RECT  1.775000 11.940000  1.945000 12.110000 ;
      RECT  1.775000 22.790000  1.945000 22.960000 ;
      RECT  1.955000  1.470000  2.125000  1.640000 ;
      RECT  1.955000 10.050000  2.125000 10.220000 ;
      RECT  1.955000 13.010000  2.125000 13.180000 ;
      RECT  1.955000 21.590000  2.125000 21.760000 ;
      RECT  2.135000  0.400000  2.305000  0.570000 ;
      RECT  2.135000 11.250000  2.305000 11.420000 ;
      RECT  2.135000 11.940000  2.305000 12.110000 ;
      RECT  2.135000 22.790000  2.305000 22.960000 ;
      RECT  2.315000  1.470000  2.485000  1.640000 ;
      RECT  2.315000 10.050000  2.485000 10.220000 ;
      RECT  2.315000 13.010000  2.485000 13.180000 ;
      RECT  2.315000 21.590000  2.485000 21.760000 ;
      RECT  2.495000  0.400000  2.665000  0.570000 ;
      RECT  2.495000 11.250000  2.665000 11.420000 ;
      RECT  2.495000 11.940000  2.665000 12.110000 ;
      RECT  2.495000 22.790000  2.665000 22.960000 ;
      RECT  2.675000  1.470000  2.845000  1.640000 ;
      RECT  2.675000 10.050000  2.845000 10.220000 ;
      RECT  2.675000 13.010000  2.845000 13.180000 ;
      RECT  2.675000 21.590000  2.845000 21.760000 ;
      RECT  2.855000  0.400000  3.025000  0.570000 ;
      RECT  2.855000 11.250000  3.025000 11.420000 ;
      RECT  2.855000 11.940000  3.025000 12.110000 ;
      RECT  2.855000 22.790000  3.025000 22.960000 ;
      RECT  3.035000  1.470000  3.205000  1.640000 ;
      RECT  3.035000 10.050000  3.205000 10.220000 ;
      RECT  3.035000 13.010000  3.205000 13.180000 ;
      RECT  3.035000 21.590000  3.205000 21.760000 ;
      RECT  3.215000  0.400000  3.385000  0.570000 ;
      RECT  3.215000 11.250000  3.385000 11.420000 ;
      RECT  3.215000 11.940000  3.385000 12.110000 ;
      RECT  3.215000 22.790000  3.385000 22.960000 ;
      RECT  3.395000  1.470000  3.565000  1.640000 ;
      RECT  3.395000 10.050000  3.565000 10.220000 ;
      RECT  3.395000 13.010000  3.565000 13.180000 ;
      RECT  3.395000 21.590000  3.565000 21.760000 ;
      RECT  3.575000  0.400000  3.745000  0.570000 ;
      RECT  3.575000 11.250000  3.745000 11.420000 ;
      RECT  3.575000 11.940000  3.745000 12.110000 ;
      RECT  3.575000 22.790000  3.745000 22.960000 ;
      RECT  3.755000  1.470000  3.925000  1.640000 ;
      RECT  3.755000 10.050000  3.925000 10.220000 ;
      RECT  3.755000 13.010000  3.925000 13.180000 ;
      RECT  3.755000 21.590000  3.925000 21.760000 ;
      RECT  3.935000  0.400000  4.105000  0.570000 ;
      RECT  3.935000 11.250000  4.105000 11.420000 ;
      RECT  3.935000 11.940000  4.105000 12.110000 ;
      RECT  3.935000 22.790000  4.105000 22.960000 ;
      RECT  4.115000  1.470000  4.285000  1.640000 ;
      RECT  4.115000 10.050000  4.285000 10.220000 ;
      RECT  4.115000 13.010000  4.285000 13.180000 ;
      RECT  4.115000 21.590000  4.285000 21.760000 ;
      RECT  4.295000  0.400000  4.465000  0.570000 ;
      RECT  4.295000 11.250000  4.465000 11.420000 ;
      RECT  4.295000 11.940000  4.465000 12.110000 ;
      RECT  4.295000 22.790000  4.465000 22.960000 ;
      RECT  4.475000  1.470000  4.645000  1.640000 ;
      RECT  4.475000 10.050000  4.645000 10.220000 ;
      RECT  4.475000 13.010000  4.645000 13.180000 ;
      RECT  4.475000 21.590000  4.645000 21.760000 ;
      RECT  4.655000  0.400000  4.825000  0.570000 ;
      RECT  4.655000 11.250000  4.825000 11.420000 ;
      RECT  4.655000 11.940000  4.825000 12.110000 ;
      RECT  4.655000 22.790000  4.825000 22.960000 ;
      RECT  4.835000  1.470000  5.005000  1.640000 ;
      RECT  4.835000 10.050000  5.005000 10.220000 ;
      RECT  4.835000 13.010000  5.005000 13.180000 ;
      RECT  4.835000 21.590000  5.005000 21.760000 ;
      RECT  5.015000  0.400000  5.185000  0.570000 ;
      RECT  5.015000 11.250000  5.185000 11.420000 ;
      RECT  5.015000 11.940000  5.185000 12.110000 ;
      RECT  5.015000 22.790000  5.185000 22.960000 ;
      RECT  5.375000  0.400000  5.545000  0.570000 ;
      RECT  5.375000 11.250000  5.545000 11.420000 ;
      RECT  5.375000 11.940000  5.545000 12.110000 ;
      RECT  5.375000 22.790000  5.545000 22.960000 ;
      RECT  5.735000  0.400000  5.905000  0.570000 ;
      RECT  5.735000 11.250000  5.905000 11.420000 ;
      RECT  5.735000 11.940000  5.905000 12.110000 ;
      RECT  5.735000 22.790000  5.905000 22.960000 ;
      RECT  6.095000  0.400000  6.265000  0.570000 ;
      RECT  6.095000 11.250000  6.265000 11.420000 ;
      RECT  6.095000 11.940000  6.265000 12.110000 ;
      RECT  6.095000 22.790000  6.265000 22.960000 ;
      RECT  6.210000  5.580000  9.620000  6.110000 ;
      RECT  6.210000 17.120000  9.620000 17.650000 ;
      RECT  6.335000  1.470000  6.505000  1.640000 ;
      RECT  6.335000 10.050000  6.505000 10.220000 ;
      RECT  6.335000 13.010000  6.505000 13.180000 ;
      RECT  6.335000 21.590000  6.505000 21.760000 ;
      RECT  6.455000  0.400000  6.625000  0.570000 ;
      RECT  6.455000 11.250000  6.625000 11.420000 ;
      RECT  6.455000 11.940000  6.625000 12.110000 ;
      RECT  6.455000 22.790000  6.625000 22.960000 ;
      RECT  6.695000  1.470000  6.865000  1.640000 ;
      RECT  6.695000 10.050000  6.865000 10.220000 ;
      RECT  6.695000 13.010000  6.865000 13.180000 ;
      RECT  6.695000 21.590000  6.865000 21.760000 ;
      RECT  6.815000  0.400000  6.985000  0.570000 ;
      RECT  6.815000 11.250000  6.985000 11.420000 ;
      RECT  6.815000 11.940000  6.985000 12.110000 ;
      RECT  6.815000 22.790000  6.985000 22.960000 ;
      RECT  7.055000  1.470000  7.225000  1.640000 ;
      RECT  7.055000 10.050000  7.225000 10.220000 ;
      RECT  7.055000 13.010000  7.225000 13.180000 ;
      RECT  7.055000 21.590000  7.225000 21.760000 ;
      RECT  7.175000  0.400000  7.345000  0.570000 ;
      RECT  7.175000 11.250000  7.345000 11.420000 ;
      RECT  7.175000 11.940000  7.345000 12.110000 ;
      RECT  7.175000 22.790000  7.345000 22.960000 ;
      RECT  7.415000  1.470000  7.585000  1.640000 ;
      RECT  7.415000 10.050000  7.585000 10.220000 ;
      RECT  7.415000 13.010000  7.585000 13.180000 ;
      RECT  7.415000 21.590000  7.585000 21.760000 ;
      RECT  7.535000  0.400000  7.705000  0.570000 ;
      RECT  7.535000 11.250000  7.705000 11.420000 ;
      RECT  7.535000 11.940000  7.705000 12.110000 ;
      RECT  7.535000 22.790000  7.705000 22.960000 ;
      RECT  7.775000  1.470000  7.945000  1.640000 ;
      RECT  7.775000 10.050000  7.945000 10.220000 ;
      RECT  7.775000 13.010000  7.945000 13.180000 ;
      RECT  7.775000 21.590000  7.945000 21.760000 ;
      RECT  7.895000  0.400000  8.065000  0.570000 ;
      RECT  7.895000 11.250000  8.065000 11.420000 ;
      RECT  7.895000 11.940000  8.065000 12.110000 ;
      RECT  7.895000 22.790000  8.065000 22.960000 ;
      RECT  8.135000  1.470000  8.305000  1.640000 ;
      RECT  8.135000 10.050000  8.305000 10.220000 ;
      RECT  8.135000 13.010000  8.305000 13.180000 ;
      RECT  8.135000 21.590000  8.305000 21.760000 ;
      RECT  8.255000  0.400000  8.425000  0.570000 ;
      RECT  8.255000 11.250000  8.425000 11.420000 ;
      RECT  8.255000 11.940000  8.425000 12.110000 ;
      RECT  8.255000 22.790000  8.425000 22.960000 ;
      RECT  8.495000  1.470000  8.665000  1.640000 ;
      RECT  8.495000 10.050000  8.665000 10.220000 ;
      RECT  8.495000 13.010000  8.665000 13.180000 ;
      RECT  8.495000 21.590000  8.665000 21.760000 ;
      RECT  8.615000  0.400000  8.785000  0.570000 ;
      RECT  8.615000 11.250000  8.785000 11.420000 ;
      RECT  8.615000 11.940000  8.785000 12.110000 ;
      RECT  8.615000 22.790000  8.785000 22.960000 ;
      RECT  8.855000  1.470000  9.025000  1.640000 ;
      RECT  8.855000 10.050000  9.025000 10.220000 ;
      RECT  8.855000 13.010000  9.025000 13.180000 ;
      RECT  8.855000 21.590000  9.025000 21.760000 ;
      RECT  8.975000  0.400000  9.145000  0.570000 ;
      RECT  8.975000 11.250000  9.145000 11.420000 ;
      RECT  8.975000 11.940000  9.145000 12.110000 ;
      RECT  8.975000 22.790000  9.145000 22.960000 ;
      RECT  9.215000  1.470000  9.385000  1.640000 ;
      RECT  9.215000 10.050000  9.385000 10.220000 ;
      RECT  9.215000 13.010000  9.385000 13.180000 ;
      RECT  9.215000 21.590000  9.385000 21.760000 ;
      RECT  9.335000  0.400000  9.505000  0.570000 ;
      RECT  9.335000 11.250000  9.505000 11.420000 ;
      RECT  9.335000 11.940000  9.505000 12.110000 ;
      RECT  9.335000 22.790000  9.505000 22.960000 ;
      RECT  9.575000  1.470000  9.745000  1.640000 ;
      RECT  9.575000 10.050000  9.745000 10.220000 ;
      RECT  9.575000 13.010000  9.745000 13.180000 ;
      RECT  9.575000 21.590000  9.745000 21.760000 ;
      RECT  9.695000  0.400000  9.865000  0.570000 ;
      RECT  9.695000 11.250000  9.865000 11.420000 ;
      RECT  9.695000 11.940000  9.865000 12.110000 ;
      RECT  9.695000 22.790000  9.865000 22.960000 ;
      RECT 10.165000  1.080000 10.695000 10.610000 ;
      RECT 10.165000 12.620000 10.695000 22.150000 ;
      RECT 11.055000  1.080000 11.585000 10.610000 ;
      RECT 11.055000 12.620000 11.585000 22.150000 ;
      RECT 11.825000  0.400000 11.995000  0.570000 ;
      RECT 11.825000 11.250000 11.995000 11.420000 ;
      RECT 11.825000 11.940000 11.995000 12.110000 ;
      RECT 11.825000 22.790000 11.995000 22.960000 ;
      RECT 12.005000  1.470000 12.175000  1.640000 ;
      RECT 12.005000 10.050000 12.175000 10.220000 ;
      RECT 12.005000 13.010000 12.175000 13.180000 ;
      RECT 12.005000 21.590000 12.175000 21.760000 ;
      RECT 12.130000  5.580000 15.540000  6.110000 ;
      RECT 12.130000 17.120000 15.540000 17.650000 ;
      RECT 12.185000  0.400000 12.355000  0.570000 ;
      RECT 12.185000 11.250000 12.355000 11.420000 ;
      RECT 12.185000 11.940000 12.355000 12.110000 ;
      RECT 12.185000 22.790000 12.355000 22.960000 ;
      RECT 12.365000  1.470000 12.535000  1.640000 ;
      RECT 12.365000 10.050000 12.535000 10.220000 ;
      RECT 12.365000 13.010000 12.535000 13.180000 ;
      RECT 12.365000 21.590000 12.535000 21.760000 ;
      RECT 12.545000  0.400000 12.715000  0.570000 ;
      RECT 12.545000 11.250000 12.715000 11.420000 ;
      RECT 12.545000 11.940000 12.715000 12.110000 ;
      RECT 12.545000 22.790000 12.715000 22.960000 ;
      RECT 12.725000  1.470000 12.895000  1.640000 ;
      RECT 12.725000 10.050000 12.895000 10.220000 ;
      RECT 12.725000 13.010000 12.895000 13.180000 ;
      RECT 12.725000 21.590000 12.895000 21.760000 ;
      RECT 12.905000  0.400000 13.075000  0.570000 ;
      RECT 12.905000 11.250000 13.075000 11.420000 ;
      RECT 12.905000 11.940000 13.075000 12.110000 ;
      RECT 12.905000 22.790000 13.075000 22.960000 ;
      RECT 13.085000  1.470000 13.255000  1.640000 ;
      RECT 13.085000 10.050000 13.255000 10.220000 ;
      RECT 13.085000 13.010000 13.255000 13.180000 ;
      RECT 13.085000 21.590000 13.255000 21.760000 ;
      RECT 13.265000  0.400000 13.435000  0.570000 ;
      RECT 13.265000 11.250000 13.435000 11.420000 ;
      RECT 13.265000 11.940000 13.435000 12.110000 ;
      RECT 13.265000 22.790000 13.435000 22.960000 ;
      RECT 13.445000  1.470000 13.615000  1.640000 ;
      RECT 13.445000 10.050000 13.615000 10.220000 ;
      RECT 13.445000 13.010000 13.615000 13.180000 ;
      RECT 13.445000 21.590000 13.615000 21.760000 ;
      RECT 13.625000  0.400000 13.795000  0.570000 ;
      RECT 13.625000 11.250000 13.795000 11.420000 ;
      RECT 13.625000 11.940000 13.795000 12.110000 ;
      RECT 13.625000 22.790000 13.795000 22.960000 ;
      RECT 13.805000  1.470000 13.975000  1.640000 ;
      RECT 13.805000 10.050000 13.975000 10.220000 ;
      RECT 13.805000 13.010000 13.975000 13.180000 ;
      RECT 13.805000 21.590000 13.975000 21.760000 ;
      RECT 13.985000  0.400000 14.155000  0.570000 ;
      RECT 13.985000 11.250000 14.155000 11.420000 ;
      RECT 13.985000 11.940000 14.155000 12.110000 ;
      RECT 13.985000 22.790000 14.155000 22.960000 ;
      RECT 14.165000  1.470000 14.335000  1.640000 ;
      RECT 14.165000 10.050000 14.335000 10.220000 ;
      RECT 14.165000 13.010000 14.335000 13.180000 ;
      RECT 14.165000 21.590000 14.335000 21.760000 ;
      RECT 14.345000  0.400000 14.515000  0.570000 ;
      RECT 14.345000 11.250000 14.515000 11.420000 ;
      RECT 14.345000 11.940000 14.515000 12.110000 ;
      RECT 14.345000 22.790000 14.515000 22.960000 ;
      RECT 14.525000  1.470000 14.695000  1.640000 ;
      RECT 14.525000 10.050000 14.695000 10.220000 ;
      RECT 14.525000 13.010000 14.695000 13.180000 ;
      RECT 14.525000 21.590000 14.695000 21.760000 ;
      RECT 14.705000  0.400000 14.875000  0.570000 ;
      RECT 14.705000 11.250000 14.875000 11.420000 ;
      RECT 14.705000 11.940000 14.875000 12.110000 ;
      RECT 14.705000 22.790000 14.875000 22.960000 ;
      RECT 14.885000  1.470000 15.055000  1.640000 ;
      RECT 14.885000 10.050000 15.055000 10.220000 ;
      RECT 14.885000 13.010000 15.055000 13.180000 ;
      RECT 14.885000 21.590000 15.055000 21.760000 ;
      RECT 15.065000  0.400000 15.235000  0.570000 ;
      RECT 15.065000 11.250000 15.235000 11.420000 ;
      RECT 15.065000 11.940000 15.235000 12.110000 ;
      RECT 15.065000 22.790000 15.235000 22.960000 ;
      RECT 15.245000  1.470000 15.415000  1.640000 ;
      RECT 15.245000 10.050000 15.415000 10.220000 ;
      RECT 15.245000 13.010000 15.415000 13.180000 ;
      RECT 15.245000 21.590000 15.415000 21.760000 ;
      RECT 15.425000  0.400000 15.595000  0.570000 ;
      RECT 15.425000 11.250000 15.595000 11.420000 ;
      RECT 15.425000 11.940000 15.595000 12.110000 ;
      RECT 15.425000 22.790000 15.595000 22.960000 ;
      RECT 15.785000  0.400000 15.955000  0.570000 ;
      RECT 15.785000 11.250000 15.955000 11.420000 ;
      RECT 15.785000 11.940000 15.955000 12.110000 ;
      RECT 15.785000 22.790000 15.955000 22.960000 ;
      RECT 16.145000  0.400000 16.315000  0.570000 ;
      RECT 16.145000 11.250000 16.315000 11.420000 ;
      RECT 16.145000 11.940000 16.315000 12.110000 ;
      RECT 16.145000 22.790000 16.315000 22.960000 ;
      RECT 16.505000  0.400000 16.675000  0.570000 ;
      RECT 16.505000 11.250000 16.675000 11.420000 ;
      RECT 16.505000 11.940000 16.675000 12.110000 ;
      RECT 16.505000 22.790000 16.675000 22.960000 ;
      RECT 16.620000  5.580000 20.030000  6.110000 ;
      RECT 16.620000 17.120000 20.030000 17.650000 ;
      RECT 16.745000  1.470000 16.915000  1.640000 ;
      RECT 16.745000 10.050000 16.915000 10.220000 ;
      RECT 16.745000 13.010000 16.915000 13.180000 ;
      RECT 16.745000 21.590000 16.915000 21.760000 ;
      RECT 16.865000  0.400000 17.035000  0.570000 ;
      RECT 16.865000 11.250000 17.035000 11.420000 ;
      RECT 16.865000 11.940000 17.035000 12.110000 ;
      RECT 16.865000 22.790000 17.035000 22.960000 ;
      RECT 17.105000  1.470000 17.275000  1.640000 ;
      RECT 17.105000 10.050000 17.275000 10.220000 ;
      RECT 17.105000 13.010000 17.275000 13.180000 ;
      RECT 17.105000 21.590000 17.275000 21.760000 ;
      RECT 17.225000  0.400000 17.395000  0.570000 ;
      RECT 17.225000 11.250000 17.395000 11.420000 ;
      RECT 17.225000 11.940000 17.395000 12.110000 ;
      RECT 17.225000 22.790000 17.395000 22.960000 ;
      RECT 17.465000  1.470000 17.635000  1.640000 ;
      RECT 17.465000 10.050000 17.635000 10.220000 ;
      RECT 17.465000 13.010000 17.635000 13.180000 ;
      RECT 17.465000 21.590000 17.635000 21.760000 ;
      RECT 17.585000  0.400000 17.755000  0.570000 ;
      RECT 17.585000 11.250000 17.755000 11.420000 ;
      RECT 17.585000 11.940000 17.755000 12.110000 ;
      RECT 17.585000 22.790000 17.755000 22.960000 ;
      RECT 17.825000  1.470000 17.995000  1.640000 ;
      RECT 17.825000 10.050000 17.995000 10.220000 ;
      RECT 17.825000 13.010000 17.995000 13.180000 ;
      RECT 17.825000 21.590000 17.995000 21.760000 ;
      RECT 17.945000  0.400000 18.115000  0.570000 ;
      RECT 17.945000 11.250000 18.115000 11.420000 ;
      RECT 17.945000 11.940000 18.115000 12.110000 ;
      RECT 17.945000 22.790000 18.115000 22.960000 ;
      RECT 18.185000  1.470000 18.355000  1.640000 ;
      RECT 18.185000 10.050000 18.355000 10.220000 ;
      RECT 18.185000 13.010000 18.355000 13.180000 ;
      RECT 18.185000 21.590000 18.355000 21.760000 ;
      RECT 18.305000  0.400000 18.475000  0.570000 ;
      RECT 18.305000 11.250000 18.475000 11.420000 ;
      RECT 18.305000 11.940000 18.475000 12.110000 ;
      RECT 18.305000 22.790000 18.475000 22.960000 ;
      RECT 18.545000  1.470000 18.715000  1.640000 ;
      RECT 18.545000 10.050000 18.715000 10.220000 ;
      RECT 18.545000 13.010000 18.715000 13.180000 ;
      RECT 18.545000 21.590000 18.715000 21.760000 ;
      RECT 18.665000  0.400000 18.835000  0.570000 ;
      RECT 18.665000 11.250000 18.835000 11.420000 ;
      RECT 18.665000 11.940000 18.835000 12.110000 ;
      RECT 18.665000 22.790000 18.835000 22.960000 ;
      RECT 18.905000  1.470000 19.075000  1.640000 ;
      RECT 18.905000 10.050000 19.075000 10.220000 ;
      RECT 18.905000 13.010000 19.075000 13.180000 ;
      RECT 18.905000 21.590000 19.075000 21.760000 ;
      RECT 19.025000  0.400000 19.195000  0.570000 ;
      RECT 19.025000 11.250000 19.195000 11.420000 ;
      RECT 19.025000 11.940000 19.195000 12.110000 ;
      RECT 19.025000 22.790000 19.195000 22.960000 ;
      RECT 19.265000  1.470000 19.435000  1.640000 ;
      RECT 19.265000 10.050000 19.435000 10.220000 ;
      RECT 19.265000 13.010000 19.435000 13.180000 ;
      RECT 19.265000 21.590000 19.435000 21.760000 ;
      RECT 19.385000  0.400000 19.555000  0.570000 ;
      RECT 19.385000 11.250000 19.555000 11.420000 ;
      RECT 19.385000 11.940000 19.555000 12.110000 ;
      RECT 19.385000 22.790000 19.555000 22.960000 ;
      RECT 19.625000  1.470000 19.795000  1.640000 ;
      RECT 19.625000 10.050000 19.795000 10.220000 ;
      RECT 19.625000 13.010000 19.795000 13.180000 ;
      RECT 19.625000 21.590000 19.795000 21.760000 ;
      RECT 19.745000  0.400000 19.915000  0.570000 ;
      RECT 19.745000 11.250000 19.915000 11.420000 ;
      RECT 19.745000 11.940000 19.915000 12.110000 ;
      RECT 19.745000 22.790000 19.915000 22.960000 ;
      RECT 19.985000  1.470000 20.155000  1.640000 ;
      RECT 19.985000 10.050000 20.155000 10.220000 ;
      RECT 19.985000 13.010000 20.155000 13.180000 ;
      RECT 19.985000 21.590000 20.155000 21.760000 ;
      RECT 20.105000  0.400000 20.275000  0.570000 ;
      RECT 20.105000 11.250000 20.275000 11.420000 ;
      RECT 20.105000 11.940000 20.275000 12.110000 ;
      RECT 20.105000 22.790000 20.275000 22.960000 ;
      RECT 20.575000  1.080000 21.105000 10.610000 ;
      RECT 20.575000 12.620000 21.105000 22.150000 ;
    LAYER met1 ;
      RECT  0.465000  0.065000 21.285000  0.215000 ;
      RECT  0.465000  0.215000  1.215000  1.420000 ;
      RECT  0.465000  1.420000  5.120000  1.690000 ;
      RECT  0.465000  1.690000  1.310000  2.140000 ;
      RECT  0.465000  2.140000  5.120000  2.280000 ;
      RECT  0.465000  2.280000  1.310000  2.700000 ;
      RECT  0.465000  2.700000  5.120000  2.840000 ;
      RECT  0.465000  2.840000  1.310000  3.260000 ;
      RECT  0.465000  3.260000  5.120000  3.400000 ;
      RECT  0.465000  3.400000  1.310000  3.820000 ;
      RECT  0.465000  3.820000  5.120000  3.960000 ;
      RECT  0.465000  3.960000  1.310000  4.380000 ;
      RECT  0.465000  4.380000  5.120000  4.520000 ;
      RECT  0.465000  4.520000  1.310000  4.940000 ;
      RECT  0.465000  4.940000  5.120000  5.080000 ;
      RECT  0.465000  5.080000  1.310000  6.610000 ;
      RECT  0.465000  6.610000  5.120000  6.750000 ;
      RECT  0.465000  6.750000  1.310000  7.170000 ;
      RECT  0.465000  7.170000  5.120000  7.310000 ;
      RECT  0.465000  7.310000  1.310000  7.730000 ;
      RECT  0.465000  7.730000  5.120000  7.870000 ;
      RECT  0.465000  7.870000  1.310000  8.290000 ;
      RECT  0.465000  8.290000  5.120000  8.430000 ;
      RECT  0.465000  8.430000  1.310000  8.850000 ;
      RECT  0.465000  8.850000  5.120000  8.990000 ;
      RECT  0.465000  8.990000  1.310000  9.410000 ;
      RECT  0.465000  9.410000  5.120000  9.550000 ;
      RECT  0.465000  9.550000  1.310000 10.000000 ;
      RECT  0.465000 10.000000  5.120000 10.270000 ;
      RECT  0.465000 10.270000  1.215000 11.605000 ;
      RECT  0.465000 11.605000 21.285000 11.755000 ;
      RECT  0.465000 11.755000  1.215000 12.960000 ;
      RECT  0.465000 12.960000  5.120000 13.230000 ;
      RECT  0.465000 13.230000  1.310000 13.680000 ;
      RECT  0.465000 13.680000  5.120000 13.820000 ;
      RECT  0.465000 13.820000  1.310000 14.240000 ;
      RECT  0.465000 14.240000  5.120000 14.380000 ;
      RECT  0.465000 14.380000  1.310000 14.800000 ;
      RECT  0.465000 14.800000  5.120000 14.940000 ;
      RECT  0.465000 14.940000  1.310000 15.360000 ;
      RECT  0.465000 15.360000  5.120000 15.500000 ;
      RECT  0.465000 15.500000  1.310000 15.920000 ;
      RECT  0.465000 15.920000  5.120000 16.060000 ;
      RECT  0.465000 16.060000  1.310000 16.480000 ;
      RECT  0.465000 16.480000  5.120000 16.620000 ;
      RECT  0.465000 16.620000  1.310000 18.150000 ;
      RECT  0.465000 18.150000  5.120000 18.290000 ;
      RECT  0.465000 18.290000  1.310000 18.710000 ;
      RECT  0.465000 18.710000  5.120000 18.850000 ;
      RECT  0.465000 18.850000  1.310000 19.270000 ;
      RECT  0.465000 19.270000  5.120000 19.410000 ;
      RECT  0.465000 19.410000  1.310000 19.830000 ;
      RECT  0.465000 19.830000  5.120000 19.970000 ;
      RECT  0.465000 19.970000  1.310000 20.390000 ;
      RECT  0.465000 20.390000  5.120000 20.530000 ;
      RECT  0.465000 20.530000  1.310000 20.950000 ;
      RECT  0.465000 20.950000  5.120000 21.090000 ;
      RECT  0.465000 21.090000  1.310000 21.540000 ;
      RECT  0.465000 21.540000  5.120000 21.810000 ;
      RECT  0.465000 21.810000  1.215000 23.145000 ;
      RECT  0.465000 23.145000 21.285000 23.295000 ;
      RECT  1.355000  0.355000  9.980000  1.270000 ;
      RECT  1.355000 10.420000  9.980000 11.465000 ;
      RECT  1.355000 11.895000  9.980000 12.810000 ;
      RECT  1.355000 21.960000  9.980000 23.005000 ;
      RECT  1.450000  1.860000  9.890000  2.000000 ;
      RECT  1.450000  2.420000  9.890000  2.560000 ;
      RECT  1.450000  2.980000  9.890000  3.120000 ;
      RECT  1.450000  3.540000  9.890000  3.680000 ;
      RECT  1.450000  4.100000  9.890000  4.240000 ;
      RECT  1.450000  4.660000  9.890000  4.800000 ;
      RECT  1.450000  5.220000  9.890000  5.360000 ;
      RECT  1.450000  5.530000  9.890000  6.160000 ;
      RECT  1.450000  6.330000  9.890000  6.470000 ;
      RECT  1.450000  6.890000  9.890000  7.030000 ;
      RECT  1.450000  7.450000  9.890000  7.590000 ;
      RECT  1.450000  8.010000  9.890000  8.150000 ;
      RECT  1.450000  8.570000  9.890000  8.710000 ;
      RECT  1.450000  9.130000  9.890000  9.270000 ;
      RECT  1.450000  9.690000  9.890000  9.830000 ;
      RECT  1.450000 13.400000  9.890000 13.540000 ;
      RECT  1.450000 13.960000  9.890000 14.100000 ;
      RECT  1.450000 14.520000  9.890000 14.660000 ;
      RECT  1.450000 15.080000  9.890000 15.220000 ;
      RECT  1.450000 15.640000  9.890000 15.780000 ;
      RECT  1.450000 16.200000  9.890000 16.340000 ;
      RECT  1.450000 16.760000  9.890000 16.900000 ;
      RECT  1.450000 17.070000  9.890000 17.700000 ;
      RECT  1.450000 17.870000  9.890000 18.010000 ;
      RECT  1.450000 18.430000  9.890000 18.570000 ;
      RECT  1.450000 18.990000  9.890000 19.130000 ;
      RECT  1.450000 19.550000  9.890000 19.690000 ;
      RECT  1.450000 20.110000  9.890000 20.250000 ;
      RECT  1.450000 20.670000  9.890000 20.810000 ;
      RECT  1.450000 21.230000  9.890000 21.370000 ;
      RECT  5.260000  1.270000  6.080000  1.860000 ;
      RECT  5.260000  2.000000  6.080000  2.420000 ;
      RECT  5.260000  2.560000  6.080000  2.980000 ;
      RECT  5.260000  3.120000  6.080000  3.540000 ;
      RECT  5.260000  3.680000  6.080000  4.100000 ;
      RECT  5.260000  4.240000  6.080000  4.660000 ;
      RECT  5.260000  4.800000  6.080000  5.220000 ;
      RECT  5.260000  5.360000  6.080000  5.530000 ;
      RECT  5.260000  6.160000  6.080000  6.330000 ;
      RECT  5.260000  6.470000  6.080000  6.890000 ;
      RECT  5.260000  7.030000  6.080000  7.450000 ;
      RECT  5.260000  7.590000  6.080000  8.010000 ;
      RECT  5.260000  8.150000  6.080000  8.570000 ;
      RECT  5.260000  8.710000  6.080000  9.130000 ;
      RECT  5.260000  9.270000  6.080000  9.690000 ;
      RECT  5.260000  9.830000  6.080000 10.420000 ;
      RECT  5.260000 12.810000  6.080000 13.400000 ;
      RECT  5.260000 13.540000  6.080000 13.960000 ;
      RECT  5.260000 14.100000  6.080000 14.520000 ;
      RECT  5.260000 14.660000  6.080000 15.080000 ;
      RECT  5.260000 15.220000  6.080000 15.640000 ;
      RECT  5.260000 15.780000  6.080000 16.200000 ;
      RECT  5.260000 16.340000  6.080000 16.760000 ;
      RECT  5.260000 16.900000  6.080000 17.070000 ;
      RECT  5.260000 17.700000  6.080000 17.870000 ;
      RECT  5.260000 18.010000  6.080000 18.430000 ;
      RECT  5.260000 18.570000  6.080000 18.990000 ;
      RECT  5.260000 19.130000  6.080000 19.550000 ;
      RECT  5.260000 19.690000  6.080000 20.110000 ;
      RECT  5.260000 20.250000  6.080000 20.670000 ;
      RECT  5.260000 20.810000  6.080000 21.230000 ;
      RECT  5.260000 21.370000  6.080000 21.960000 ;
      RECT  6.220000  1.420000 15.530000  1.690000 ;
      RECT  6.220000  2.140000 15.530000  2.280000 ;
      RECT  6.220000  2.700000 15.530000  2.840000 ;
      RECT  6.220000  3.260000 15.530000  3.400000 ;
      RECT  6.220000  3.820000 15.530000  3.960000 ;
      RECT  6.220000  4.380000 15.530000  4.520000 ;
      RECT  6.220000  4.940000 15.530000  5.080000 ;
      RECT  6.220000  6.610000 15.530000  6.750000 ;
      RECT  6.220000  7.170000 15.530000  7.310000 ;
      RECT  6.220000  7.730000 15.530000  7.870000 ;
      RECT  6.220000  8.290000 15.530000  8.430000 ;
      RECT  6.220000  8.850000 15.530000  8.990000 ;
      RECT  6.220000  9.410000 15.530000  9.550000 ;
      RECT  6.220000 10.000000 15.530000 10.270000 ;
      RECT  6.220000 12.960000 15.530000 13.230000 ;
      RECT  6.220000 13.680000 15.530000 13.820000 ;
      RECT  6.220000 14.240000 15.530000 14.380000 ;
      RECT  6.220000 14.800000 15.530000 14.940000 ;
      RECT  6.220000 15.360000 15.530000 15.500000 ;
      RECT  6.220000 15.920000 15.530000 16.060000 ;
      RECT  6.220000 16.480000 15.530000 16.620000 ;
      RECT  6.220000 18.150000 15.530000 18.290000 ;
      RECT  6.220000 18.710000 15.530000 18.850000 ;
      RECT  6.220000 19.270000 15.530000 19.410000 ;
      RECT  6.220000 19.830000 15.530000 19.970000 ;
      RECT  6.220000 20.390000 15.530000 20.530000 ;
      RECT  6.220000 20.950000 15.530000 21.090000 ;
      RECT  6.220000 21.540000 15.530000 21.810000 ;
      RECT 10.030000  1.690000 11.720000  2.140000 ;
      RECT 10.030000  2.280000 11.720000  2.700000 ;
      RECT 10.030000  2.840000 11.720000  3.260000 ;
      RECT 10.030000  3.400000 11.720000  3.820000 ;
      RECT 10.030000  3.960000 11.720000  4.380000 ;
      RECT 10.030000  4.520000 11.720000  4.940000 ;
      RECT 10.030000  5.080000 11.720000  6.610000 ;
      RECT 10.030000  6.750000 11.720000  7.170000 ;
      RECT 10.030000  7.310000 11.720000  7.730000 ;
      RECT 10.030000  7.870000 11.720000  8.290000 ;
      RECT 10.030000  8.430000 11.720000  8.850000 ;
      RECT 10.030000  8.990000 11.720000  9.410000 ;
      RECT 10.030000  9.550000 11.720000 10.000000 ;
      RECT 10.030000 13.230000 11.720000 13.680000 ;
      RECT 10.030000 13.820000 11.720000 14.240000 ;
      RECT 10.030000 14.380000 11.720000 14.800000 ;
      RECT 10.030000 14.940000 11.720000 15.360000 ;
      RECT 10.030000 15.500000 11.720000 15.920000 ;
      RECT 10.030000 16.060000 11.720000 16.480000 ;
      RECT 10.030000 16.620000 11.720000 18.150000 ;
      RECT 10.030000 18.290000 11.720000 18.710000 ;
      RECT 10.030000 18.850000 11.720000 19.270000 ;
      RECT 10.030000 19.410000 11.720000 19.830000 ;
      RECT 10.030000 19.970000 11.720000 20.390000 ;
      RECT 10.030000 20.530000 11.720000 20.950000 ;
      RECT 10.030000 21.090000 11.720000 21.540000 ;
      RECT 10.120000  0.215000 11.625000  1.420000 ;
      RECT 10.120000 10.270000 11.625000 11.605000 ;
      RECT 10.120000 11.755000 11.625000 12.960000 ;
      RECT 10.120000 21.810000 11.625000 23.145000 ;
      RECT 11.765000  0.355000 20.390000  1.270000 ;
      RECT 11.765000 10.420000 20.390000 11.465000 ;
      RECT 11.765000 11.895000 20.390000 12.810000 ;
      RECT 11.765000 21.960000 20.390000 23.005000 ;
      RECT 11.860000  1.860000 20.300000  2.000000 ;
      RECT 11.860000  2.420000 20.300000  2.560000 ;
      RECT 11.860000  2.980000 20.300000  3.120000 ;
      RECT 11.860000  3.540000 20.300000  3.680000 ;
      RECT 11.860000  4.100000 20.300000  4.240000 ;
      RECT 11.860000  4.660000 20.300000  4.800000 ;
      RECT 11.860000  5.220000 20.300000  5.360000 ;
      RECT 11.860000  5.530000 20.300000  6.160000 ;
      RECT 11.860000  6.330000 20.300000  6.470000 ;
      RECT 11.860000  6.890000 20.300000  7.030000 ;
      RECT 11.860000  7.450000 20.300000  7.590000 ;
      RECT 11.860000  8.010000 20.300000  8.150000 ;
      RECT 11.860000  8.570000 20.300000  8.710000 ;
      RECT 11.860000  9.130000 20.300000  9.270000 ;
      RECT 11.860000  9.690000 20.300000  9.830000 ;
      RECT 11.860000 13.400000 20.300000 13.540000 ;
      RECT 11.860000 13.960000 20.300000 14.100000 ;
      RECT 11.860000 14.520000 20.300000 14.660000 ;
      RECT 11.860000 15.080000 20.300000 15.220000 ;
      RECT 11.860000 15.640000 20.300000 15.780000 ;
      RECT 11.860000 16.200000 20.300000 16.340000 ;
      RECT 11.860000 16.760000 20.300000 16.900000 ;
      RECT 11.860000 17.070000 20.300000 17.700000 ;
      RECT 11.860000 17.870000 20.300000 18.010000 ;
      RECT 11.860000 18.430000 20.300000 18.570000 ;
      RECT 11.860000 18.990000 20.300000 19.130000 ;
      RECT 11.860000 19.550000 20.300000 19.690000 ;
      RECT 11.860000 20.110000 20.300000 20.250000 ;
      RECT 11.860000 20.670000 20.300000 20.810000 ;
      RECT 11.860000 21.230000 20.300000 21.370000 ;
      RECT 15.670000  1.270000 16.490000  1.860000 ;
      RECT 15.670000  2.000000 16.490000  2.420000 ;
      RECT 15.670000  2.560000 16.490000  2.980000 ;
      RECT 15.670000  3.120000 16.490000  3.540000 ;
      RECT 15.670000  3.680000 16.490000  4.100000 ;
      RECT 15.670000  4.240000 16.490000  4.660000 ;
      RECT 15.670000  4.800000 16.490000  5.220000 ;
      RECT 15.670000  5.360000 16.490000  5.530000 ;
      RECT 15.670000  6.160000 16.490000  6.330000 ;
      RECT 15.670000  6.470000 16.490000  6.890000 ;
      RECT 15.670000  7.030000 16.490000  7.450000 ;
      RECT 15.670000  7.590000 16.490000  8.010000 ;
      RECT 15.670000  8.150000 16.490000  8.570000 ;
      RECT 15.670000  8.710000 16.490000  9.130000 ;
      RECT 15.670000  9.270000 16.490000  9.690000 ;
      RECT 15.670000  9.830000 16.490000 10.420000 ;
      RECT 15.670000 12.810000 16.490000 13.400000 ;
      RECT 15.670000 13.540000 16.490000 13.960000 ;
      RECT 15.670000 14.100000 16.490000 14.520000 ;
      RECT 15.670000 14.660000 16.490000 15.080000 ;
      RECT 15.670000 15.220000 16.490000 15.640000 ;
      RECT 15.670000 15.780000 16.490000 16.200000 ;
      RECT 15.670000 16.340000 16.490000 16.760000 ;
      RECT 15.670000 16.900000 16.490000 17.070000 ;
      RECT 15.670000 17.700000 16.490000 17.870000 ;
      RECT 15.670000 18.010000 16.490000 18.430000 ;
      RECT 15.670000 18.570000 16.490000 18.990000 ;
      RECT 15.670000 19.130000 16.490000 19.550000 ;
      RECT 15.670000 19.690000 16.490000 20.110000 ;
      RECT 15.670000 20.250000 16.490000 20.670000 ;
      RECT 15.670000 20.810000 16.490000 21.230000 ;
      RECT 15.670000 21.370000 16.490000 21.960000 ;
      RECT 16.630000  1.420000 21.285000  1.690000 ;
      RECT 16.630000  2.140000 21.285000  2.280000 ;
      RECT 16.630000  2.700000 21.285000  2.840000 ;
      RECT 16.630000  3.260000 21.285000  3.400000 ;
      RECT 16.630000  3.820000 21.285000  3.960000 ;
      RECT 16.630000  4.380000 21.285000  4.520000 ;
      RECT 16.630000  4.940000 21.285000  5.080000 ;
      RECT 16.630000  6.610000 21.285000  6.750000 ;
      RECT 16.630000  7.170000 21.285000  7.310000 ;
      RECT 16.630000  7.730000 21.285000  7.870000 ;
      RECT 16.630000  8.290000 21.285000  8.430000 ;
      RECT 16.630000  8.850000 21.285000  8.990000 ;
      RECT 16.630000  9.410000 21.285000  9.550000 ;
      RECT 16.630000 10.000000 21.285000 10.270000 ;
      RECT 16.630000 12.960000 21.285000 13.230000 ;
      RECT 16.630000 13.680000 21.285000 13.820000 ;
      RECT 16.630000 14.240000 21.285000 14.380000 ;
      RECT 16.630000 14.800000 21.285000 14.940000 ;
      RECT 16.630000 15.360000 21.285000 15.500000 ;
      RECT 16.630000 15.920000 21.285000 16.060000 ;
      RECT 16.630000 16.480000 21.285000 16.620000 ;
      RECT 16.630000 18.150000 21.285000 18.290000 ;
      RECT 16.630000 18.710000 21.285000 18.850000 ;
      RECT 16.630000 19.270000 21.285000 19.410000 ;
      RECT 16.630000 19.830000 21.285000 19.970000 ;
      RECT 16.630000 20.390000 21.285000 20.530000 ;
      RECT 16.630000 20.950000 21.285000 21.090000 ;
      RECT 16.630000 21.540000 21.285000 21.810000 ;
      RECT 20.440000  1.690000 21.285000  2.140000 ;
      RECT 20.440000  2.280000 21.285000  2.700000 ;
      RECT 20.440000  2.840000 21.285000  3.260000 ;
      RECT 20.440000  3.400000 21.285000  3.820000 ;
      RECT 20.440000  3.960000 21.285000  4.380000 ;
      RECT 20.440000  4.520000 21.285000  4.940000 ;
      RECT 20.440000  5.080000 21.285000  6.610000 ;
      RECT 20.440000  6.750000 21.285000  7.170000 ;
      RECT 20.440000  7.310000 21.285000  7.730000 ;
      RECT 20.440000  7.870000 21.285000  8.290000 ;
      RECT 20.440000  8.430000 21.285000  8.850000 ;
      RECT 20.440000  8.990000 21.285000  9.410000 ;
      RECT 20.440000  9.550000 21.285000 10.000000 ;
      RECT 20.440000 13.230000 21.285000 13.680000 ;
      RECT 20.440000 13.820000 21.285000 14.240000 ;
      RECT 20.440000 14.380000 21.285000 14.800000 ;
      RECT 20.440000 14.940000 21.285000 15.360000 ;
      RECT 20.440000 15.500000 21.285000 15.920000 ;
      RECT 20.440000 16.060000 21.285000 16.480000 ;
      RECT 20.440000 16.620000 21.285000 18.150000 ;
      RECT 20.440000 18.290000 21.285000 18.710000 ;
      RECT 20.440000 18.850000 21.285000 19.270000 ;
      RECT 20.440000 19.410000 21.285000 19.830000 ;
      RECT 20.440000 19.970000 21.285000 20.390000 ;
      RECT 20.440000 20.530000 21.285000 20.950000 ;
      RECT 20.440000 21.090000 21.285000 21.540000 ;
      RECT 20.530000  0.215000 21.285000  1.420000 ;
      RECT 20.530000 10.270000 21.285000 11.605000 ;
      RECT 20.530000 11.755000 21.285000 12.960000 ;
      RECT 20.530000 21.810000 21.285000 23.145000 ;
    LAYER met2 ;
      RECT  0.325000  0.140000 21.425000  1.270000 ;
      RECT  0.325000  1.270000  0.845000 10.420000 ;
      RECT  0.325000 10.420000 21.425000 12.810000 ;
      RECT  0.325000 12.810000  0.845000 21.960000 ;
      RECT  0.325000 21.960000 21.425000 23.220000 ;
      RECT  0.990000  1.420000  5.120000  1.690000 ;
      RECT  0.990000  1.690000  1.310000  1.860000 ;
      RECT  0.990000  1.860000  5.120000  2.000000 ;
      RECT  0.990000  2.000000  1.310000  2.420000 ;
      RECT  0.990000  2.420000  5.120000  2.560000 ;
      RECT  0.990000  2.560000  1.310000  2.980000 ;
      RECT  0.990000  2.980000  5.120000  3.120000 ;
      RECT  0.990000  3.120000  1.310000  3.540000 ;
      RECT  0.990000  3.540000  5.120000  3.680000 ;
      RECT  0.990000  3.680000  1.310000  4.100000 ;
      RECT  0.990000  4.100000  5.120000  4.240000 ;
      RECT  0.990000  4.240000  1.310000  4.660000 ;
      RECT  0.990000  4.660000  5.120000  4.800000 ;
      RECT  0.990000  4.800000  1.310000  5.220000 ;
      RECT  0.990000  5.220000  5.120000  5.360000 ;
      RECT  0.990000  5.360000  1.310000  6.330000 ;
      RECT  0.990000  6.330000  5.120000  6.470000 ;
      RECT  0.990000  6.470000  1.310000  6.890000 ;
      RECT  0.990000  6.890000  5.120000  7.030000 ;
      RECT  0.990000  7.030000  1.310000  7.450000 ;
      RECT  0.990000  7.450000  5.120000  7.590000 ;
      RECT  0.990000  7.590000  1.310000  8.010000 ;
      RECT  0.990000  8.010000  5.120000  8.150000 ;
      RECT  0.990000  8.150000  1.310000  8.570000 ;
      RECT  0.990000  8.570000  5.120000  8.710000 ;
      RECT  0.990000  8.710000  1.310000  9.130000 ;
      RECT  0.990000  9.130000  5.120000  9.270000 ;
      RECT  0.990000  9.270000  1.310000  9.690000 ;
      RECT  0.990000  9.690000  5.120000  9.830000 ;
      RECT  0.990000  9.830000  1.310000 10.000000 ;
      RECT  0.990000 10.000000  5.120000 10.270000 ;
      RECT  0.990000 12.960000  5.120000 13.230000 ;
      RECT  0.990000 13.230000  1.310000 13.400000 ;
      RECT  0.990000 13.400000  5.120000 13.540000 ;
      RECT  0.990000 13.540000  1.310000 13.960000 ;
      RECT  0.990000 13.960000  5.120000 14.100000 ;
      RECT  0.990000 14.100000  1.310000 14.520000 ;
      RECT  0.990000 14.520000  5.120000 14.660000 ;
      RECT  0.990000 14.660000  1.310000 15.080000 ;
      RECT  0.990000 15.080000  5.120000 15.220000 ;
      RECT  0.990000 15.220000  1.310000 15.640000 ;
      RECT  0.990000 15.640000  5.120000 15.780000 ;
      RECT  0.990000 15.780000  1.310000 16.200000 ;
      RECT  0.990000 16.200000  5.120000 16.340000 ;
      RECT  0.990000 16.340000  1.310000 16.760000 ;
      RECT  0.990000 16.760000  5.120000 16.900000 ;
      RECT  0.990000 16.900000  1.310000 17.870000 ;
      RECT  0.990000 17.870000  5.120000 18.010000 ;
      RECT  0.990000 18.010000  1.310000 18.430000 ;
      RECT  0.990000 18.430000  5.120000 18.570000 ;
      RECT  0.990000 18.570000  1.310000 18.990000 ;
      RECT  0.990000 18.990000  5.120000 19.130000 ;
      RECT  0.990000 19.130000  1.310000 19.550000 ;
      RECT  0.990000 19.550000  5.120000 19.690000 ;
      RECT  0.990000 19.690000  1.310000 20.110000 ;
      RECT  0.990000 20.110000  5.120000 20.250000 ;
      RECT  0.990000 20.250000  1.310000 20.670000 ;
      RECT  0.990000 20.670000  5.120000 20.810000 ;
      RECT  0.990000 20.810000  1.310000 21.230000 ;
      RECT  0.990000 21.230000  5.120000 21.370000 ;
      RECT  0.990000 21.370000  1.310000 21.540000 ;
      RECT  0.990000 21.540000  5.120000 21.810000 ;
      RECT  1.450000  2.140000  9.890000  2.280000 ;
      RECT  1.450000  2.700000  9.890000  2.840000 ;
      RECT  1.450000  3.260000  9.890000  3.400000 ;
      RECT  1.450000  3.820000  9.890000  3.960000 ;
      RECT  1.450000  4.380000  9.890000  4.520000 ;
      RECT  1.450000  4.940000  9.890000  5.080000 ;
      RECT  1.450000  5.530000  9.890000  6.160000 ;
      RECT  1.450000  6.610000  9.890000  6.750000 ;
      RECT  1.450000  7.170000  9.890000  7.310000 ;
      RECT  1.450000  7.730000  9.890000  7.870000 ;
      RECT  1.450000  8.290000  9.890000  8.430000 ;
      RECT  1.450000  8.850000  9.890000  8.990000 ;
      RECT  1.450000  9.410000  9.890000  9.550000 ;
      RECT  1.450000 13.680000  9.890000 13.820000 ;
      RECT  1.450000 14.240000  9.890000 14.380000 ;
      RECT  1.450000 14.800000  9.890000 14.940000 ;
      RECT  1.450000 15.360000  9.890000 15.500000 ;
      RECT  1.450000 15.920000  9.890000 16.060000 ;
      RECT  1.450000 16.480000  9.890000 16.620000 ;
      RECT  1.450000 17.070000  9.890000 17.700000 ;
      RECT  1.450000 18.150000  9.890000 18.290000 ;
      RECT  1.450000 18.710000  9.890000 18.850000 ;
      RECT  1.450000 19.270000  9.890000 19.410000 ;
      RECT  1.450000 19.830000  9.890000 19.970000 ;
      RECT  1.450000 20.390000  9.890000 20.530000 ;
      RECT  1.450000 20.950000  9.890000 21.090000 ;
      RECT  5.260000  1.270000  6.080000  2.140000 ;
      RECT  5.260000  2.280000  6.080000  2.700000 ;
      RECT  5.260000  2.840000  6.080000  3.260000 ;
      RECT  5.260000  3.400000  6.080000  3.820000 ;
      RECT  5.260000  3.960000  6.080000  4.380000 ;
      RECT  5.260000  4.520000  6.080000  4.940000 ;
      RECT  5.260000  5.080000  6.080000  5.530000 ;
      RECT  5.260000  6.160000  6.080000  6.610000 ;
      RECT  5.260000  6.750000  6.080000  7.170000 ;
      RECT  5.260000  7.310000  6.080000  7.730000 ;
      RECT  5.260000  7.870000  6.080000  8.290000 ;
      RECT  5.260000  8.430000  6.080000  8.850000 ;
      RECT  5.260000  8.990000  6.080000  9.410000 ;
      RECT  5.260000  9.550000  6.080000 10.420000 ;
      RECT  5.260000 12.810000  6.080000 13.680000 ;
      RECT  5.260000 13.820000  6.080000 14.240000 ;
      RECT  5.260000 14.380000  6.080000 14.800000 ;
      RECT  5.260000 14.940000  6.080000 15.360000 ;
      RECT  5.260000 15.500000  6.080000 15.920000 ;
      RECT  5.260000 16.060000  6.080000 16.480000 ;
      RECT  5.260000 16.620000  6.080000 17.070000 ;
      RECT  5.260000 17.700000  6.080000 18.150000 ;
      RECT  5.260000 18.290000  6.080000 18.710000 ;
      RECT  5.260000 18.850000  6.080000 19.270000 ;
      RECT  5.260000 19.410000  6.080000 19.830000 ;
      RECT  5.260000 19.970000  6.080000 20.390000 ;
      RECT  5.260000 20.530000  6.080000 20.950000 ;
      RECT  5.260000 21.090000  6.080000 21.960000 ;
      RECT  6.220000  1.420000 10.350000  1.690000 ;
      RECT  6.220000  1.860000 10.350000  2.000000 ;
      RECT  6.220000  2.420000 10.350000  2.560000 ;
      RECT  6.220000  2.980000 10.350000  3.120000 ;
      RECT  6.220000  3.540000 10.350000  3.680000 ;
      RECT  6.220000  4.100000 10.350000  4.240000 ;
      RECT  6.220000  4.660000 10.350000  4.800000 ;
      RECT  6.220000  5.220000 10.350000  5.360000 ;
      RECT  6.220000  6.330000 10.350000  6.470000 ;
      RECT  6.220000  6.890000 10.350000  7.030000 ;
      RECT  6.220000  7.450000 10.350000  7.590000 ;
      RECT  6.220000  8.010000 10.350000  8.150000 ;
      RECT  6.220000  8.570000 10.350000  8.710000 ;
      RECT  6.220000  9.130000 10.350000  9.270000 ;
      RECT  6.220000  9.690000 10.350000  9.830000 ;
      RECT  6.220000 10.000000 10.350000 10.270000 ;
      RECT  6.220000 12.960000 10.350000 13.230000 ;
      RECT  6.220000 13.400000 10.350000 13.540000 ;
      RECT  6.220000 13.960000 10.350000 14.100000 ;
      RECT  6.220000 14.520000 10.350000 14.660000 ;
      RECT  6.220000 15.080000 10.350000 15.220000 ;
      RECT  6.220000 15.640000 10.350000 15.780000 ;
      RECT  6.220000 16.200000 10.350000 16.340000 ;
      RECT  6.220000 16.760000 10.350000 16.900000 ;
      RECT  6.220000 17.870000 10.350000 18.010000 ;
      RECT  6.220000 18.430000 10.350000 18.570000 ;
      RECT  6.220000 18.990000 10.350000 19.130000 ;
      RECT  6.220000 19.550000 10.350000 19.690000 ;
      RECT  6.220000 20.110000 10.350000 20.250000 ;
      RECT  6.220000 20.670000 10.350000 20.810000 ;
      RECT  6.220000 21.230000 10.350000 21.370000 ;
      RECT  6.220000 21.540000 10.350000 21.810000 ;
      RECT 10.030000  1.690000 10.350000  1.860000 ;
      RECT 10.030000  2.000000 10.350000  2.420000 ;
      RECT 10.030000  2.560000 10.350000  2.980000 ;
      RECT 10.030000  3.120000 10.350000  3.540000 ;
      RECT 10.030000  3.680000 10.350000  4.100000 ;
      RECT 10.030000  4.240000 10.350000  4.660000 ;
      RECT 10.030000  4.800000 10.350000  5.220000 ;
      RECT 10.030000  5.360000 10.350000  6.330000 ;
      RECT 10.030000  6.470000 10.350000  6.890000 ;
      RECT 10.030000  7.030000 10.350000  7.450000 ;
      RECT 10.030000  7.590000 10.350000  8.010000 ;
      RECT 10.030000  8.150000 10.350000  8.570000 ;
      RECT 10.030000  8.710000 10.350000  9.130000 ;
      RECT 10.030000  9.270000 10.350000  9.690000 ;
      RECT 10.030000  9.830000 10.350000 10.000000 ;
      RECT 10.030000 13.230000 10.350000 13.400000 ;
      RECT 10.030000 13.540000 10.350000 13.960000 ;
      RECT 10.030000 14.100000 10.350000 14.520000 ;
      RECT 10.030000 14.660000 10.350000 15.080000 ;
      RECT 10.030000 15.220000 10.350000 15.640000 ;
      RECT 10.030000 15.780000 10.350000 16.200000 ;
      RECT 10.030000 16.340000 10.350000 16.760000 ;
      RECT 10.030000 16.900000 10.350000 17.870000 ;
      RECT 10.030000 18.010000 10.350000 18.430000 ;
      RECT 10.030000 18.570000 10.350000 18.990000 ;
      RECT 10.030000 19.130000 10.350000 19.550000 ;
      RECT 10.030000 19.690000 10.350000 20.110000 ;
      RECT 10.030000 20.250000 10.350000 20.670000 ;
      RECT 10.030000 20.810000 10.350000 21.230000 ;
      RECT 10.030000 21.370000 10.350000 21.540000 ;
      RECT 10.490000  1.270000 11.255000 10.420000 ;
      RECT 10.490000 12.810000 11.255000 21.960000 ;
      RECT 11.400000  1.420000 15.530000  1.690000 ;
      RECT 11.400000  1.690000 11.720000  1.860000 ;
      RECT 11.400000  1.860000 15.530000  2.000000 ;
      RECT 11.400000  2.000000 11.720000  2.420000 ;
      RECT 11.400000  2.420000 15.530000  2.560000 ;
      RECT 11.400000  2.560000 11.720000  2.980000 ;
      RECT 11.400000  2.980000 15.530000  3.120000 ;
      RECT 11.400000  3.120000 11.720000  3.540000 ;
      RECT 11.400000  3.540000 15.530000  3.680000 ;
      RECT 11.400000  3.680000 11.720000  4.100000 ;
      RECT 11.400000  4.100000 15.530000  4.240000 ;
      RECT 11.400000  4.240000 11.720000  4.660000 ;
      RECT 11.400000  4.660000 15.530000  4.800000 ;
      RECT 11.400000  4.800000 11.720000  5.220000 ;
      RECT 11.400000  5.220000 15.530000  5.360000 ;
      RECT 11.400000  5.360000 11.720000  6.330000 ;
      RECT 11.400000  6.330000 15.530000  6.470000 ;
      RECT 11.400000  6.470000 11.720000  6.890000 ;
      RECT 11.400000  6.890000 15.530000  7.030000 ;
      RECT 11.400000  7.030000 11.720000  7.450000 ;
      RECT 11.400000  7.450000 15.530000  7.590000 ;
      RECT 11.400000  7.590000 11.720000  8.010000 ;
      RECT 11.400000  8.010000 15.530000  8.150000 ;
      RECT 11.400000  8.150000 11.720000  8.570000 ;
      RECT 11.400000  8.570000 15.530000  8.710000 ;
      RECT 11.400000  8.710000 11.720000  9.130000 ;
      RECT 11.400000  9.130000 15.530000  9.270000 ;
      RECT 11.400000  9.270000 11.720000  9.690000 ;
      RECT 11.400000  9.690000 15.530000  9.830000 ;
      RECT 11.400000  9.830000 11.720000 10.000000 ;
      RECT 11.400000 10.000000 15.530000 10.270000 ;
      RECT 11.400000 12.960000 15.530000 13.230000 ;
      RECT 11.400000 13.230000 11.720000 13.400000 ;
      RECT 11.400000 13.400000 15.530000 13.540000 ;
      RECT 11.400000 13.540000 11.720000 13.960000 ;
      RECT 11.400000 13.960000 15.530000 14.100000 ;
      RECT 11.400000 14.100000 11.720000 14.520000 ;
      RECT 11.400000 14.520000 15.530000 14.660000 ;
      RECT 11.400000 14.660000 11.720000 15.080000 ;
      RECT 11.400000 15.080000 15.530000 15.220000 ;
      RECT 11.400000 15.220000 11.720000 15.640000 ;
      RECT 11.400000 15.640000 15.530000 15.780000 ;
      RECT 11.400000 15.780000 11.720000 16.200000 ;
      RECT 11.400000 16.200000 15.530000 16.340000 ;
      RECT 11.400000 16.340000 11.720000 16.760000 ;
      RECT 11.400000 16.760000 15.530000 16.900000 ;
      RECT 11.400000 16.900000 11.720000 17.870000 ;
      RECT 11.400000 17.870000 15.530000 18.010000 ;
      RECT 11.400000 18.010000 11.720000 18.430000 ;
      RECT 11.400000 18.430000 15.530000 18.570000 ;
      RECT 11.400000 18.570000 11.720000 18.990000 ;
      RECT 11.400000 18.990000 15.530000 19.130000 ;
      RECT 11.400000 19.130000 11.720000 19.550000 ;
      RECT 11.400000 19.550000 15.530000 19.690000 ;
      RECT 11.400000 19.690000 11.720000 20.110000 ;
      RECT 11.400000 20.110000 15.530000 20.250000 ;
      RECT 11.400000 20.250000 11.720000 20.670000 ;
      RECT 11.400000 20.670000 15.530000 20.810000 ;
      RECT 11.400000 20.810000 11.720000 21.230000 ;
      RECT 11.400000 21.230000 15.530000 21.370000 ;
      RECT 11.400000 21.370000 11.720000 21.540000 ;
      RECT 11.400000 21.540000 15.530000 21.810000 ;
      RECT 11.860000  2.140000 20.300000  2.280000 ;
      RECT 11.860000  2.700000 20.300000  2.840000 ;
      RECT 11.860000  3.260000 20.300000  3.400000 ;
      RECT 11.860000  3.820000 20.300000  3.960000 ;
      RECT 11.860000  4.380000 20.300000  4.520000 ;
      RECT 11.860000  4.940000 20.300000  5.080000 ;
      RECT 11.860000  5.530000 20.300000  6.160000 ;
      RECT 11.860000  6.610000 20.300000  6.750000 ;
      RECT 11.860000  7.170000 20.300000  7.310000 ;
      RECT 11.860000  7.730000 20.300000  7.870000 ;
      RECT 11.860000  8.290000 20.300000  8.430000 ;
      RECT 11.860000  8.850000 20.300000  8.990000 ;
      RECT 11.860000  9.410000 20.300000  9.550000 ;
      RECT 11.860000 13.680000 20.300000 13.820000 ;
      RECT 11.860000 14.240000 20.300000 14.380000 ;
      RECT 11.860000 14.800000 20.300000 14.940000 ;
      RECT 11.860000 15.360000 20.300000 15.500000 ;
      RECT 11.860000 15.920000 20.300000 16.060000 ;
      RECT 11.860000 16.480000 20.300000 16.620000 ;
      RECT 11.860000 17.070000 20.300000 17.700000 ;
      RECT 11.860000 18.150000 20.300000 18.290000 ;
      RECT 11.860000 18.710000 20.300000 18.850000 ;
      RECT 11.860000 19.270000 20.300000 19.410000 ;
      RECT 11.860000 19.830000 20.300000 19.970000 ;
      RECT 11.860000 20.390000 20.300000 20.530000 ;
      RECT 11.860000 20.950000 20.300000 21.090000 ;
      RECT 15.670000  1.270000 16.490000  2.140000 ;
      RECT 15.670000  2.280000 16.490000  2.700000 ;
      RECT 15.670000  2.840000 16.490000  3.260000 ;
      RECT 15.670000  3.400000 16.490000  3.820000 ;
      RECT 15.670000  3.960000 16.490000  4.380000 ;
      RECT 15.670000  4.520000 16.490000  4.940000 ;
      RECT 15.670000  5.080000 16.490000  5.530000 ;
      RECT 15.670000  6.160000 16.490000  6.610000 ;
      RECT 15.670000  6.750000 16.490000  7.170000 ;
      RECT 15.670000  7.310000 16.490000  7.730000 ;
      RECT 15.670000  7.870000 16.490000  8.290000 ;
      RECT 15.670000  8.430000 16.490000  8.850000 ;
      RECT 15.670000  8.990000 16.490000  9.410000 ;
      RECT 15.670000  9.550000 16.490000 10.420000 ;
      RECT 15.670000 12.810000 16.490000 13.680000 ;
      RECT 15.670000 13.820000 16.490000 14.240000 ;
      RECT 15.670000 14.380000 16.490000 14.800000 ;
      RECT 15.670000 14.940000 16.490000 15.360000 ;
      RECT 15.670000 15.500000 16.490000 15.920000 ;
      RECT 15.670000 16.060000 16.490000 16.480000 ;
      RECT 15.670000 16.620000 16.490000 17.070000 ;
      RECT 15.670000 17.700000 16.490000 18.150000 ;
      RECT 15.670000 18.290000 16.490000 18.710000 ;
      RECT 15.670000 18.850000 16.490000 19.270000 ;
      RECT 15.670000 19.410000 16.490000 19.830000 ;
      RECT 15.670000 19.970000 16.490000 20.390000 ;
      RECT 15.670000 20.530000 16.490000 20.950000 ;
      RECT 15.670000 21.090000 16.490000 21.960000 ;
      RECT 16.630000  1.420000 20.760000  1.690000 ;
      RECT 16.630000  1.860000 20.760000  2.000000 ;
      RECT 16.630000  2.420000 20.760000  2.560000 ;
      RECT 16.630000  2.980000 20.760000  3.120000 ;
      RECT 16.630000  3.540000 20.760000  3.680000 ;
      RECT 16.630000  4.100000 20.760000  4.240000 ;
      RECT 16.630000  4.660000 20.760000  4.800000 ;
      RECT 16.630000  5.220000 20.760000  5.360000 ;
      RECT 16.630000  6.330000 20.760000  6.470000 ;
      RECT 16.630000  6.890000 20.760000  7.030000 ;
      RECT 16.630000  7.450000 20.760000  7.590000 ;
      RECT 16.630000  8.010000 20.760000  8.150000 ;
      RECT 16.630000  8.570000 20.760000  8.710000 ;
      RECT 16.630000  9.130000 20.760000  9.270000 ;
      RECT 16.630000  9.690000 20.760000  9.830000 ;
      RECT 16.630000 10.000000 20.760000 10.270000 ;
      RECT 16.630000 12.960000 20.760000 13.230000 ;
      RECT 16.630000 13.400000 20.760000 13.540000 ;
      RECT 16.630000 13.960000 20.760000 14.100000 ;
      RECT 16.630000 14.520000 20.760000 14.660000 ;
      RECT 16.630000 15.080000 20.760000 15.220000 ;
      RECT 16.630000 15.640000 20.760000 15.780000 ;
      RECT 16.630000 16.200000 20.760000 16.340000 ;
      RECT 16.630000 16.760000 20.760000 16.900000 ;
      RECT 16.630000 17.870000 20.760000 18.010000 ;
      RECT 16.630000 18.430000 20.760000 18.570000 ;
      RECT 16.630000 18.990000 20.760000 19.130000 ;
      RECT 16.630000 19.550000 20.760000 19.690000 ;
      RECT 16.630000 20.110000 20.760000 20.250000 ;
      RECT 16.630000 20.670000 20.760000 20.810000 ;
      RECT 16.630000 21.230000 20.760000 21.370000 ;
      RECT 16.630000 21.540000 20.760000 21.810000 ;
      RECT 20.440000  1.690000 20.760000  1.860000 ;
      RECT 20.440000  2.000000 20.760000  2.420000 ;
      RECT 20.440000  2.560000 20.760000  2.980000 ;
      RECT 20.440000  3.120000 20.760000  3.540000 ;
      RECT 20.440000  3.680000 20.760000  4.100000 ;
      RECT 20.440000  4.240000 20.760000  4.660000 ;
      RECT 20.440000  4.800000 20.760000  5.220000 ;
      RECT 20.440000  5.360000 20.760000  6.330000 ;
      RECT 20.440000  6.470000 20.760000  6.890000 ;
      RECT 20.440000  7.030000 20.760000  7.450000 ;
      RECT 20.440000  7.590000 20.760000  8.010000 ;
      RECT 20.440000  8.150000 20.760000  8.570000 ;
      RECT 20.440000  8.710000 20.760000  9.130000 ;
      RECT 20.440000  9.270000 20.760000  9.690000 ;
      RECT 20.440000  9.830000 20.760000 10.000000 ;
      RECT 20.440000 13.230000 20.760000 13.400000 ;
      RECT 20.440000 13.540000 20.760000 13.960000 ;
      RECT 20.440000 14.100000 20.760000 14.520000 ;
      RECT 20.440000 14.660000 20.760000 15.080000 ;
      RECT 20.440000 15.220000 20.760000 15.640000 ;
      RECT 20.440000 15.780000 20.760000 16.200000 ;
      RECT 20.440000 16.340000 20.760000 16.760000 ;
      RECT 20.440000 16.900000 20.760000 17.870000 ;
      RECT 20.440000 18.010000 20.760000 18.430000 ;
      RECT 20.440000 18.570000 20.760000 18.990000 ;
      RECT 20.440000 19.130000 20.760000 19.550000 ;
      RECT 20.440000 19.690000 20.760000 20.110000 ;
      RECT 20.440000 20.250000 20.760000 20.670000 ;
      RECT 20.440000 20.810000 20.760000 21.230000 ;
      RECT 20.440000 21.370000 20.760000 21.540000 ;
      RECT 20.900000  1.270000 21.425000 10.420000 ;
      RECT 20.900000 12.810000 21.425000 21.960000 ;
    LAYER met3 ;
      RECT  0.300000  0.140000  0.630000 23.220000 ;
      RECT  0.965000  0.235000 10.375000  0.565000 ;
      RECT  0.965000  0.565000  1.295000  1.465000 ;
      RECT  0.965000  1.465000  5.205000  1.765000 ;
      RECT  0.965000  1.765000  1.295000  2.665000 ;
      RECT  0.965000  2.665000  5.205000  2.965000 ;
      RECT  0.965000  2.965000  1.295000  3.865000 ;
      RECT  0.965000  3.865000  5.205000  4.165000 ;
      RECT  0.965000  4.165000  1.295000  5.065000 ;
      RECT  0.965000  5.065000  5.205000  5.365000 ;
      RECT  0.965000  5.365000  1.295000  6.295000 ;
      RECT  0.965000  6.295000  5.205000  6.595000 ;
      RECT  0.965000  6.595000  1.295000  7.495000 ;
      RECT  0.965000  7.495000  5.205000  7.795000 ;
      RECT  0.965000  7.795000  1.295000  8.695000 ;
      RECT  0.965000  8.695000  5.205000  8.995000 ;
      RECT  0.965000  8.995000  1.295000  9.895000 ;
      RECT  0.965000  9.895000  5.205000 10.195000 ;
      RECT  0.965000 10.195000  1.295000 11.095000 ;
      RECT  0.965000 11.095000 10.375000 11.425000 ;
      RECT  0.965000 11.775000 10.375000 12.105000 ;
      RECT  0.965000 12.105000  1.295000 13.005000 ;
      RECT  0.965000 13.005000  5.205000 13.305000 ;
      RECT  0.965000 13.305000  1.295000 14.205000 ;
      RECT  0.965000 14.205000  5.205000 14.505000 ;
      RECT  0.965000 14.505000  1.295000 15.405000 ;
      RECT  0.965000 15.405000  5.205000 15.705000 ;
      RECT  0.965000 15.705000  1.295000 16.605000 ;
      RECT  0.965000 16.605000  5.205000 16.905000 ;
      RECT  0.965000 16.905000  1.295000 17.835000 ;
      RECT  0.965000 17.835000  5.205000 18.135000 ;
      RECT  0.965000 18.135000  1.295000 19.035000 ;
      RECT  0.965000 19.035000  5.205000 19.335000 ;
      RECT  0.965000 19.335000  1.295000 20.235000 ;
      RECT  0.965000 20.235000  5.205000 20.535000 ;
      RECT  0.965000 20.535000  1.295000 21.435000 ;
      RECT  0.965000 21.435000  5.205000 21.735000 ;
      RECT  0.965000 21.735000  1.295000 22.635000 ;
      RECT  0.965000 22.635000 10.375000 22.965000 ;
      RECT  1.595000  0.865000  9.745000  1.165000 ;
      RECT  1.595000  2.065000  9.745000  2.365000 ;
      RECT  1.595000  3.265000  9.745000  3.565000 ;
      RECT  1.595000  4.465000  9.745000  4.765000 ;
      RECT  1.595000  5.665000  9.745000  5.995000 ;
      RECT  1.595000  6.895000  9.745000  7.195000 ;
      RECT  1.595000  8.095000  9.745000  8.395000 ;
      RECT  1.595000  9.295000  9.745000  9.595000 ;
      RECT  1.595000 10.495000  9.745000 10.795000 ;
      RECT  1.595000 12.405000  9.745000 12.705000 ;
      RECT  1.595000 13.605000  9.745000 13.905000 ;
      RECT  1.595000 14.805000  9.745000 15.105000 ;
      RECT  1.595000 16.005000  9.745000 16.305000 ;
      RECT  1.595000 17.205000  9.745000 17.535000 ;
      RECT  1.595000 18.435000  9.745000 18.735000 ;
      RECT  1.595000 19.635000  9.745000 19.935000 ;
      RECT  1.595000 20.835000  9.745000 21.135000 ;
      RECT  1.595000 22.035000  9.745000 22.335000 ;
      RECT  5.505000  1.165000  5.835000  2.065000 ;
      RECT  5.505000  2.365000  5.835000  3.265000 ;
      RECT  5.505000  3.565000  5.835000  4.465000 ;
      RECT  5.505000  4.765000  5.835000  5.665000 ;
      RECT  5.505000  5.995000  5.835000  6.895000 ;
      RECT  5.505000  7.195000  5.835000  8.095000 ;
      RECT  5.505000  8.395000  5.835000  9.295000 ;
      RECT  5.505000  9.595000  5.835000 10.495000 ;
      RECT  5.505000 12.705000  5.835000 13.605000 ;
      RECT  5.505000 13.905000  5.835000 14.805000 ;
      RECT  5.505000 15.105000  5.835000 16.005000 ;
      RECT  5.505000 16.305000  5.835000 17.205000 ;
      RECT  5.505000 17.535000  5.835000 18.435000 ;
      RECT  5.505000 18.735000  5.835000 19.635000 ;
      RECT  5.505000 19.935000  5.835000 20.835000 ;
      RECT  5.505000 21.135000  5.835000 22.035000 ;
      RECT  6.135000  1.465000 10.375000  1.765000 ;
      RECT  6.135000  2.665000 10.375000  2.965000 ;
      RECT  6.135000  3.865000 10.375000  4.165000 ;
      RECT  6.135000  5.065000 10.375000  5.365000 ;
      RECT  6.135000  6.295000 10.375000  6.595000 ;
      RECT  6.135000  7.495000 10.375000  7.795000 ;
      RECT  6.135000  8.695000 10.375000  8.995000 ;
      RECT  6.135000  9.895000 10.375000 10.195000 ;
      RECT  6.135000 13.005000 10.375000 13.305000 ;
      RECT  6.135000 14.205000 10.375000 14.505000 ;
      RECT  6.135000 15.405000 10.375000 15.705000 ;
      RECT  6.135000 16.605000 10.375000 16.905000 ;
      RECT  6.135000 17.835000 10.375000 18.135000 ;
      RECT  6.135000 19.035000 10.375000 19.335000 ;
      RECT  6.135000 20.235000 10.375000 20.535000 ;
      RECT  6.135000 21.435000 10.375000 21.735000 ;
      RECT 10.045000  0.565000 10.375000  1.465000 ;
      RECT 10.045000  1.765000 10.375000  2.665000 ;
      RECT 10.045000  2.965000 10.375000  3.865000 ;
      RECT 10.045000  4.165000 10.375000  5.065000 ;
      RECT 10.045000  5.365000 10.375000  6.295000 ;
      RECT 10.045000  6.595000 10.375000  7.495000 ;
      RECT 10.045000  7.795000 10.375000  8.695000 ;
      RECT 10.045000  8.995000 10.375000  9.895000 ;
      RECT 10.045000 10.195000 10.375000 11.095000 ;
      RECT 10.045000 12.105000 10.375000 13.005000 ;
      RECT 10.045000 13.305000 10.375000 14.205000 ;
      RECT 10.045000 14.505000 10.375000 15.405000 ;
      RECT 10.045000 15.705000 10.375000 16.605000 ;
      RECT 10.045000 16.905000 10.375000 17.835000 ;
      RECT 10.045000 18.135000 10.375000 19.035000 ;
      RECT 10.045000 19.335000 10.375000 20.235000 ;
      RECT 10.045000 20.535000 10.375000 21.435000 ;
      RECT 10.045000 21.735000 10.375000 22.635000 ;
      RECT 10.710000  0.140000 11.040000 23.220000 ;
      RECT 11.375000  0.235000 20.785000  0.565000 ;
      RECT 11.375000  0.565000 11.705000  1.465000 ;
      RECT 11.375000  1.465000 15.615000  1.765000 ;
      RECT 11.375000  1.765000 11.705000  2.665000 ;
      RECT 11.375000  2.665000 15.615000  2.965000 ;
      RECT 11.375000  2.965000 11.705000  3.865000 ;
      RECT 11.375000  3.865000 15.615000  4.165000 ;
      RECT 11.375000  4.165000 11.705000  5.065000 ;
      RECT 11.375000  5.065000 15.615000  5.365000 ;
      RECT 11.375000  5.365000 11.705000  6.295000 ;
      RECT 11.375000  6.295000 15.615000  6.595000 ;
      RECT 11.375000  6.595000 11.705000  7.495000 ;
      RECT 11.375000  7.495000 15.615000  7.795000 ;
      RECT 11.375000  7.795000 11.705000  8.695000 ;
      RECT 11.375000  8.695000 15.615000  8.995000 ;
      RECT 11.375000  8.995000 11.705000  9.895000 ;
      RECT 11.375000  9.895000 15.615000 10.195000 ;
      RECT 11.375000 10.195000 11.705000 11.095000 ;
      RECT 11.375000 11.095000 20.785000 11.425000 ;
      RECT 11.375000 11.775000 20.785000 12.105000 ;
      RECT 11.375000 12.105000 11.705000 13.005000 ;
      RECT 11.375000 13.005000 15.615000 13.305000 ;
      RECT 11.375000 13.305000 11.705000 14.205000 ;
      RECT 11.375000 14.205000 15.615000 14.505000 ;
      RECT 11.375000 14.505000 11.705000 15.405000 ;
      RECT 11.375000 15.405000 15.615000 15.705000 ;
      RECT 11.375000 15.705000 11.705000 16.605000 ;
      RECT 11.375000 16.605000 15.615000 16.905000 ;
      RECT 11.375000 16.905000 11.705000 17.835000 ;
      RECT 11.375000 17.835000 15.615000 18.135000 ;
      RECT 11.375000 18.135000 11.705000 19.035000 ;
      RECT 11.375000 19.035000 15.615000 19.335000 ;
      RECT 11.375000 19.335000 11.705000 20.235000 ;
      RECT 11.375000 20.235000 15.615000 20.535000 ;
      RECT 11.375000 20.535000 11.705000 21.435000 ;
      RECT 11.375000 21.435000 15.615000 21.735000 ;
      RECT 11.375000 21.735000 11.705000 22.635000 ;
      RECT 11.375000 22.635000 20.785000 22.965000 ;
      RECT 12.005000  0.865000 20.155000  1.165000 ;
      RECT 12.005000  2.065000 20.155000  2.365000 ;
      RECT 12.005000  3.265000 20.155000  3.565000 ;
      RECT 12.005000  4.465000 20.155000  4.765000 ;
      RECT 12.005000  5.665000 20.155000  5.995000 ;
      RECT 12.005000  6.895000 20.155000  7.195000 ;
      RECT 12.005000  8.095000 20.155000  8.395000 ;
      RECT 12.005000  9.295000 20.155000  9.595000 ;
      RECT 12.005000 10.495000 20.155000 10.795000 ;
      RECT 12.005000 12.405000 20.155000 12.705000 ;
      RECT 12.005000 13.605000 20.155000 13.905000 ;
      RECT 12.005000 14.805000 20.155000 15.105000 ;
      RECT 12.005000 16.005000 20.155000 16.305000 ;
      RECT 12.005000 17.205000 20.155000 17.535000 ;
      RECT 12.005000 18.435000 20.155000 18.735000 ;
      RECT 12.005000 19.635000 20.155000 19.935000 ;
      RECT 12.005000 20.835000 20.155000 21.135000 ;
      RECT 12.005000 22.035000 20.155000 22.335000 ;
      RECT 15.915000  1.165000 16.245000  2.065000 ;
      RECT 15.915000  2.365000 16.245000  3.265000 ;
      RECT 15.915000  3.565000 16.245000  4.465000 ;
      RECT 15.915000  4.765000 16.245000  5.665000 ;
      RECT 15.915000  5.995000 16.245000  6.895000 ;
      RECT 15.915000  7.195000 16.245000  8.095000 ;
      RECT 15.915000  8.395000 16.245000  9.295000 ;
      RECT 15.915000  9.595000 16.245000 10.495000 ;
      RECT 15.915000 12.705000 16.245000 13.605000 ;
      RECT 15.915000 13.905000 16.245000 14.805000 ;
      RECT 15.915000 15.105000 16.245000 16.005000 ;
      RECT 15.915000 16.305000 16.245000 17.205000 ;
      RECT 15.915000 17.535000 16.245000 18.435000 ;
      RECT 15.915000 18.735000 16.245000 19.635000 ;
      RECT 15.915000 19.935000 16.245000 20.835000 ;
      RECT 15.915000 21.135000 16.245000 22.035000 ;
      RECT 16.545000  1.465000 20.785000  1.765000 ;
      RECT 16.545000  2.665000 20.785000  2.965000 ;
      RECT 16.545000  3.865000 20.785000  4.165000 ;
      RECT 16.545000  5.065000 20.785000  5.365000 ;
      RECT 16.545000  6.295000 20.785000  6.595000 ;
      RECT 16.545000  7.495000 20.785000  7.795000 ;
      RECT 16.545000  8.695000 20.785000  8.995000 ;
      RECT 16.545000  9.895000 20.785000 10.195000 ;
      RECT 16.545000 13.005000 20.785000 13.305000 ;
      RECT 16.545000 14.205000 20.785000 14.505000 ;
      RECT 16.545000 15.405000 20.785000 15.705000 ;
      RECT 16.545000 16.605000 20.785000 16.905000 ;
      RECT 16.545000 17.835000 20.785000 18.135000 ;
      RECT 16.545000 19.035000 20.785000 19.335000 ;
      RECT 16.545000 20.235000 20.785000 20.535000 ;
      RECT 16.545000 21.435000 20.785000 21.735000 ;
      RECT 20.455000  0.565000 20.785000  1.465000 ;
      RECT 20.455000  1.765000 20.785000  2.665000 ;
      RECT 20.455000  2.965000 20.785000  3.865000 ;
      RECT 20.455000  4.165000 20.785000  5.065000 ;
      RECT 20.455000  5.365000 20.785000  6.295000 ;
      RECT 20.455000  6.595000 20.785000  7.495000 ;
      RECT 20.455000  7.795000 20.785000  8.695000 ;
      RECT 20.455000  8.995000 20.785000  9.895000 ;
      RECT 20.455000 10.195000 20.785000 11.095000 ;
      RECT 20.455000 12.105000 20.785000 13.005000 ;
      RECT 20.455000 13.305000 20.785000 14.205000 ;
      RECT 20.455000 14.505000 20.785000 15.405000 ;
      RECT 20.455000 15.705000 20.785000 16.605000 ;
      RECT 20.455000 16.905000 20.785000 17.835000 ;
      RECT 20.455000 18.135000 20.785000 19.035000 ;
      RECT 20.455000 19.335000 20.785000 20.235000 ;
      RECT 20.455000 20.535000 20.785000 21.435000 ;
      RECT 20.455000 21.735000 20.785000 22.635000 ;
      RECT 21.120000  0.140000 21.450000 23.220000 ;
    LAYER pwell ;
      RECT 9.960000 18.440000 10.720000 19.220000 ;
    LAYER via ;
      RECT  1.020000  1.960000  1.280000  2.220000 ;
      RECT  1.020000  2.280000  1.280000  2.540000 ;
      RECT  1.020000  2.600000  1.280000  2.860000 ;
      RECT  1.020000  2.920000  1.280000  3.180000 ;
      RECT  1.020000  3.240000  1.280000  3.500000 ;
      RECT  1.020000  3.560000  1.280000  3.820000 ;
      RECT  1.020000  3.880000  1.280000  4.140000 ;
      RECT  1.020000  4.200000  1.280000  4.460000 ;
      RECT  1.020000  4.520000  1.280000  4.780000 ;
      RECT  1.020000  4.840000  1.280000  5.100000 ;
      RECT  1.020000  5.160000  1.280000  5.420000 ;
      RECT  1.020000  6.270000  1.280000  6.530000 ;
      RECT  1.020000  6.590000  1.280000  6.850000 ;
      RECT  1.020000  6.910000  1.280000  7.170000 ;
      RECT  1.020000  7.230000  1.280000  7.490000 ;
      RECT  1.020000  7.550000  1.280000  7.810000 ;
      RECT  1.020000  7.870000  1.280000  8.130000 ;
      RECT  1.020000  8.190000  1.280000  8.450000 ;
      RECT  1.020000  8.510000  1.280000  8.770000 ;
      RECT  1.020000  8.830000  1.280000  9.090000 ;
      RECT  1.020000  9.150000  1.280000  9.410000 ;
      RECT  1.020000  9.470000  1.280000  9.730000 ;
      RECT  1.020000 13.500000  1.280000 13.760000 ;
      RECT  1.020000 13.820000  1.280000 14.080000 ;
      RECT  1.020000 14.140000  1.280000 14.400000 ;
      RECT  1.020000 14.460000  1.280000 14.720000 ;
      RECT  1.020000 14.780000  1.280000 15.040000 ;
      RECT  1.020000 15.100000  1.280000 15.360000 ;
      RECT  1.020000 15.420000  1.280000 15.680000 ;
      RECT  1.020000 15.740000  1.280000 16.000000 ;
      RECT  1.020000 16.060000  1.280000 16.320000 ;
      RECT  1.020000 16.380000  1.280000 16.640000 ;
      RECT  1.020000 16.700000  1.280000 16.960000 ;
      RECT  1.020000 17.810000  1.280000 18.070000 ;
      RECT  1.020000 18.130000  1.280000 18.390000 ;
      RECT  1.020000 18.450000  1.280000 18.710000 ;
      RECT  1.020000 18.770000  1.280000 19.030000 ;
      RECT  1.020000 19.090000  1.280000 19.350000 ;
      RECT  1.020000 19.410000  1.280000 19.670000 ;
      RECT  1.020000 19.730000  1.280000 19.990000 ;
      RECT  1.020000 20.050000  1.280000 20.310000 ;
      RECT  1.020000 20.370000  1.280000 20.630000 ;
      RECT  1.020000 20.690000  1.280000 20.950000 ;
      RECT  1.020000 21.010000  1.280000 21.270000 ;
      RECT  1.385000  0.355000  1.645000  0.615000 ;
      RECT  1.385000 11.205000  1.645000 11.465000 ;
      RECT  1.385000 11.895000  1.645000 12.155000 ;
      RECT  1.385000 22.745000  1.645000 23.005000 ;
      RECT  1.535000  5.535000  1.795000  5.795000 ;
      RECT  1.535000  5.895000  1.795000  6.155000 ;
      RECT  1.535000 17.075000  1.795000 17.335000 ;
      RECT  1.535000 17.435000  1.795000 17.695000 ;
      RECT  1.630000  1.425000  1.890000  1.685000 ;
      RECT  1.630000 10.005000  1.890000 10.265000 ;
      RECT  1.630000 12.965000  1.890000 13.225000 ;
      RECT  1.630000 21.545000  1.890000 21.805000 ;
      RECT  1.705000  0.355000  1.965000  0.615000 ;
      RECT  1.705000 11.205000  1.965000 11.465000 ;
      RECT  1.705000 11.895000  1.965000 12.155000 ;
      RECT  1.705000 22.745000  1.965000 23.005000 ;
      RECT  1.855000  5.535000  2.115000  5.795000 ;
      RECT  1.855000  5.895000  2.115000  6.155000 ;
      RECT  1.855000 17.075000  2.115000 17.335000 ;
      RECT  1.855000 17.435000  2.115000 17.695000 ;
      RECT  1.950000  1.425000  2.210000  1.685000 ;
      RECT  1.950000 10.005000  2.210000 10.265000 ;
      RECT  1.950000 12.965000  2.210000 13.225000 ;
      RECT  1.950000 21.545000  2.210000 21.805000 ;
      RECT  2.025000  0.355000  2.285000  0.615000 ;
      RECT  2.025000 11.205000  2.285000 11.465000 ;
      RECT  2.025000 11.895000  2.285000 12.155000 ;
      RECT  2.025000 22.745000  2.285000 23.005000 ;
      RECT  2.175000  5.535000  2.435000  5.795000 ;
      RECT  2.175000  5.895000  2.435000  6.155000 ;
      RECT  2.175000 17.075000  2.435000 17.335000 ;
      RECT  2.175000 17.435000  2.435000 17.695000 ;
      RECT  2.270000  1.425000  2.530000  1.685000 ;
      RECT  2.270000 10.005000  2.530000 10.265000 ;
      RECT  2.270000 12.965000  2.530000 13.225000 ;
      RECT  2.270000 21.545000  2.530000 21.805000 ;
      RECT  2.345000  0.355000  2.605000  0.615000 ;
      RECT  2.345000 11.205000  2.605000 11.465000 ;
      RECT  2.345000 11.895000  2.605000 12.155000 ;
      RECT  2.345000 22.745000  2.605000 23.005000 ;
      RECT  2.495000  5.535000  2.755000  5.795000 ;
      RECT  2.495000  5.895000  2.755000  6.155000 ;
      RECT  2.495000 17.075000  2.755000 17.335000 ;
      RECT  2.495000 17.435000  2.755000 17.695000 ;
      RECT  2.590000  1.425000  2.850000  1.685000 ;
      RECT  2.590000 10.005000  2.850000 10.265000 ;
      RECT  2.590000 12.965000  2.850000 13.225000 ;
      RECT  2.590000 21.545000  2.850000 21.805000 ;
      RECT  2.665000  0.355000  2.925000  0.615000 ;
      RECT  2.665000 11.205000  2.925000 11.465000 ;
      RECT  2.665000 11.895000  2.925000 12.155000 ;
      RECT  2.665000 22.745000  2.925000 23.005000 ;
      RECT  2.815000  5.535000  3.075000  5.795000 ;
      RECT  2.815000  5.895000  3.075000  6.155000 ;
      RECT  2.815000 17.075000  3.075000 17.335000 ;
      RECT  2.815000 17.435000  3.075000 17.695000 ;
      RECT  2.910000  1.425000  3.170000  1.685000 ;
      RECT  2.910000 10.005000  3.170000 10.265000 ;
      RECT  2.910000 12.965000  3.170000 13.225000 ;
      RECT  2.910000 21.545000  3.170000 21.805000 ;
      RECT  2.985000  0.355000  3.245000  0.615000 ;
      RECT  2.985000 11.205000  3.245000 11.465000 ;
      RECT  2.985000 11.895000  3.245000 12.155000 ;
      RECT  2.985000 22.745000  3.245000 23.005000 ;
      RECT  3.135000  5.535000  3.395000  5.795000 ;
      RECT  3.135000  5.895000  3.395000  6.155000 ;
      RECT  3.135000 17.075000  3.395000 17.335000 ;
      RECT  3.135000 17.435000  3.395000 17.695000 ;
      RECT  3.230000  1.425000  3.490000  1.685000 ;
      RECT  3.230000 10.005000  3.490000 10.265000 ;
      RECT  3.230000 12.965000  3.490000 13.225000 ;
      RECT  3.230000 21.545000  3.490000 21.805000 ;
      RECT  3.305000  0.355000  3.565000  0.615000 ;
      RECT  3.305000 11.205000  3.565000 11.465000 ;
      RECT  3.305000 11.895000  3.565000 12.155000 ;
      RECT  3.305000 22.745000  3.565000 23.005000 ;
      RECT  3.455000  5.535000  3.715000  5.795000 ;
      RECT  3.455000  5.895000  3.715000  6.155000 ;
      RECT  3.455000 17.075000  3.715000 17.335000 ;
      RECT  3.455000 17.435000  3.715000 17.695000 ;
      RECT  3.550000  1.425000  3.810000  1.685000 ;
      RECT  3.550000 10.005000  3.810000 10.265000 ;
      RECT  3.550000 12.965000  3.810000 13.225000 ;
      RECT  3.550000 21.545000  3.810000 21.805000 ;
      RECT  3.625000  0.355000  3.885000  0.615000 ;
      RECT  3.625000 11.205000  3.885000 11.465000 ;
      RECT  3.625000 11.895000  3.885000 12.155000 ;
      RECT  3.625000 22.745000  3.885000 23.005000 ;
      RECT  3.775000  5.535000  4.035000  5.795000 ;
      RECT  3.775000  5.895000  4.035000  6.155000 ;
      RECT  3.775000 17.075000  4.035000 17.335000 ;
      RECT  3.775000 17.435000  4.035000 17.695000 ;
      RECT  3.870000  1.425000  4.130000  1.685000 ;
      RECT  3.870000 10.005000  4.130000 10.265000 ;
      RECT  3.870000 12.965000  4.130000 13.225000 ;
      RECT  3.870000 21.545000  4.130000 21.805000 ;
      RECT  3.945000  0.355000  4.205000  0.615000 ;
      RECT  3.945000 11.205000  4.205000 11.465000 ;
      RECT  3.945000 11.895000  4.205000 12.155000 ;
      RECT  3.945000 22.745000  4.205000 23.005000 ;
      RECT  4.095000  5.535000  4.355000  5.795000 ;
      RECT  4.095000  5.895000  4.355000  6.155000 ;
      RECT  4.095000 17.075000  4.355000 17.335000 ;
      RECT  4.095000 17.435000  4.355000 17.695000 ;
      RECT  4.190000  1.425000  4.450000  1.685000 ;
      RECT  4.190000 10.005000  4.450000 10.265000 ;
      RECT  4.190000 12.965000  4.450000 13.225000 ;
      RECT  4.190000 21.545000  4.450000 21.805000 ;
      RECT  4.265000  0.355000  4.525000  0.615000 ;
      RECT  4.265000 11.205000  4.525000 11.465000 ;
      RECT  4.265000 11.895000  4.525000 12.155000 ;
      RECT  4.265000 22.745000  4.525000 23.005000 ;
      RECT  4.415000  5.535000  4.675000  5.795000 ;
      RECT  4.415000  5.895000  4.675000  6.155000 ;
      RECT  4.415000 17.075000  4.675000 17.335000 ;
      RECT  4.415000 17.435000  4.675000 17.695000 ;
      RECT  4.510000  1.425000  4.770000  1.685000 ;
      RECT  4.510000 10.005000  4.770000 10.265000 ;
      RECT  4.510000 12.965000  4.770000 13.225000 ;
      RECT  4.510000 21.545000  4.770000 21.805000 ;
      RECT  4.585000  0.355000  4.845000  0.615000 ;
      RECT  4.585000 11.205000  4.845000 11.465000 ;
      RECT  4.585000 11.895000  4.845000 12.155000 ;
      RECT  4.585000 22.745000  4.845000 23.005000 ;
      RECT  4.735000  5.535000  4.995000  5.795000 ;
      RECT  4.735000  5.895000  4.995000  6.155000 ;
      RECT  4.735000 17.075000  4.995000 17.335000 ;
      RECT  4.735000 17.435000  4.995000 17.695000 ;
      RECT  4.830000  1.425000  5.090000  1.685000 ;
      RECT  4.830000 10.005000  5.090000 10.265000 ;
      RECT  4.830000 12.965000  5.090000 13.225000 ;
      RECT  4.830000 21.545000  5.090000 21.805000 ;
      RECT  4.905000  0.355000  5.165000  0.615000 ;
      RECT  4.905000 11.205000  5.165000 11.465000 ;
      RECT  4.905000 11.895000  5.165000 12.155000 ;
      RECT  4.905000 22.745000  5.165000 23.005000 ;
      RECT  5.055000  5.535000  5.315000  5.795000 ;
      RECT  5.055000  5.895000  5.315000  6.155000 ;
      RECT  5.055000 17.075000  5.315000 17.335000 ;
      RECT  5.055000 17.435000  5.315000 17.695000 ;
      RECT  5.225000  0.355000  5.485000  0.615000 ;
      RECT  5.225000 11.205000  5.485000 11.465000 ;
      RECT  5.225000 11.895000  5.485000 12.155000 ;
      RECT  5.225000 22.745000  5.485000 23.005000 ;
      RECT  5.290000  1.960000  5.550000  2.220000 ;
      RECT  5.290000  2.280000  5.550000  2.540000 ;
      RECT  5.290000  2.600000  5.550000  2.860000 ;
      RECT  5.290000  2.920000  5.550000  3.180000 ;
      RECT  5.290000  3.240000  5.550000  3.500000 ;
      RECT  5.290000  3.560000  5.550000  3.820000 ;
      RECT  5.290000  3.880000  5.550000  4.140000 ;
      RECT  5.290000  4.200000  5.550000  4.460000 ;
      RECT  5.290000  4.520000  5.550000  4.780000 ;
      RECT  5.290000  4.840000  5.550000  5.100000 ;
      RECT  5.290000  5.160000  5.550000  5.420000 ;
      RECT  5.290000  6.270000  5.550000  6.530000 ;
      RECT  5.290000  6.590000  5.550000  6.850000 ;
      RECT  5.290000  6.910000  5.550000  7.170000 ;
      RECT  5.290000  7.230000  5.550000  7.490000 ;
      RECT  5.290000  7.550000  5.550000  7.810000 ;
      RECT  5.290000  7.870000  5.550000  8.130000 ;
      RECT  5.290000  8.190000  5.550000  8.450000 ;
      RECT  5.290000  8.510000  5.550000  8.770000 ;
      RECT  5.290000  8.830000  5.550000  9.090000 ;
      RECT  5.290000  9.150000  5.550000  9.410000 ;
      RECT  5.290000  9.470000  5.550000  9.730000 ;
      RECT  5.290000 13.500000  5.550000 13.760000 ;
      RECT  5.290000 13.820000  5.550000 14.080000 ;
      RECT  5.290000 14.140000  5.550000 14.400000 ;
      RECT  5.290000 14.460000  5.550000 14.720000 ;
      RECT  5.290000 14.780000  5.550000 15.040000 ;
      RECT  5.290000 15.100000  5.550000 15.360000 ;
      RECT  5.290000 15.420000  5.550000 15.680000 ;
      RECT  5.290000 15.740000  5.550000 16.000000 ;
      RECT  5.290000 16.060000  5.550000 16.320000 ;
      RECT  5.290000 16.380000  5.550000 16.640000 ;
      RECT  5.290000 16.700000  5.550000 16.960000 ;
      RECT  5.290000 17.810000  5.550000 18.070000 ;
      RECT  5.290000 18.130000  5.550000 18.390000 ;
      RECT  5.290000 18.450000  5.550000 18.710000 ;
      RECT  5.290000 18.770000  5.550000 19.030000 ;
      RECT  5.290000 19.090000  5.550000 19.350000 ;
      RECT  5.290000 19.410000  5.550000 19.670000 ;
      RECT  5.290000 19.730000  5.550000 19.990000 ;
      RECT  5.290000 20.050000  5.550000 20.310000 ;
      RECT  5.290000 20.370000  5.550000 20.630000 ;
      RECT  5.290000 20.690000  5.550000 20.950000 ;
      RECT  5.290000 21.010000  5.550000 21.270000 ;
      RECT  5.545000  0.355000  5.805000  0.615000 ;
      RECT  5.545000 11.205000  5.805000 11.465000 ;
      RECT  5.545000 11.895000  5.805000 12.155000 ;
      RECT  5.545000 22.745000  5.805000 23.005000 ;
      RECT  5.790000  1.960000  6.050000  2.220000 ;
      RECT  5.790000  2.280000  6.050000  2.540000 ;
      RECT  5.790000  2.600000  6.050000  2.860000 ;
      RECT  5.790000  2.920000  6.050000  3.180000 ;
      RECT  5.790000  3.240000  6.050000  3.500000 ;
      RECT  5.790000  3.560000  6.050000  3.820000 ;
      RECT  5.790000  3.880000  6.050000  4.140000 ;
      RECT  5.790000  4.200000  6.050000  4.460000 ;
      RECT  5.790000  4.520000  6.050000  4.780000 ;
      RECT  5.790000  4.840000  6.050000  5.100000 ;
      RECT  5.790000  5.160000  6.050000  5.420000 ;
      RECT  5.790000  6.270000  6.050000  6.530000 ;
      RECT  5.790000  6.590000  6.050000  6.850000 ;
      RECT  5.790000  6.910000  6.050000  7.170000 ;
      RECT  5.790000  7.230000  6.050000  7.490000 ;
      RECT  5.790000  7.550000  6.050000  7.810000 ;
      RECT  5.790000  7.870000  6.050000  8.130000 ;
      RECT  5.790000  8.190000  6.050000  8.450000 ;
      RECT  5.790000  8.510000  6.050000  8.770000 ;
      RECT  5.790000  8.830000  6.050000  9.090000 ;
      RECT  5.790000  9.150000  6.050000  9.410000 ;
      RECT  5.790000  9.470000  6.050000  9.730000 ;
      RECT  5.790000 13.500000  6.050000 13.760000 ;
      RECT  5.790000 13.820000  6.050000 14.080000 ;
      RECT  5.790000 14.140000  6.050000 14.400000 ;
      RECT  5.790000 14.460000  6.050000 14.720000 ;
      RECT  5.790000 14.780000  6.050000 15.040000 ;
      RECT  5.790000 15.100000  6.050000 15.360000 ;
      RECT  5.790000 15.420000  6.050000 15.680000 ;
      RECT  5.790000 15.740000  6.050000 16.000000 ;
      RECT  5.790000 16.060000  6.050000 16.320000 ;
      RECT  5.790000 16.380000  6.050000 16.640000 ;
      RECT  5.790000 16.700000  6.050000 16.960000 ;
      RECT  5.790000 17.810000  6.050000 18.070000 ;
      RECT  5.790000 18.130000  6.050000 18.390000 ;
      RECT  5.790000 18.450000  6.050000 18.710000 ;
      RECT  5.790000 18.770000  6.050000 19.030000 ;
      RECT  5.790000 19.090000  6.050000 19.350000 ;
      RECT  5.790000 19.410000  6.050000 19.670000 ;
      RECT  5.790000 19.730000  6.050000 19.990000 ;
      RECT  5.790000 20.050000  6.050000 20.310000 ;
      RECT  5.790000 20.370000  6.050000 20.630000 ;
      RECT  5.790000 20.690000  6.050000 20.950000 ;
      RECT  5.790000 21.010000  6.050000 21.270000 ;
      RECT  5.865000  0.355000  6.125000  0.615000 ;
      RECT  5.865000 11.205000  6.125000 11.465000 ;
      RECT  5.865000 11.895000  6.125000 12.155000 ;
      RECT  5.865000 22.745000  6.125000 23.005000 ;
      RECT  6.025000  5.535000  6.285000  5.795000 ;
      RECT  6.025000  5.895000  6.285000  6.155000 ;
      RECT  6.025000 17.075000  6.285000 17.335000 ;
      RECT  6.025000 17.435000  6.285000 17.695000 ;
      RECT  6.185000  0.355000  6.445000  0.615000 ;
      RECT  6.185000 11.205000  6.445000 11.465000 ;
      RECT  6.185000 11.895000  6.445000 12.155000 ;
      RECT  6.185000 22.745000  6.445000 23.005000 ;
      RECT  6.250000  1.425000  6.510000  1.685000 ;
      RECT  6.250000 10.005000  6.510000 10.265000 ;
      RECT  6.250000 12.965000  6.510000 13.225000 ;
      RECT  6.250000 21.545000  6.510000 21.805000 ;
      RECT  6.345000  5.535000  6.605000  5.795000 ;
      RECT  6.345000  5.895000  6.605000  6.155000 ;
      RECT  6.345000 17.075000  6.605000 17.335000 ;
      RECT  6.345000 17.435000  6.605000 17.695000 ;
      RECT  6.505000  0.355000  6.765000  0.615000 ;
      RECT  6.505000 11.205000  6.765000 11.465000 ;
      RECT  6.505000 11.895000  6.765000 12.155000 ;
      RECT  6.505000 22.745000  6.765000 23.005000 ;
      RECT  6.570000  1.425000  6.830000  1.685000 ;
      RECT  6.570000 10.005000  6.830000 10.265000 ;
      RECT  6.570000 12.965000  6.830000 13.225000 ;
      RECT  6.570000 21.545000  6.830000 21.805000 ;
      RECT  6.665000  5.535000  6.925000  5.795000 ;
      RECT  6.665000  5.895000  6.925000  6.155000 ;
      RECT  6.665000 17.075000  6.925000 17.335000 ;
      RECT  6.665000 17.435000  6.925000 17.695000 ;
      RECT  6.825000  0.355000  7.085000  0.615000 ;
      RECT  6.825000 11.205000  7.085000 11.465000 ;
      RECT  6.825000 11.895000  7.085000 12.155000 ;
      RECT  6.825000 22.745000  7.085000 23.005000 ;
      RECT  6.890000  1.425000  7.150000  1.685000 ;
      RECT  6.890000 10.005000  7.150000 10.265000 ;
      RECT  6.890000 12.965000  7.150000 13.225000 ;
      RECT  6.890000 21.545000  7.150000 21.805000 ;
      RECT  6.985000  5.535000  7.245000  5.795000 ;
      RECT  6.985000  5.895000  7.245000  6.155000 ;
      RECT  6.985000 17.075000  7.245000 17.335000 ;
      RECT  6.985000 17.435000  7.245000 17.695000 ;
      RECT  7.145000  0.355000  7.405000  0.615000 ;
      RECT  7.145000 11.205000  7.405000 11.465000 ;
      RECT  7.145000 11.895000  7.405000 12.155000 ;
      RECT  7.145000 22.745000  7.405000 23.005000 ;
      RECT  7.210000  1.425000  7.470000  1.685000 ;
      RECT  7.210000 10.005000  7.470000 10.265000 ;
      RECT  7.210000 12.965000  7.470000 13.225000 ;
      RECT  7.210000 21.545000  7.470000 21.805000 ;
      RECT  7.305000  5.535000  7.565000  5.795000 ;
      RECT  7.305000  5.895000  7.565000  6.155000 ;
      RECT  7.305000 17.075000  7.565000 17.335000 ;
      RECT  7.305000 17.435000  7.565000 17.695000 ;
      RECT  7.465000  0.355000  7.725000  0.615000 ;
      RECT  7.465000 11.205000  7.725000 11.465000 ;
      RECT  7.465000 11.895000  7.725000 12.155000 ;
      RECT  7.465000 22.745000  7.725000 23.005000 ;
      RECT  7.530000  1.425000  7.790000  1.685000 ;
      RECT  7.530000 10.005000  7.790000 10.265000 ;
      RECT  7.530000 12.965000  7.790000 13.225000 ;
      RECT  7.530000 21.545000  7.790000 21.805000 ;
      RECT  7.625000  5.535000  7.885000  5.795000 ;
      RECT  7.625000  5.895000  7.885000  6.155000 ;
      RECT  7.625000 17.075000  7.885000 17.335000 ;
      RECT  7.625000 17.435000  7.885000 17.695000 ;
      RECT  7.785000  0.355000  8.045000  0.615000 ;
      RECT  7.785000 11.205000  8.045000 11.465000 ;
      RECT  7.785000 11.895000  8.045000 12.155000 ;
      RECT  7.785000 22.745000  8.045000 23.005000 ;
      RECT  7.850000  1.425000  8.110000  1.685000 ;
      RECT  7.850000 10.005000  8.110000 10.265000 ;
      RECT  7.850000 12.965000  8.110000 13.225000 ;
      RECT  7.850000 21.545000  8.110000 21.805000 ;
      RECT  7.945000  5.535000  8.205000  5.795000 ;
      RECT  7.945000  5.895000  8.205000  6.155000 ;
      RECT  7.945000 17.075000  8.205000 17.335000 ;
      RECT  7.945000 17.435000  8.205000 17.695000 ;
      RECT  8.105000  0.355000  8.365000  0.615000 ;
      RECT  8.105000 11.205000  8.365000 11.465000 ;
      RECT  8.105000 11.895000  8.365000 12.155000 ;
      RECT  8.105000 22.745000  8.365000 23.005000 ;
      RECT  8.170000  1.425000  8.430000  1.685000 ;
      RECT  8.170000 10.005000  8.430000 10.265000 ;
      RECT  8.170000 12.965000  8.430000 13.225000 ;
      RECT  8.170000 21.545000  8.430000 21.805000 ;
      RECT  8.265000  5.535000  8.525000  5.795000 ;
      RECT  8.265000  5.895000  8.525000  6.155000 ;
      RECT  8.265000 17.075000  8.525000 17.335000 ;
      RECT  8.265000 17.435000  8.525000 17.695000 ;
      RECT  8.425000  0.355000  8.685000  0.615000 ;
      RECT  8.425000 11.205000  8.685000 11.465000 ;
      RECT  8.425000 11.895000  8.685000 12.155000 ;
      RECT  8.425000 22.745000  8.685000 23.005000 ;
      RECT  8.490000  1.425000  8.750000  1.685000 ;
      RECT  8.490000 10.005000  8.750000 10.265000 ;
      RECT  8.490000 12.965000  8.750000 13.225000 ;
      RECT  8.490000 21.545000  8.750000 21.805000 ;
      RECT  8.585000  5.535000  8.845000  5.795000 ;
      RECT  8.585000  5.895000  8.845000  6.155000 ;
      RECT  8.585000 17.075000  8.845000 17.335000 ;
      RECT  8.585000 17.435000  8.845000 17.695000 ;
      RECT  8.745000  0.355000  9.005000  0.615000 ;
      RECT  8.745000 11.205000  9.005000 11.465000 ;
      RECT  8.745000 11.895000  9.005000 12.155000 ;
      RECT  8.745000 22.745000  9.005000 23.005000 ;
      RECT  8.810000  1.425000  9.070000  1.685000 ;
      RECT  8.810000 10.005000  9.070000 10.265000 ;
      RECT  8.810000 12.965000  9.070000 13.225000 ;
      RECT  8.810000 21.545000  9.070000 21.805000 ;
      RECT  8.905000  5.535000  9.165000  5.795000 ;
      RECT  8.905000  5.895000  9.165000  6.155000 ;
      RECT  8.905000 17.075000  9.165000 17.335000 ;
      RECT  8.905000 17.435000  9.165000 17.695000 ;
      RECT  9.065000  0.355000  9.325000  0.615000 ;
      RECT  9.065000 11.205000  9.325000 11.465000 ;
      RECT  9.065000 11.895000  9.325000 12.155000 ;
      RECT  9.065000 22.745000  9.325000 23.005000 ;
      RECT  9.130000  1.425000  9.390000  1.685000 ;
      RECT  9.130000 10.005000  9.390000 10.265000 ;
      RECT  9.130000 12.965000  9.390000 13.225000 ;
      RECT  9.130000 21.545000  9.390000 21.805000 ;
      RECT  9.225000  5.535000  9.485000  5.795000 ;
      RECT  9.225000  5.895000  9.485000  6.155000 ;
      RECT  9.225000 17.075000  9.485000 17.335000 ;
      RECT  9.225000 17.435000  9.485000 17.695000 ;
      RECT  9.385000  0.355000  9.645000  0.615000 ;
      RECT  9.385000 11.205000  9.645000 11.465000 ;
      RECT  9.385000 11.895000  9.645000 12.155000 ;
      RECT  9.385000 22.745000  9.645000 23.005000 ;
      RECT  9.450000  1.425000  9.710000  1.685000 ;
      RECT  9.450000 10.005000  9.710000 10.265000 ;
      RECT  9.450000 12.965000  9.710000 13.225000 ;
      RECT  9.450000 21.545000  9.710000 21.805000 ;
      RECT  9.545000  5.535000  9.805000  5.795000 ;
      RECT  9.545000  5.895000  9.805000  6.155000 ;
      RECT  9.545000 17.075000  9.805000 17.335000 ;
      RECT  9.545000 17.435000  9.805000 17.695000 ;
      RECT 10.060000  1.960000 10.320000  2.220000 ;
      RECT 10.060000  2.280000 10.320000  2.540000 ;
      RECT 10.060000  2.600000 10.320000  2.860000 ;
      RECT 10.060000  2.920000 10.320000  3.180000 ;
      RECT 10.060000  3.240000 10.320000  3.500000 ;
      RECT 10.060000  3.560000 10.320000  3.820000 ;
      RECT 10.060000  3.880000 10.320000  4.140000 ;
      RECT 10.060000  4.200000 10.320000  4.460000 ;
      RECT 10.060000  4.520000 10.320000  4.780000 ;
      RECT 10.060000  4.840000 10.320000  5.100000 ;
      RECT 10.060000  5.160000 10.320000  5.420000 ;
      RECT 10.060000  6.270000 10.320000  6.530000 ;
      RECT 10.060000  6.590000 10.320000  6.850000 ;
      RECT 10.060000  6.910000 10.320000  7.170000 ;
      RECT 10.060000  7.230000 10.320000  7.490000 ;
      RECT 10.060000  7.550000 10.320000  7.810000 ;
      RECT 10.060000  7.870000 10.320000  8.130000 ;
      RECT 10.060000  8.190000 10.320000  8.450000 ;
      RECT 10.060000  8.510000 10.320000  8.770000 ;
      RECT 10.060000  8.830000 10.320000  9.090000 ;
      RECT 10.060000  9.150000 10.320000  9.410000 ;
      RECT 10.060000  9.470000 10.320000  9.730000 ;
      RECT 10.060000 13.500000 10.320000 13.760000 ;
      RECT 10.060000 13.820000 10.320000 14.080000 ;
      RECT 10.060000 14.140000 10.320000 14.400000 ;
      RECT 10.060000 14.460000 10.320000 14.720000 ;
      RECT 10.060000 14.780000 10.320000 15.040000 ;
      RECT 10.060000 15.100000 10.320000 15.360000 ;
      RECT 10.060000 15.420000 10.320000 15.680000 ;
      RECT 10.060000 15.740000 10.320000 16.000000 ;
      RECT 10.060000 16.060000 10.320000 16.320000 ;
      RECT 10.060000 16.380000 10.320000 16.640000 ;
      RECT 10.060000 16.700000 10.320000 16.960000 ;
      RECT 10.060000 17.810000 10.320000 18.070000 ;
      RECT 10.060000 18.130000 10.320000 18.390000 ;
      RECT 10.060000 18.450000 10.320000 18.710000 ;
      RECT 10.060000 18.770000 10.320000 19.030000 ;
      RECT 10.060000 19.090000 10.320000 19.350000 ;
      RECT 10.060000 19.410000 10.320000 19.670000 ;
      RECT 10.060000 19.730000 10.320000 19.990000 ;
      RECT 10.060000 20.050000 10.320000 20.310000 ;
      RECT 10.060000 20.370000 10.320000 20.630000 ;
      RECT 10.060000 20.690000 10.320000 20.950000 ;
      RECT 10.060000 21.010000 10.320000 21.270000 ;
      RECT 11.430000  1.960000 11.690000  2.220000 ;
      RECT 11.430000  2.280000 11.690000  2.540000 ;
      RECT 11.430000  2.600000 11.690000  2.860000 ;
      RECT 11.430000  2.920000 11.690000  3.180000 ;
      RECT 11.430000  3.240000 11.690000  3.500000 ;
      RECT 11.430000  3.560000 11.690000  3.820000 ;
      RECT 11.430000  3.880000 11.690000  4.140000 ;
      RECT 11.430000  4.200000 11.690000  4.460000 ;
      RECT 11.430000  4.520000 11.690000  4.780000 ;
      RECT 11.430000  4.840000 11.690000  5.100000 ;
      RECT 11.430000  5.160000 11.690000  5.420000 ;
      RECT 11.430000  6.270000 11.690000  6.530000 ;
      RECT 11.430000  6.590000 11.690000  6.850000 ;
      RECT 11.430000  6.910000 11.690000  7.170000 ;
      RECT 11.430000  7.230000 11.690000  7.490000 ;
      RECT 11.430000  7.550000 11.690000  7.810000 ;
      RECT 11.430000  7.870000 11.690000  8.130000 ;
      RECT 11.430000  8.190000 11.690000  8.450000 ;
      RECT 11.430000  8.510000 11.690000  8.770000 ;
      RECT 11.430000  8.830000 11.690000  9.090000 ;
      RECT 11.430000  9.150000 11.690000  9.410000 ;
      RECT 11.430000  9.470000 11.690000  9.730000 ;
      RECT 11.430000 13.500000 11.690000 13.760000 ;
      RECT 11.430000 13.820000 11.690000 14.080000 ;
      RECT 11.430000 14.140000 11.690000 14.400000 ;
      RECT 11.430000 14.460000 11.690000 14.720000 ;
      RECT 11.430000 14.780000 11.690000 15.040000 ;
      RECT 11.430000 15.100000 11.690000 15.360000 ;
      RECT 11.430000 15.420000 11.690000 15.680000 ;
      RECT 11.430000 15.740000 11.690000 16.000000 ;
      RECT 11.430000 16.060000 11.690000 16.320000 ;
      RECT 11.430000 16.380000 11.690000 16.640000 ;
      RECT 11.430000 16.700000 11.690000 16.960000 ;
      RECT 11.430000 17.810000 11.690000 18.070000 ;
      RECT 11.430000 18.130000 11.690000 18.390000 ;
      RECT 11.430000 18.450000 11.690000 18.710000 ;
      RECT 11.430000 18.770000 11.690000 19.030000 ;
      RECT 11.430000 19.090000 11.690000 19.350000 ;
      RECT 11.430000 19.410000 11.690000 19.670000 ;
      RECT 11.430000 19.730000 11.690000 19.990000 ;
      RECT 11.430000 20.050000 11.690000 20.310000 ;
      RECT 11.430000 20.370000 11.690000 20.630000 ;
      RECT 11.430000 20.690000 11.690000 20.950000 ;
      RECT 11.430000 21.010000 11.690000 21.270000 ;
      RECT 11.795000  0.355000 12.055000  0.615000 ;
      RECT 11.795000 11.205000 12.055000 11.465000 ;
      RECT 11.795000 11.895000 12.055000 12.155000 ;
      RECT 11.795000 22.745000 12.055000 23.005000 ;
      RECT 11.945000  5.535000 12.205000  5.795000 ;
      RECT 11.945000  5.895000 12.205000  6.155000 ;
      RECT 11.945000 17.075000 12.205000 17.335000 ;
      RECT 11.945000 17.435000 12.205000 17.695000 ;
      RECT 12.040000  1.425000 12.300000  1.685000 ;
      RECT 12.040000 10.005000 12.300000 10.265000 ;
      RECT 12.040000 12.965000 12.300000 13.225000 ;
      RECT 12.040000 21.545000 12.300000 21.805000 ;
      RECT 12.115000  0.355000 12.375000  0.615000 ;
      RECT 12.115000 11.205000 12.375000 11.465000 ;
      RECT 12.115000 11.895000 12.375000 12.155000 ;
      RECT 12.115000 22.745000 12.375000 23.005000 ;
      RECT 12.265000  5.535000 12.525000  5.795000 ;
      RECT 12.265000  5.895000 12.525000  6.155000 ;
      RECT 12.265000 17.075000 12.525000 17.335000 ;
      RECT 12.265000 17.435000 12.525000 17.695000 ;
      RECT 12.360000  1.425000 12.620000  1.685000 ;
      RECT 12.360000 10.005000 12.620000 10.265000 ;
      RECT 12.360000 12.965000 12.620000 13.225000 ;
      RECT 12.360000 21.545000 12.620000 21.805000 ;
      RECT 12.435000  0.355000 12.695000  0.615000 ;
      RECT 12.435000 11.205000 12.695000 11.465000 ;
      RECT 12.435000 11.895000 12.695000 12.155000 ;
      RECT 12.435000 22.745000 12.695000 23.005000 ;
      RECT 12.585000  5.535000 12.845000  5.795000 ;
      RECT 12.585000  5.895000 12.845000  6.155000 ;
      RECT 12.585000 17.075000 12.845000 17.335000 ;
      RECT 12.585000 17.435000 12.845000 17.695000 ;
      RECT 12.680000  1.425000 12.940000  1.685000 ;
      RECT 12.680000 10.005000 12.940000 10.265000 ;
      RECT 12.680000 12.965000 12.940000 13.225000 ;
      RECT 12.680000 21.545000 12.940000 21.805000 ;
      RECT 12.755000  0.355000 13.015000  0.615000 ;
      RECT 12.755000 11.205000 13.015000 11.465000 ;
      RECT 12.755000 11.895000 13.015000 12.155000 ;
      RECT 12.755000 22.745000 13.015000 23.005000 ;
      RECT 12.905000  5.535000 13.165000  5.795000 ;
      RECT 12.905000  5.895000 13.165000  6.155000 ;
      RECT 12.905000 17.075000 13.165000 17.335000 ;
      RECT 12.905000 17.435000 13.165000 17.695000 ;
      RECT 13.000000  1.425000 13.260000  1.685000 ;
      RECT 13.000000 10.005000 13.260000 10.265000 ;
      RECT 13.000000 12.965000 13.260000 13.225000 ;
      RECT 13.000000 21.545000 13.260000 21.805000 ;
      RECT 13.075000  0.355000 13.335000  0.615000 ;
      RECT 13.075000 11.205000 13.335000 11.465000 ;
      RECT 13.075000 11.895000 13.335000 12.155000 ;
      RECT 13.075000 22.745000 13.335000 23.005000 ;
      RECT 13.225000  5.535000 13.485000  5.795000 ;
      RECT 13.225000  5.895000 13.485000  6.155000 ;
      RECT 13.225000 17.075000 13.485000 17.335000 ;
      RECT 13.225000 17.435000 13.485000 17.695000 ;
      RECT 13.320000  1.425000 13.580000  1.685000 ;
      RECT 13.320000 10.005000 13.580000 10.265000 ;
      RECT 13.320000 12.965000 13.580000 13.225000 ;
      RECT 13.320000 21.545000 13.580000 21.805000 ;
      RECT 13.395000  0.355000 13.655000  0.615000 ;
      RECT 13.395000 11.205000 13.655000 11.465000 ;
      RECT 13.395000 11.895000 13.655000 12.155000 ;
      RECT 13.395000 22.745000 13.655000 23.005000 ;
      RECT 13.545000  5.535000 13.805000  5.795000 ;
      RECT 13.545000  5.895000 13.805000  6.155000 ;
      RECT 13.545000 17.075000 13.805000 17.335000 ;
      RECT 13.545000 17.435000 13.805000 17.695000 ;
      RECT 13.640000  1.425000 13.900000  1.685000 ;
      RECT 13.640000 10.005000 13.900000 10.265000 ;
      RECT 13.640000 12.965000 13.900000 13.225000 ;
      RECT 13.640000 21.545000 13.900000 21.805000 ;
      RECT 13.715000  0.355000 13.975000  0.615000 ;
      RECT 13.715000 11.205000 13.975000 11.465000 ;
      RECT 13.715000 11.895000 13.975000 12.155000 ;
      RECT 13.715000 22.745000 13.975000 23.005000 ;
      RECT 13.865000  5.535000 14.125000  5.795000 ;
      RECT 13.865000  5.895000 14.125000  6.155000 ;
      RECT 13.865000 17.075000 14.125000 17.335000 ;
      RECT 13.865000 17.435000 14.125000 17.695000 ;
      RECT 13.960000  1.425000 14.220000  1.685000 ;
      RECT 13.960000 10.005000 14.220000 10.265000 ;
      RECT 13.960000 12.965000 14.220000 13.225000 ;
      RECT 13.960000 21.545000 14.220000 21.805000 ;
      RECT 14.035000  0.355000 14.295000  0.615000 ;
      RECT 14.035000 11.205000 14.295000 11.465000 ;
      RECT 14.035000 11.895000 14.295000 12.155000 ;
      RECT 14.035000 22.745000 14.295000 23.005000 ;
      RECT 14.185000  5.535000 14.445000  5.795000 ;
      RECT 14.185000  5.895000 14.445000  6.155000 ;
      RECT 14.185000 17.075000 14.445000 17.335000 ;
      RECT 14.185000 17.435000 14.445000 17.695000 ;
      RECT 14.280000  1.425000 14.540000  1.685000 ;
      RECT 14.280000 10.005000 14.540000 10.265000 ;
      RECT 14.280000 12.965000 14.540000 13.225000 ;
      RECT 14.280000 21.545000 14.540000 21.805000 ;
      RECT 14.355000  0.355000 14.615000  0.615000 ;
      RECT 14.355000 11.205000 14.615000 11.465000 ;
      RECT 14.355000 11.895000 14.615000 12.155000 ;
      RECT 14.355000 22.745000 14.615000 23.005000 ;
      RECT 14.505000  5.535000 14.765000  5.795000 ;
      RECT 14.505000  5.895000 14.765000  6.155000 ;
      RECT 14.505000 17.075000 14.765000 17.335000 ;
      RECT 14.505000 17.435000 14.765000 17.695000 ;
      RECT 14.600000  1.425000 14.860000  1.685000 ;
      RECT 14.600000 10.005000 14.860000 10.265000 ;
      RECT 14.600000 12.965000 14.860000 13.225000 ;
      RECT 14.600000 21.545000 14.860000 21.805000 ;
      RECT 14.675000  0.355000 14.935000  0.615000 ;
      RECT 14.675000 11.205000 14.935000 11.465000 ;
      RECT 14.675000 11.895000 14.935000 12.155000 ;
      RECT 14.675000 22.745000 14.935000 23.005000 ;
      RECT 14.825000  5.535000 15.085000  5.795000 ;
      RECT 14.825000  5.895000 15.085000  6.155000 ;
      RECT 14.825000 17.075000 15.085000 17.335000 ;
      RECT 14.825000 17.435000 15.085000 17.695000 ;
      RECT 14.920000  1.425000 15.180000  1.685000 ;
      RECT 14.920000 10.005000 15.180000 10.265000 ;
      RECT 14.920000 12.965000 15.180000 13.225000 ;
      RECT 14.920000 21.545000 15.180000 21.805000 ;
      RECT 14.995000  0.355000 15.255000  0.615000 ;
      RECT 14.995000 11.205000 15.255000 11.465000 ;
      RECT 14.995000 11.895000 15.255000 12.155000 ;
      RECT 14.995000 22.745000 15.255000 23.005000 ;
      RECT 15.145000  5.535000 15.405000  5.795000 ;
      RECT 15.145000  5.895000 15.405000  6.155000 ;
      RECT 15.145000 17.075000 15.405000 17.335000 ;
      RECT 15.145000 17.435000 15.405000 17.695000 ;
      RECT 15.240000  1.425000 15.500000  1.685000 ;
      RECT 15.240000 10.005000 15.500000 10.265000 ;
      RECT 15.240000 12.965000 15.500000 13.225000 ;
      RECT 15.240000 21.545000 15.500000 21.805000 ;
      RECT 15.315000  0.355000 15.575000  0.615000 ;
      RECT 15.315000 11.205000 15.575000 11.465000 ;
      RECT 15.315000 11.895000 15.575000 12.155000 ;
      RECT 15.315000 22.745000 15.575000 23.005000 ;
      RECT 15.465000  5.535000 15.725000  5.795000 ;
      RECT 15.465000  5.895000 15.725000  6.155000 ;
      RECT 15.465000 17.075000 15.725000 17.335000 ;
      RECT 15.465000 17.435000 15.725000 17.695000 ;
      RECT 15.635000  0.355000 15.895000  0.615000 ;
      RECT 15.635000 11.205000 15.895000 11.465000 ;
      RECT 15.635000 11.895000 15.895000 12.155000 ;
      RECT 15.635000 22.745000 15.895000 23.005000 ;
      RECT 15.700000  1.960000 15.960000  2.220000 ;
      RECT 15.700000  2.280000 15.960000  2.540000 ;
      RECT 15.700000  2.600000 15.960000  2.860000 ;
      RECT 15.700000  2.920000 15.960000  3.180000 ;
      RECT 15.700000  3.240000 15.960000  3.500000 ;
      RECT 15.700000  3.560000 15.960000  3.820000 ;
      RECT 15.700000  3.880000 15.960000  4.140000 ;
      RECT 15.700000  4.200000 15.960000  4.460000 ;
      RECT 15.700000  4.520000 15.960000  4.780000 ;
      RECT 15.700000  4.840000 15.960000  5.100000 ;
      RECT 15.700000  5.160000 15.960000  5.420000 ;
      RECT 15.700000  6.270000 15.960000  6.530000 ;
      RECT 15.700000  6.590000 15.960000  6.850000 ;
      RECT 15.700000  6.910000 15.960000  7.170000 ;
      RECT 15.700000  7.230000 15.960000  7.490000 ;
      RECT 15.700000  7.550000 15.960000  7.810000 ;
      RECT 15.700000  7.870000 15.960000  8.130000 ;
      RECT 15.700000  8.190000 15.960000  8.450000 ;
      RECT 15.700000  8.510000 15.960000  8.770000 ;
      RECT 15.700000  8.830000 15.960000  9.090000 ;
      RECT 15.700000  9.150000 15.960000  9.410000 ;
      RECT 15.700000  9.470000 15.960000  9.730000 ;
      RECT 15.700000 13.500000 15.960000 13.760000 ;
      RECT 15.700000 13.820000 15.960000 14.080000 ;
      RECT 15.700000 14.140000 15.960000 14.400000 ;
      RECT 15.700000 14.460000 15.960000 14.720000 ;
      RECT 15.700000 14.780000 15.960000 15.040000 ;
      RECT 15.700000 15.100000 15.960000 15.360000 ;
      RECT 15.700000 15.420000 15.960000 15.680000 ;
      RECT 15.700000 15.740000 15.960000 16.000000 ;
      RECT 15.700000 16.060000 15.960000 16.320000 ;
      RECT 15.700000 16.380000 15.960000 16.640000 ;
      RECT 15.700000 16.700000 15.960000 16.960000 ;
      RECT 15.700000 17.810000 15.960000 18.070000 ;
      RECT 15.700000 18.130000 15.960000 18.390000 ;
      RECT 15.700000 18.450000 15.960000 18.710000 ;
      RECT 15.700000 18.770000 15.960000 19.030000 ;
      RECT 15.700000 19.090000 15.960000 19.350000 ;
      RECT 15.700000 19.410000 15.960000 19.670000 ;
      RECT 15.700000 19.730000 15.960000 19.990000 ;
      RECT 15.700000 20.050000 15.960000 20.310000 ;
      RECT 15.700000 20.370000 15.960000 20.630000 ;
      RECT 15.700000 20.690000 15.960000 20.950000 ;
      RECT 15.700000 21.010000 15.960000 21.270000 ;
      RECT 15.955000  0.355000 16.215000  0.615000 ;
      RECT 15.955000 11.205000 16.215000 11.465000 ;
      RECT 15.955000 11.895000 16.215000 12.155000 ;
      RECT 15.955000 22.745000 16.215000 23.005000 ;
      RECT 16.200000  1.960000 16.460000  2.220000 ;
      RECT 16.200000  2.280000 16.460000  2.540000 ;
      RECT 16.200000  2.600000 16.460000  2.860000 ;
      RECT 16.200000  2.920000 16.460000  3.180000 ;
      RECT 16.200000  3.240000 16.460000  3.500000 ;
      RECT 16.200000  3.560000 16.460000  3.820000 ;
      RECT 16.200000  3.880000 16.460000  4.140000 ;
      RECT 16.200000  4.200000 16.460000  4.460000 ;
      RECT 16.200000  4.520000 16.460000  4.780000 ;
      RECT 16.200000  4.840000 16.460000  5.100000 ;
      RECT 16.200000  5.160000 16.460000  5.420000 ;
      RECT 16.200000  6.270000 16.460000  6.530000 ;
      RECT 16.200000  6.590000 16.460000  6.850000 ;
      RECT 16.200000  6.910000 16.460000  7.170000 ;
      RECT 16.200000  7.230000 16.460000  7.490000 ;
      RECT 16.200000  7.550000 16.460000  7.810000 ;
      RECT 16.200000  7.870000 16.460000  8.130000 ;
      RECT 16.200000  8.190000 16.460000  8.450000 ;
      RECT 16.200000  8.510000 16.460000  8.770000 ;
      RECT 16.200000  8.830000 16.460000  9.090000 ;
      RECT 16.200000  9.150000 16.460000  9.410000 ;
      RECT 16.200000  9.470000 16.460000  9.730000 ;
      RECT 16.200000 13.500000 16.460000 13.760000 ;
      RECT 16.200000 13.820000 16.460000 14.080000 ;
      RECT 16.200000 14.140000 16.460000 14.400000 ;
      RECT 16.200000 14.460000 16.460000 14.720000 ;
      RECT 16.200000 14.780000 16.460000 15.040000 ;
      RECT 16.200000 15.100000 16.460000 15.360000 ;
      RECT 16.200000 15.420000 16.460000 15.680000 ;
      RECT 16.200000 15.740000 16.460000 16.000000 ;
      RECT 16.200000 16.060000 16.460000 16.320000 ;
      RECT 16.200000 16.380000 16.460000 16.640000 ;
      RECT 16.200000 16.700000 16.460000 16.960000 ;
      RECT 16.200000 17.810000 16.460000 18.070000 ;
      RECT 16.200000 18.130000 16.460000 18.390000 ;
      RECT 16.200000 18.450000 16.460000 18.710000 ;
      RECT 16.200000 18.770000 16.460000 19.030000 ;
      RECT 16.200000 19.090000 16.460000 19.350000 ;
      RECT 16.200000 19.410000 16.460000 19.670000 ;
      RECT 16.200000 19.730000 16.460000 19.990000 ;
      RECT 16.200000 20.050000 16.460000 20.310000 ;
      RECT 16.200000 20.370000 16.460000 20.630000 ;
      RECT 16.200000 20.690000 16.460000 20.950000 ;
      RECT 16.200000 21.010000 16.460000 21.270000 ;
      RECT 16.275000  0.355000 16.535000  0.615000 ;
      RECT 16.275000 11.205000 16.535000 11.465000 ;
      RECT 16.275000 11.895000 16.535000 12.155000 ;
      RECT 16.275000 22.745000 16.535000 23.005000 ;
      RECT 16.435000  5.535000 16.695000  5.795000 ;
      RECT 16.435000  5.895000 16.695000  6.155000 ;
      RECT 16.435000 17.075000 16.695000 17.335000 ;
      RECT 16.435000 17.435000 16.695000 17.695000 ;
      RECT 16.595000  0.355000 16.855000  0.615000 ;
      RECT 16.595000 11.205000 16.855000 11.465000 ;
      RECT 16.595000 11.895000 16.855000 12.155000 ;
      RECT 16.595000 22.745000 16.855000 23.005000 ;
      RECT 16.660000  1.425000 16.920000  1.685000 ;
      RECT 16.660000 10.005000 16.920000 10.265000 ;
      RECT 16.660000 12.965000 16.920000 13.225000 ;
      RECT 16.660000 21.545000 16.920000 21.805000 ;
      RECT 16.755000  5.535000 17.015000  5.795000 ;
      RECT 16.755000  5.895000 17.015000  6.155000 ;
      RECT 16.755000 17.075000 17.015000 17.335000 ;
      RECT 16.755000 17.435000 17.015000 17.695000 ;
      RECT 16.915000  0.355000 17.175000  0.615000 ;
      RECT 16.915000 11.205000 17.175000 11.465000 ;
      RECT 16.915000 11.895000 17.175000 12.155000 ;
      RECT 16.915000 22.745000 17.175000 23.005000 ;
      RECT 16.980000  1.425000 17.240000  1.685000 ;
      RECT 16.980000 10.005000 17.240000 10.265000 ;
      RECT 16.980000 12.965000 17.240000 13.225000 ;
      RECT 16.980000 21.545000 17.240000 21.805000 ;
      RECT 17.075000  5.535000 17.335000  5.795000 ;
      RECT 17.075000  5.895000 17.335000  6.155000 ;
      RECT 17.075000 17.075000 17.335000 17.335000 ;
      RECT 17.075000 17.435000 17.335000 17.695000 ;
      RECT 17.235000  0.355000 17.495000  0.615000 ;
      RECT 17.235000 11.205000 17.495000 11.465000 ;
      RECT 17.235000 11.895000 17.495000 12.155000 ;
      RECT 17.235000 22.745000 17.495000 23.005000 ;
      RECT 17.300000  1.425000 17.560000  1.685000 ;
      RECT 17.300000 10.005000 17.560000 10.265000 ;
      RECT 17.300000 12.965000 17.560000 13.225000 ;
      RECT 17.300000 21.545000 17.560000 21.805000 ;
      RECT 17.395000  5.535000 17.655000  5.795000 ;
      RECT 17.395000  5.895000 17.655000  6.155000 ;
      RECT 17.395000 17.075000 17.655000 17.335000 ;
      RECT 17.395000 17.435000 17.655000 17.695000 ;
      RECT 17.555000  0.355000 17.815000  0.615000 ;
      RECT 17.555000 11.205000 17.815000 11.465000 ;
      RECT 17.555000 11.895000 17.815000 12.155000 ;
      RECT 17.555000 22.745000 17.815000 23.005000 ;
      RECT 17.620000  1.425000 17.880000  1.685000 ;
      RECT 17.620000 10.005000 17.880000 10.265000 ;
      RECT 17.620000 12.965000 17.880000 13.225000 ;
      RECT 17.620000 21.545000 17.880000 21.805000 ;
      RECT 17.715000  5.535000 17.975000  5.795000 ;
      RECT 17.715000  5.895000 17.975000  6.155000 ;
      RECT 17.715000 17.075000 17.975000 17.335000 ;
      RECT 17.715000 17.435000 17.975000 17.695000 ;
      RECT 17.875000  0.355000 18.135000  0.615000 ;
      RECT 17.875000 11.205000 18.135000 11.465000 ;
      RECT 17.875000 11.895000 18.135000 12.155000 ;
      RECT 17.875000 22.745000 18.135000 23.005000 ;
      RECT 17.940000  1.425000 18.200000  1.685000 ;
      RECT 17.940000 10.005000 18.200000 10.265000 ;
      RECT 17.940000 12.965000 18.200000 13.225000 ;
      RECT 17.940000 21.545000 18.200000 21.805000 ;
      RECT 18.035000  5.535000 18.295000  5.795000 ;
      RECT 18.035000  5.895000 18.295000  6.155000 ;
      RECT 18.035000 17.075000 18.295000 17.335000 ;
      RECT 18.035000 17.435000 18.295000 17.695000 ;
      RECT 18.195000  0.355000 18.455000  0.615000 ;
      RECT 18.195000 11.205000 18.455000 11.465000 ;
      RECT 18.195000 11.895000 18.455000 12.155000 ;
      RECT 18.195000 22.745000 18.455000 23.005000 ;
      RECT 18.260000  1.425000 18.520000  1.685000 ;
      RECT 18.260000 10.005000 18.520000 10.265000 ;
      RECT 18.260000 12.965000 18.520000 13.225000 ;
      RECT 18.260000 21.545000 18.520000 21.805000 ;
      RECT 18.355000  5.535000 18.615000  5.795000 ;
      RECT 18.355000  5.895000 18.615000  6.155000 ;
      RECT 18.355000 17.075000 18.615000 17.335000 ;
      RECT 18.355000 17.435000 18.615000 17.695000 ;
      RECT 18.515000  0.355000 18.775000  0.615000 ;
      RECT 18.515000 11.205000 18.775000 11.465000 ;
      RECT 18.515000 11.895000 18.775000 12.155000 ;
      RECT 18.515000 22.745000 18.775000 23.005000 ;
      RECT 18.580000  1.425000 18.840000  1.685000 ;
      RECT 18.580000 10.005000 18.840000 10.265000 ;
      RECT 18.580000 12.965000 18.840000 13.225000 ;
      RECT 18.580000 21.545000 18.840000 21.805000 ;
      RECT 18.675000  5.535000 18.935000  5.795000 ;
      RECT 18.675000  5.895000 18.935000  6.155000 ;
      RECT 18.675000 17.075000 18.935000 17.335000 ;
      RECT 18.675000 17.435000 18.935000 17.695000 ;
      RECT 18.835000  0.355000 19.095000  0.615000 ;
      RECT 18.835000 11.205000 19.095000 11.465000 ;
      RECT 18.835000 11.895000 19.095000 12.155000 ;
      RECT 18.835000 22.745000 19.095000 23.005000 ;
      RECT 18.900000  1.425000 19.160000  1.685000 ;
      RECT 18.900000 10.005000 19.160000 10.265000 ;
      RECT 18.900000 12.965000 19.160000 13.225000 ;
      RECT 18.900000 21.545000 19.160000 21.805000 ;
      RECT 18.995000  5.535000 19.255000  5.795000 ;
      RECT 18.995000  5.895000 19.255000  6.155000 ;
      RECT 18.995000 17.075000 19.255000 17.335000 ;
      RECT 18.995000 17.435000 19.255000 17.695000 ;
      RECT 19.155000  0.355000 19.415000  0.615000 ;
      RECT 19.155000 11.205000 19.415000 11.465000 ;
      RECT 19.155000 11.895000 19.415000 12.155000 ;
      RECT 19.155000 22.745000 19.415000 23.005000 ;
      RECT 19.220000  1.425000 19.480000  1.685000 ;
      RECT 19.220000 10.005000 19.480000 10.265000 ;
      RECT 19.220000 12.965000 19.480000 13.225000 ;
      RECT 19.220000 21.545000 19.480000 21.805000 ;
      RECT 19.315000  5.535000 19.575000  5.795000 ;
      RECT 19.315000  5.895000 19.575000  6.155000 ;
      RECT 19.315000 17.075000 19.575000 17.335000 ;
      RECT 19.315000 17.435000 19.575000 17.695000 ;
      RECT 19.475000  0.355000 19.735000  0.615000 ;
      RECT 19.475000 11.205000 19.735000 11.465000 ;
      RECT 19.475000 11.895000 19.735000 12.155000 ;
      RECT 19.475000 22.745000 19.735000 23.005000 ;
      RECT 19.540000  1.425000 19.800000  1.685000 ;
      RECT 19.540000 10.005000 19.800000 10.265000 ;
      RECT 19.540000 12.965000 19.800000 13.225000 ;
      RECT 19.540000 21.545000 19.800000 21.805000 ;
      RECT 19.635000  5.535000 19.895000  5.795000 ;
      RECT 19.635000  5.895000 19.895000  6.155000 ;
      RECT 19.635000 17.075000 19.895000 17.335000 ;
      RECT 19.635000 17.435000 19.895000 17.695000 ;
      RECT 19.795000  0.355000 20.055000  0.615000 ;
      RECT 19.795000 11.205000 20.055000 11.465000 ;
      RECT 19.795000 11.895000 20.055000 12.155000 ;
      RECT 19.795000 22.745000 20.055000 23.005000 ;
      RECT 19.860000  1.425000 20.120000  1.685000 ;
      RECT 19.860000 10.005000 20.120000 10.265000 ;
      RECT 19.860000 12.965000 20.120000 13.225000 ;
      RECT 19.860000 21.545000 20.120000 21.805000 ;
      RECT 19.955000  5.535000 20.215000  5.795000 ;
      RECT 19.955000  5.895000 20.215000  6.155000 ;
      RECT 19.955000 17.075000 20.215000 17.335000 ;
      RECT 19.955000 17.435000 20.215000 17.695000 ;
      RECT 20.470000  1.960000 20.730000  2.220000 ;
      RECT 20.470000  2.280000 20.730000  2.540000 ;
      RECT 20.470000  2.600000 20.730000  2.860000 ;
      RECT 20.470000  2.920000 20.730000  3.180000 ;
      RECT 20.470000  3.240000 20.730000  3.500000 ;
      RECT 20.470000  3.560000 20.730000  3.820000 ;
      RECT 20.470000  3.880000 20.730000  4.140000 ;
      RECT 20.470000  4.200000 20.730000  4.460000 ;
      RECT 20.470000  4.520000 20.730000  4.780000 ;
      RECT 20.470000  4.840000 20.730000  5.100000 ;
      RECT 20.470000  5.160000 20.730000  5.420000 ;
      RECT 20.470000  6.270000 20.730000  6.530000 ;
      RECT 20.470000  6.590000 20.730000  6.850000 ;
      RECT 20.470000  6.910000 20.730000  7.170000 ;
      RECT 20.470000  7.230000 20.730000  7.490000 ;
      RECT 20.470000  7.550000 20.730000  7.810000 ;
      RECT 20.470000  7.870000 20.730000  8.130000 ;
      RECT 20.470000  8.190000 20.730000  8.450000 ;
      RECT 20.470000  8.510000 20.730000  8.770000 ;
      RECT 20.470000  8.830000 20.730000  9.090000 ;
      RECT 20.470000  9.150000 20.730000  9.410000 ;
      RECT 20.470000  9.470000 20.730000  9.730000 ;
      RECT 20.470000 13.500000 20.730000 13.760000 ;
      RECT 20.470000 13.820000 20.730000 14.080000 ;
      RECT 20.470000 14.140000 20.730000 14.400000 ;
      RECT 20.470000 14.460000 20.730000 14.720000 ;
      RECT 20.470000 14.780000 20.730000 15.040000 ;
      RECT 20.470000 15.100000 20.730000 15.360000 ;
      RECT 20.470000 15.420000 20.730000 15.680000 ;
      RECT 20.470000 15.740000 20.730000 16.000000 ;
      RECT 20.470000 16.060000 20.730000 16.320000 ;
      RECT 20.470000 16.380000 20.730000 16.640000 ;
      RECT 20.470000 16.700000 20.730000 16.960000 ;
      RECT 20.470000 17.810000 20.730000 18.070000 ;
      RECT 20.470000 18.130000 20.730000 18.390000 ;
      RECT 20.470000 18.450000 20.730000 18.710000 ;
      RECT 20.470000 18.770000 20.730000 19.030000 ;
      RECT 20.470000 19.090000 20.730000 19.350000 ;
      RECT 20.470000 19.410000 20.730000 19.670000 ;
      RECT 20.470000 19.730000 20.730000 19.990000 ;
      RECT 20.470000 20.050000 20.730000 20.310000 ;
      RECT 20.470000 20.370000 20.730000 20.630000 ;
      RECT 20.470000 20.690000 20.730000 20.950000 ;
      RECT 20.470000 21.010000 20.730000 21.270000 ;
    LAYER via2 ;
      RECT  0.325000  0.485000  0.605000  0.765000 ;
      RECT  0.325000  0.885000  0.605000  1.165000 ;
      RECT  0.325000  1.285000  0.605000  1.565000 ;
      RECT  0.325000  1.685000  0.605000  1.965000 ;
      RECT  0.325000  2.085000  0.605000  2.365000 ;
      RECT  0.325000  2.485000  0.605000  2.765000 ;
      RECT  0.325000  2.885000  0.605000  3.165000 ;
      RECT  0.325000  3.285000  0.605000  3.565000 ;
      RECT  0.325000  3.685000  0.605000  3.965000 ;
      RECT  0.325000  4.085000  0.605000  4.365000 ;
      RECT  0.325000  4.485000  0.605000  4.765000 ;
      RECT  0.325000  4.885000  0.605000  5.165000 ;
      RECT  0.325000  5.285000  0.605000  5.565000 ;
      RECT  0.325000  5.685000  0.605000  5.965000 ;
      RECT  0.325000  6.085000  0.605000  6.365000 ;
      RECT  0.325000  6.485000  0.605000  6.765000 ;
      RECT  0.325000  6.885000  0.605000  7.165000 ;
      RECT  0.325000  7.285000  0.605000  7.565000 ;
      RECT  0.325000  7.685000  0.605000  7.965000 ;
      RECT  0.325000  8.085000  0.605000  8.365000 ;
      RECT  0.325000  8.485000  0.605000  8.765000 ;
      RECT  0.325000  8.885000  0.605000  9.165000 ;
      RECT  0.325000  9.285000  0.605000  9.565000 ;
      RECT  0.325000  9.685000  0.605000  9.965000 ;
      RECT  0.325000 10.085000  0.605000 10.365000 ;
      RECT  0.325000 10.485000  0.605000 10.765000 ;
      RECT  0.325000 10.885000  0.605000 11.165000 ;
      RECT  0.325000 11.285000  0.605000 11.565000 ;
      RECT  0.325000 12.025000  0.605000 12.305000 ;
      RECT  0.325000 12.425000  0.605000 12.705000 ;
      RECT  0.325000 12.825000  0.605000 13.105000 ;
      RECT  0.325000 13.225000  0.605000 13.505000 ;
      RECT  0.325000 13.625000  0.605000 13.905000 ;
      RECT  0.325000 14.025000  0.605000 14.305000 ;
      RECT  0.325000 14.425000  0.605000 14.705000 ;
      RECT  0.325000 14.825000  0.605000 15.105000 ;
      RECT  0.325000 15.225000  0.605000 15.505000 ;
      RECT  0.325000 15.625000  0.605000 15.905000 ;
      RECT  0.325000 16.025000  0.605000 16.305000 ;
      RECT  0.325000 16.425000  0.605000 16.705000 ;
      RECT  0.325000 16.825000  0.605000 17.105000 ;
      RECT  0.325000 17.225000  0.605000 17.505000 ;
      RECT  0.325000 17.625000  0.605000 17.905000 ;
      RECT  0.325000 18.025000  0.605000 18.305000 ;
      RECT  0.325000 18.425000  0.605000 18.705000 ;
      RECT  0.325000 18.825000  0.605000 19.105000 ;
      RECT  0.325000 19.225000  0.605000 19.505000 ;
      RECT  0.325000 19.625000  0.605000 19.905000 ;
      RECT  0.325000 20.025000  0.605000 20.305000 ;
      RECT  0.325000 20.425000  0.605000 20.705000 ;
      RECT  0.325000 20.825000  0.605000 21.105000 ;
      RECT  0.325000 21.225000  0.605000 21.505000 ;
      RECT  0.325000 21.625000  0.605000 21.905000 ;
      RECT  0.325000 22.025000  0.605000 22.305000 ;
      RECT  0.325000 22.425000  0.605000 22.705000 ;
      RECT  0.325000 22.825000  0.605000 23.105000 ;
      RECT  0.990000  1.490000  1.270000  1.770000 ;
      RECT  0.990000  1.890000  1.270000  2.170000 ;
      RECT  0.990000  2.290000  1.270000  2.570000 ;
      RECT  0.990000  2.690000  1.270000  2.970000 ;
      RECT  0.990000  3.090000  1.270000  3.370000 ;
      RECT  0.990000  3.490000  1.270000  3.770000 ;
      RECT  0.990000  3.890000  1.270000  4.170000 ;
      RECT  0.990000  4.290000  1.270000  4.570000 ;
      RECT  0.990000  4.690000  1.270000  4.970000 ;
      RECT  0.990000  5.090000  1.270000  5.370000 ;
      RECT  0.990000  5.490000  1.270000  5.770000 ;
      RECT  0.990000  5.890000  1.270000  6.170000 ;
      RECT  0.990000  6.290000  1.270000  6.570000 ;
      RECT  0.990000  6.690000  1.270000  6.970000 ;
      RECT  0.990000  7.090000  1.270000  7.370000 ;
      RECT  0.990000  7.490000  1.270000  7.770000 ;
      RECT  0.990000  7.890000  1.270000  8.170000 ;
      RECT  0.990000  8.290000  1.270000  8.570000 ;
      RECT  0.990000  8.690000  1.270000  8.970000 ;
      RECT  0.990000  9.090000  1.270000  9.370000 ;
      RECT  0.990000  9.490000  1.270000  9.770000 ;
      RECT  0.990000  9.890000  1.270000 10.170000 ;
      RECT  0.990000 13.030000  1.270000 13.310000 ;
      RECT  0.990000 13.430000  1.270000 13.710000 ;
      RECT  0.990000 13.830000  1.270000 14.110000 ;
      RECT  0.990000 14.230000  1.270000 14.510000 ;
      RECT  0.990000 14.630000  1.270000 14.910000 ;
      RECT  0.990000 15.030000  1.270000 15.310000 ;
      RECT  0.990000 15.430000  1.270000 15.710000 ;
      RECT  0.990000 15.830000  1.270000 16.110000 ;
      RECT  0.990000 16.230000  1.270000 16.510000 ;
      RECT  0.990000 16.630000  1.270000 16.910000 ;
      RECT  0.990000 17.030000  1.270000 17.310000 ;
      RECT  0.990000 17.430000  1.270000 17.710000 ;
      RECT  0.990000 17.830000  1.270000 18.110000 ;
      RECT  0.990000 18.230000  1.270000 18.510000 ;
      RECT  0.990000 18.630000  1.270000 18.910000 ;
      RECT  0.990000 19.030000  1.270000 19.310000 ;
      RECT  0.990000 19.430000  1.270000 19.710000 ;
      RECT  0.990000 19.830000  1.270000 20.110000 ;
      RECT  0.990000 20.230000  1.270000 20.510000 ;
      RECT  0.990000 20.630000  1.270000 20.910000 ;
      RECT  0.990000 21.030000  1.270000 21.310000 ;
      RECT  0.990000 21.430000  1.270000 21.710000 ;
      RECT  1.620000  5.690000  1.900000  5.970000 ;
      RECT  1.620000 17.230000  1.900000 17.510000 ;
      RECT  2.020000  5.690000  2.300000  5.970000 ;
      RECT  2.020000 17.230000  2.300000 17.510000 ;
      RECT  2.420000  5.690000  2.700000  5.970000 ;
      RECT  2.420000 17.230000  2.700000 17.510000 ;
      RECT  2.820000  5.690000  3.100000  5.970000 ;
      RECT  2.820000 17.230000  3.100000 17.510000 ;
      RECT  3.220000  5.690000  3.500000  5.970000 ;
      RECT  3.220000 17.230000  3.500000 17.510000 ;
      RECT  3.620000  5.690000  3.900000  5.970000 ;
      RECT  3.620000 17.230000  3.900000 17.510000 ;
      RECT  4.020000  5.690000  4.300000  5.970000 ;
      RECT  4.020000 17.230000  4.300000 17.510000 ;
      RECT  4.420000  5.690000  4.700000  5.970000 ;
      RECT  4.420000 17.230000  4.700000 17.510000 ;
      RECT  4.820000  5.690000  5.100000  5.970000 ;
      RECT  4.820000 17.230000  5.100000 17.510000 ;
      RECT  5.530000  0.890000  5.810000  1.170000 ;
      RECT  5.530000  1.290000  5.810000  1.570000 ;
      RECT  5.530000  1.690000  5.810000  1.970000 ;
      RECT  5.530000  2.090000  5.810000  2.370000 ;
      RECT  5.530000  2.490000  5.810000  2.770000 ;
      RECT  5.530000  2.890000  5.810000  3.170000 ;
      RECT  5.530000  3.290000  5.810000  3.570000 ;
      RECT  5.530000  3.690000  5.810000  3.970000 ;
      RECT  5.530000  4.090000  5.810000  4.370000 ;
      RECT  5.530000  4.490000  5.810000  4.770000 ;
      RECT  5.530000  4.890000  5.810000  5.170000 ;
      RECT  5.530000  5.290000  5.810000  5.570000 ;
      RECT  5.530000  5.690000  5.810000  5.970000 ;
      RECT  5.530000  6.090000  5.810000  6.370000 ;
      RECT  5.530000  6.490000  5.810000  6.770000 ;
      RECT  5.530000  6.890000  5.810000  7.170000 ;
      RECT  5.530000  7.290000  5.810000  7.570000 ;
      RECT  5.530000  7.690000  5.810000  7.970000 ;
      RECT  5.530000  8.090000  5.810000  8.370000 ;
      RECT  5.530000  8.490000  5.810000  8.770000 ;
      RECT  5.530000  8.890000  5.810000  9.170000 ;
      RECT  5.530000  9.290000  5.810000  9.570000 ;
      RECT  5.530000  9.690000  5.810000  9.970000 ;
      RECT  5.530000 10.090000  5.810000 10.370000 ;
      RECT  5.530000 10.490000  5.810000 10.770000 ;
      RECT  5.530000 12.430000  5.810000 12.710000 ;
      RECT  5.530000 12.830000  5.810000 13.110000 ;
      RECT  5.530000 13.230000  5.810000 13.510000 ;
      RECT  5.530000 13.630000  5.810000 13.910000 ;
      RECT  5.530000 14.030000  5.810000 14.310000 ;
      RECT  5.530000 14.430000  5.810000 14.710000 ;
      RECT  5.530000 14.830000  5.810000 15.110000 ;
      RECT  5.530000 15.230000  5.810000 15.510000 ;
      RECT  5.530000 15.630000  5.810000 15.910000 ;
      RECT  5.530000 16.030000  5.810000 16.310000 ;
      RECT  5.530000 16.430000  5.810000 16.710000 ;
      RECT  5.530000 16.830000  5.810000 17.110000 ;
      RECT  5.530000 17.230000  5.810000 17.510000 ;
      RECT  5.530000 17.630000  5.810000 17.910000 ;
      RECT  5.530000 18.030000  5.810000 18.310000 ;
      RECT  5.530000 18.430000  5.810000 18.710000 ;
      RECT  5.530000 18.830000  5.810000 19.110000 ;
      RECT  5.530000 19.230000  5.810000 19.510000 ;
      RECT  5.530000 19.630000  5.810000 19.910000 ;
      RECT  5.530000 20.030000  5.810000 20.310000 ;
      RECT  5.530000 20.430000  5.810000 20.710000 ;
      RECT  5.530000 20.830000  5.810000 21.110000 ;
      RECT  5.530000 21.230000  5.810000 21.510000 ;
      RECT  5.530000 21.630000  5.810000 21.910000 ;
      RECT  5.530000 22.030000  5.810000 22.310000 ;
      RECT  6.240000  5.690000  6.520000  5.970000 ;
      RECT  6.240000 17.230000  6.520000 17.510000 ;
      RECT  6.640000  5.690000  6.920000  5.970000 ;
      RECT  6.640000 17.230000  6.920000 17.510000 ;
      RECT  7.040000  5.690000  7.320000  5.970000 ;
      RECT  7.040000 17.230000  7.320000 17.510000 ;
      RECT  7.440000  5.690000  7.720000  5.970000 ;
      RECT  7.440000 17.230000  7.720000 17.510000 ;
      RECT  7.840000  5.690000  8.120000  5.970000 ;
      RECT  7.840000 17.230000  8.120000 17.510000 ;
      RECT  8.240000  5.690000  8.520000  5.970000 ;
      RECT  8.240000 17.230000  8.520000 17.510000 ;
      RECT  8.640000  5.690000  8.920000  5.970000 ;
      RECT  8.640000 17.230000  8.920000 17.510000 ;
      RECT  9.040000  5.690000  9.320000  5.970000 ;
      RECT  9.040000 17.230000  9.320000 17.510000 ;
      RECT  9.440000  5.690000  9.720000  5.970000 ;
      RECT  9.440000 17.230000  9.720000 17.510000 ;
      RECT 10.070000  1.490000 10.350000  1.770000 ;
      RECT 10.070000  1.890000 10.350000  2.170000 ;
      RECT 10.070000  2.290000 10.350000  2.570000 ;
      RECT 10.070000  2.690000 10.350000  2.970000 ;
      RECT 10.070000  3.090000 10.350000  3.370000 ;
      RECT 10.070000  3.490000 10.350000  3.770000 ;
      RECT 10.070000  3.890000 10.350000  4.170000 ;
      RECT 10.070000  4.290000 10.350000  4.570000 ;
      RECT 10.070000  4.690000 10.350000  4.970000 ;
      RECT 10.070000  5.090000 10.350000  5.370000 ;
      RECT 10.070000  5.490000 10.350000  5.770000 ;
      RECT 10.070000  5.890000 10.350000  6.170000 ;
      RECT 10.070000  6.290000 10.350000  6.570000 ;
      RECT 10.070000  6.690000 10.350000  6.970000 ;
      RECT 10.070000  7.090000 10.350000  7.370000 ;
      RECT 10.070000  7.490000 10.350000  7.770000 ;
      RECT 10.070000  7.890000 10.350000  8.170000 ;
      RECT 10.070000  8.290000 10.350000  8.570000 ;
      RECT 10.070000  8.690000 10.350000  8.970000 ;
      RECT 10.070000  9.090000 10.350000  9.370000 ;
      RECT 10.070000  9.490000 10.350000  9.770000 ;
      RECT 10.070000  9.890000 10.350000 10.170000 ;
      RECT 10.070000 13.030000 10.350000 13.310000 ;
      RECT 10.070000 13.430000 10.350000 13.710000 ;
      RECT 10.070000 13.830000 10.350000 14.110000 ;
      RECT 10.070000 14.230000 10.350000 14.510000 ;
      RECT 10.070000 14.630000 10.350000 14.910000 ;
      RECT 10.070000 15.030000 10.350000 15.310000 ;
      RECT 10.070000 15.430000 10.350000 15.710000 ;
      RECT 10.070000 15.830000 10.350000 16.110000 ;
      RECT 10.070000 16.230000 10.350000 16.510000 ;
      RECT 10.070000 16.630000 10.350000 16.910000 ;
      RECT 10.070000 17.030000 10.350000 17.310000 ;
      RECT 10.070000 17.430000 10.350000 17.710000 ;
      RECT 10.070000 17.830000 10.350000 18.110000 ;
      RECT 10.070000 18.230000 10.350000 18.510000 ;
      RECT 10.070000 18.630000 10.350000 18.910000 ;
      RECT 10.070000 19.030000 10.350000 19.310000 ;
      RECT 10.070000 19.430000 10.350000 19.710000 ;
      RECT 10.070000 19.830000 10.350000 20.110000 ;
      RECT 10.070000 20.230000 10.350000 20.510000 ;
      RECT 10.070000 20.630000 10.350000 20.910000 ;
      RECT 10.070000 21.030000 10.350000 21.310000 ;
      RECT 10.070000 21.430000 10.350000 21.710000 ;
      RECT 10.735000  0.485000 11.015000  0.765000 ;
      RECT 10.735000  0.885000 11.015000  1.165000 ;
      RECT 10.735000  1.285000 11.015000  1.565000 ;
      RECT 10.735000  1.685000 11.015000  1.965000 ;
      RECT 10.735000  2.085000 11.015000  2.365000 ;
      RECT 10.735000  2.485000 11.015000  2.765000 ;
      RECT 10.735000  2.885000 11.015000  3.165000 ;
      RECT 10.735000  3.285000 11.015000  3.565000 ;
      RECT 10.735000  3.685000 11.015000  3.965000 ;
      RECT 10.735000  4.085000 11.015000  4.365000 ;
      RECT 10.735000  4.485000 11.015000  4.765000 ;
      RECT 10.735000  4.885000 11.015000  5.165000 ;
      RECT 10.735000  5.285000 11.015000  5.565000 ;
      RECT 10.735000  5.685000 11.015000  5.965000 ;
      RECT 10.735000  6.085000 11.015000  6.365000 ;
      RECT 10.735000  6.485000 11.015000  6.765000 ;
      RECT 10.735000  6.885000 11.015000  7.165000 ;
      RECT 10.735000  7.285000 11.015000  7.565000 ;
      RECT 10.735000  7.685000 11.015000  7.965000 ;
      RECT 10.735000  8.085000 11.015000  8.365000 ;
      RECT 10.735000  8.485000 11.015000  8.765000 ;
      RECT 10.735000  8.885000 11.015000  9.165000 ;
      RECT 10.735000  9.285000 11.015000  9.565000 ;
      RECT 10.735000  9.685000 11.015000  9.965000 ;
      RECT 10.735000 10.085000 11.015000 10.365000 ;
      RECT 10.735000 10.485000 11.015000 10.765000 ;
      RECT 10.735000 10.885000 11.015000 11.165000 ;
      RECT 10.735000 11.285000 11.015000 11.565000 ;
      RECT 10.735000 12.025000 11.015000 12.305000 ;
      RECT 10.735000 12.425000 11.015000 12.705000 ;
      RECT 10.735000 12.825000 11.015000 13.105000 ;
      RECT 10.735000 13.225000 11.015000 13.505000 ;
      RECT 10.735000 13.625000 11.015000 13.905000 ;
      RECT 10.735000 14.025000 11.015000 14.305000 ;
      RECT 10.735000 14.425000 11.015000 14.705000 ;
      RECT 10.735000 14.825000 11.015000 15.105000 ;
      RECT 10.735000 15.225000 11.015000 15.505000 ;
      RECT 10.735000 15.625000 11.015000 15.905000 ;
      RECT 10.735000 16.025000 11.015000 16.305000 ;
      RECT 10.735000 16.425000 11.015000 16.705000 ;
      RECT 10.735000 16.825000 11.015000 17.105000 ;
      RECT 10.735000 17.225000 11.015000 17.505000 ;
      RECT 10.735000 17.625000 11.015000 17.905000 ;
      RECT 10.735000 18.025000 11.015000 18.305000 ;
      RECT 10.735000 18.425000 11.015000 18.705000 ;
      RECT 10.735000 18.825000 11.015000 19.105000 ;
      RECT 10.735000 19.225000 11.015000 19.505000 ;
      RECT 10.735000 19.625000 11.015000 19.905000 ;
      RECT 10.735000 20.025000 11.015000 20.305000 ;
      RECT 10.735000 20.425000 11.015000 20.705000 ;
      RECT 10.735000 20.825000 11.015000 21.105000 ;
      RECT 10.735000 21.225000 11.015000 21.505000 ;
      RECT 10.735000 21.625000 11.015000 21.905000 ;
      RECT 10.735000 22.025000 11.015000 22.305000 ;
      RECT 10.735000 22.425000 11.015000 22.705000 ;
      RECT 10.735000 22.825000 11.015000 23.105000 ;
      RECT 11.400000  1.490000 11.680000  1.770000 ;
      RECT 11.400000  1.890000 11.680000  2.170000 ;
      RECT 11.400000  2.290000 11.680000  2.570000 ;
      RECT 11.400000  2.690000 11.680000  2.970000 ;
      RECT 11.400000  3.090000 11.680000  3.370000 ;
      RECT 11.400000  3.490000 11.680000  3.770000 ;
      RECT 11.400000  3.890000 11.680000  4.170000 ;
      RECT 11.400000  4.290000 11.680000  4.570000 ;
      RECT 11.400000  4.690000 11.680000  4.970000 ;
      RECT 11.400000  5.090000 11.680000  5.370000 ;
      RECT 11.400000  5.490000 11.680000  5.770000 ;
      RECT 11.400000  5.890000 11.680000  6.170000 ;
      RECT 11.400000  6.290000 11.680000  6.570000 ;
      RECT 11.400000  6.690000 11.680000  6.970000 ;
      RECT 11.400000  7.090000 11.680000  7.370000 ;
      RECT 11.400000  7.490000 11.680000  7.770000 ;
      RECT 11.400000  7.890000 11.680000  8.170000 ;
      RECT 11.400000  8.290000 11.680000  8.570000 ;
      RECT 11.400000  8.690000 11.680000  8.970000 ;
      RECT 11.400000  9.090000 11.680000  9.370000 ;
      RECT 11.400000  9.490000 11.680000  9.770000 ;
      RECT 11.400000  9.890000 11.680000 10.170000 ;
      RECT 11.400000 13.030000 11.680000 13.310000 ;
      RECT 11.400000 13.430000 11.680000 13.710000 ;
      RECT 11.400000 13.830000 11.680000 14.110000 ;
      RECT 11.400000 14.230000 11.680000 14.510000 ;
      RECT 11.400000 14.630000 11.680000 14.910000 ;
      RECT 11.400000 15.030000 11.680000 15.310000 ;
      RECT 11.400000 15.430000 11.680000 15.710000 ;
      RECT 11.400000 15.830000 11.680000 16.110000 ;
      RECT 11.400000 16.230000 11.680000 16.510000 ;
      RECT 11.400000 16.630000 11.680000 16.910000 ;
      RECT 11.400000 17.030000 11.680000 17.310000 ;
      RECT 11.400000 17.430000 11.680000 17.710000 ;
      RECT 11.400000 17.830000 11.680000 18.110000 ;
      RECT 11.400000 18.230000 11.680000 18.510000 ;
      RECT 11.400000 18.630000 11.680000 18.910000 ;
      RECT 11.400000 19.030000 11.680000 19.310000 ;
      RECT 11.400000 19.430000 11.680000 19.710000 ;
      RECT 11.400000 19.830000 11.680000 20.110000 ;
      RECT 11.400000 20.230000 11.680000 20.510000 ;
      RECT 11.400000 20.630000 11.680000 20.910000 ;
      RECT 11.400000 21.030000 11.680000 21.310000 ;
      RECT 11.400000 21.430000 11.680000 21.710000 ;
      RECT 12.030000  5.690000 12.310000  5.970000 ;
      RECT 12.030000 17.230000 12.310000 17.510000 ;
      RECT 12.430000  5.690000 12.710000  5.970000 ;
      RECT 12.430000 17.230000 12.710000 17.510000 ;
      RECT 12.830000  5.690000 13.110000  5.970000 ;
      RECT 12.830000 17.230000 13.110000 17.510000 ;
      RECT 13.230000  5.690000 13.510000  5.970000 ;
      RECT 13.230000 17.230000 13.510000 17.510000 ;
      RECT 13.630000  5.690000 13.910000  5.970000 ;
      RECT 13.630000 17.230000 13.910000 17.510000 ;
      RECT 14.030000  5.690000 14.310000  5.970000 ;
      RECT 14.030000 17.230000 14.310000 17.510000 ;
      RECT 14.430000  5.690000 14.710000  5.970000 ;
      RECT 14.430000 17.230000 14.710000 17.510000 ;
      RECT 14.830000  5.690000 15.110000  5.970000 ;
      RECT 14.830000 17.230000 15.110000 17.510000 ;
      RECT 15.230000  5.690000 15.510000  5.970000 ;
      RECT 15.230000 17.230000 15.510000 17.510000 ;
      RECT 15.940000  0.890000 16.220000  1.170000 ;
      RECT 15.940000  1.290000 16.220000  1.570000 ;
      RECT 15.940000  1.690000 16.220000  1.970000 ;
      RECT 15.940000  2.090000 16.220000  2.370000 ;
      RECT 15.940000  2.490000 16.220000  2.770000 ;
      RECT 15.940000  2.890000 16.220000  3.170000 ;
      RECT 15.940000  3.290000 16.220000  3.570000 ;
      RECT 15.940000  3.690000 16.220000  3.970000 ;
      RECT 15.940000  4.090000 16.220000  4.370000 ;
      RECT 15.940000  4.490000 16.220000  4.770000 ;
      RECT 15.940000  4.890000 16.220000  5.170000 ;
      RECT 15.940000  5.290000 16.220000  5.570000 ;
      RECT 15.940000  5.690000 16.220000  5.970000 ;
      RECT 15.940000  6.090000 16.220000  6.370000 ;
      RECT 15.940000  6.490000 16.220000  6.770000 ;
      RECT 15.940000  6.890000 16.220000  7.170000 ;
      RECT 15.940000  7.290000 16.220000  7.570000 ;
      RECT 15.940000  7.690000 16.220000  7.970000 ;
      RECT 15.940000  8.090000 16.220000  8.370000 ;
      RECT 15.940000  8.490000 16.220000  8.770000 ;
      RECT 15.940000  8.890000 16.220000  9.170000 ;
      RECT 15.940000  9.290000 16.220000  9.570000 ;
      RECT 15.940000  9.690000 16.220000  9.970000 ;
      RECT 15.940000 10.090000 16.220000 10.370000 ;
      RECT 15.940000 10.490000 16.220000 10.770000 ;
      RECT 15.940000 12.430000 16.220000 12.710000 ;
      RECT 15.940000 12.830000 16.220000 13.110000 ;
      RECT 15.940000 13.230000 16.220000 13.510000 ;
      RECT 15.940000 13.630000 16.220000 13.910000 ;
      RECT 15.940000 14.030000 16.220000 14.310000 ;
      RECT 15.940000 14.430000 16.220000 14.710000 ;
      RECT 15.940000 14.830000 16.220000 15.110000 ;
      RECT 15.940000 15.230000 16.220000 15.510000 ;
      RECT 15.940000 15.630000 16.220000 15.910000 ;
      RECT 15.940000 16.030000 16.220000 16.310000 ;
      RECT 15.940000 16.430000 16.220000 16.710000 ;
      RECT 15.940000 16.830000 16.220000 17.110000 ;
      RECT 15.940000 17.230000 16.220000 17.510000 ;
      RECT 15.940000 17.630000 16.220000 17.910000 ;
      RECT 15.940000 18.030000 16.220000 18.310000 ;
      RECT 15.940000 18.430000 16.220000 18.710000 ;
      RECT 15.940000 18.830000 16.220000 19.110000 ;
      RECT 15.940000 19.230000 16.220000 19.510000 ;
      RECT 15.940000 19.630000 16.220000 19.910000 ;
      RECT 15.940000 20.030000 16.220000 20.310000 ;
      RECT 15.940000 20.430000 16.220000 20.710000 ;
      RECT 15.940000 20.830000 16.220000 21.110000 ;
      RECT 15.940000 21.230000 16.220000 21.510000 ;
      RECT 15.940000 21.630000 16.220000 21.910000 ;
      RECT 15.940000 22.030000 16.220000 22.310000 ;
      RECT 16.650000  5.690000 16.930000  5.970000 ;
      RECT 16.650000 17.230000 16.930000 17.510000 ;
      RECT 17.050000  5.690000 17.330000  5.970000 ;
      RECT 17.050000 17.230000 17.330000 17.510000 ;
      RECT 17.450000  5.690000 17.730000  5.970000 ;
      RECT 17.450000 17.230000 17.730000 17.510000 ;
      RECT 17.850000  5.690000 18.130000  5.970000 ;
      RECT 17.850000 17.230000 18.130000 17.510000 ;
      RECT 18.250000  5.690000 18.530000  5.970000 ;
      RECT 18.250000 17.230000 18.530000 17.510000 ;
      RECT 18.650000  5.690000 18.930000  5.970000 ;
      RECT 18.650000 17.230000 18.930000 17.510000 ;
      RECT 19.050000  5.690000 19.330000  5.970000 ;
      RECT 19.050000 17.230000 19.330000 17.510000 ;
      RECT 19.450000  5.690000 19.730000  5.970000 ;
      RECT 19.450000 17.230000 19.730000 17.510000 ;
      RECT 19.850000  5.690000 20.130000  5.970000 ;
      RECT 19.850000 17.230000 20.130000 17.510000 ;
      RECT 20.480000  1.490000 20.760000  1.770000 ;
      RECT 20.480000  1.890000 20.760000  2.170000 ;
      RECT 20.480000  2.290000 20.760000  2.570000 ;
      RECT 20.480000  2.690000 20.760000  2.970000 ;
      RECT 20.480000  3.090000 20.760000  3.370000 ;
      RECT 20.480000  3.490000 20.760000  3.770000 ;
      RECT 20.480000  3.890000 20.760000  4.170000 ;
      RECT 20.480000  4.290000 20.760000  4.570000 ;
      RECT 20.480000  4.690000 20.760000  4.970000 ;
      RECT 20.480000  5.090000 20.760000  5.370000 ;
      RECT 20.480000  5.490000 20.760000  5.770000 ;
      RECT 20.480000  5.890000 20.760000  6.170000 ;
      RECT 20.480000  6.290000 20.760000  6.570000 ;
      RECT 20.480000  6.690000 20.760000  6.970000 ;
      RECT 20.480000  7.090000 20.760000  7.370000 ;
      RECT 20.480000  7.490000 20.760000  7.770000 ;
      RECT 20.480000  7.890000 20.760000  8.170000 ;
      RECT 20.480000  8.290000 20.760000  8.570000 ;
      RECT 20.480000  8.690000 20.760000  8.970000 ;
      RECT 20.480000  9.090000 20.760000  9.370000 ;
      RECT 20.480000  9.490000 20.760000  9.770000 ;
      RECT 20.480000  9.890000 20.760000 10.170000 ;
      RECT 20.480000 13.030000 20.760000 13.310000 ;
      RECT 20.480000 13.430000 20.760000 13.710000 ;
      RECT 20.480000 13.830000 20.760000 14.110000 ;
      RECT 20.480000 14.230000 20.760000 14.510000 ;
      RECT 20.480000 14.630000 20.760000 14.910000 ;
      RECT 20.480000 15.030000 20.760000 15.310000 ;
      RECT 20.480000 15.430000 20.760000 15.710000 ;
      RECT 20.480000 15.830000 20.760000 16.110000 ;
      RECT 20.480000 16.230000 20.760000 16.510000 ;
      RECT 20.480000 16.630000 20.760000 16.910000 ;
      RECT 20.480000 17.030000 20.760000 17.310000 ;
      RECT 20.480000 17.430000 20.760000 17.710000 ;
      RECT 20.480000 17.830000 20.760000 18.110000 ;
      RECT 20.480000 18.230000 20.760000 18.510000 ;
      RECT 20.480000 18.630000 20.760000 18.910000 ;
      RECT 20.480000 19.030000 20.760000 19.310000 ;
      RECT 20.480000 19.430000 20.760000 19.710000 ;
      RECT 20.480000 19.830000 20.760000 20.110000 ;
      RECT 20.480000 20.230000 20.760000 20.510000 ;
      RECT 20.480000 20.630000 20.760000 20.910000 ;
      RECT 20.480000 21.030000 20.760000 21.310000 ;
      RECT 20.480000 21.430000 20.760000 21.710000 ;
      RECT 21.145000  0.485000 21.425000  0.765000 ;
      RECT 21.145000  0.885000 21.425000  1.165000 ;
      RECT 21.145000  1.285000 21.425000  1.565000 ;
      RECT 21.145000  1.685000 21.425000  1.965000 ;
      RECT 21.145000  2.085000 21.425000  2.365000 ;
      RECT 21.145000  2.485000 21.425000  2.765000 ;
      RECT 21.145000  2.885000 21.425000  3.165000 ;
      RECT 21.145000  3.285000 21.425000  3.565000 ;
      RECT 21.145000  3.685000 21.425000  3.965000 ;
      RECT 21.145000  4.085000 21.425000  4.365000 ;
      RECT 21.145000  4.485000 21.425000  4.765000 ;
      RECT 21.145000  4.885000 21.425000  5.165000 ;
      RECT 21.145000  5.285000 21.425000  5.565000 ;
      RECT 21.145000  5.685000 21.425000  5.965000 ;
      RECT 21.145000  6.085000 21.425000  6.365000 ;
      RECT 21.145000  6.485000 21.425000  6.765000 ;
      RECT 21.145000  6.885000 21.425000  7.165000 ;
      RECT 21.145000  7.285000 21.425000  7.565000 ;
      RECT 21.145000  7.685000 21.425000  7.965000 ;
      RECT 21.145000  8.085000 21.425000  8.365000 ;
      RECT 21.145000  8.485000 21.425000  8.765000 ;
      RECT 21.145000  8.885000 21.425000  9.165000 ;
      RECT 21.145000  9.285000 21.425000  9.565000 ;
      RECT 21.145000  9.685000 21.425000  9.965000 ;
      RECT 21.145000 10.085000 21.425000 10.365000 ;
      RECT 21.145000 10.485000 21.425000 10.765000 ;
      RECT 21.145000 10.885000 21.425000 11.165000 ;
      RECT 21.145000 11.285000 21.425000 11.565000 ;
      RECT 21.145000 12.025000 21.425000 12.305000 ;
      RECT 21.145000 12.425000 21.425000 12.705000 ;
      RECT 21.145000 12.825000 21.425000 13.105000 ;
      RECT 21.145000 13.225000 21.425000 13.505000 ;
      RECT 21.145000 13.625000 21.425000 13.905000 ;
      RECT 21.145000 14.025000 21.425000 14.305000 ;
      RECT 21.145000 14.425000 21.425000 14.705000 ;
      RECT 21.145000 14.825000 21.425000 15.105000 ;
      RECT 21.145000 15.225000 21.425000 15.505000 ;
      RECT 21.145000 15.625000 21.425000 15.905000 ;
      RECT 21.145000 16.025000 21.425000 16.305000 ;
      RECT 21.145000 16.425000 21.425000 16.705000 ;
      RECT 21.145000 16.825000 21.425000 17.105000 ;
      RECT 21.145000 17.225000 21.425000 17.505000 ;
      RECT 21.145000 17.625000 21.425000 17.905000 ;
      RECT 21.145000 18.025000 21.425000 18.305000 ;
      RECT 21.145000 18.425000 21.425000 18.705000 ;
      RECT 21.145000 18.825000 21.425000 19.105000 ;
      RECT 21.145000 19.225000 21.425000 19.505000 ;
      RECT 21.145000 19.625000 21.425000 19.905000 ;
      RECT 21.145000 20.025000 21.425000 20.305000 ;
      RECT 21.145000 20.425000 21.425000 20.705000 ;
      RECT 21.145000 20.825000 21.425000 21.105000 ;
      RECT 21.145000 21.225000 21.425000 21.505000 ;
      RECT 21.145000 21.625000 21.425000 21.905000 ;
      RECT 21.145000 22.025000 21.425000 22.305000 ;
      RECT 21.145000 22.425000 21.425000 22.705000 ;
      RECT 21.145000 22.825000 21.425000 23.105000 ;
    LAYER via3 ;
      RECT  0.305000  0.465000  0.625000  0.785000 ;
      RECT  0.305000  0.865000  0.625000  1.185000 ;
      RECT  0.305000  1.265000  0.625000  1.585000 ;
      RECT  0.305000  1.665000  0.625000  1.985000 ;
      RECT  0.305000  2.065000  0.625000  2.385000 ;
      RECT  0.305000  2.465000  0.625000  2.785000 ;
      RECT  0.305000  2.865000  0.625000  3.185000 ;
      RECT  0.305000  3.265000  0.625000  3.585000 ;
      RECT  0.305000  3.665000  0.625000  3.985000 ;
      RECT  0.305000  4.065000  0.625000  4.385000 ;
      RECT  0.305000  4.465000  0.625000  4.785000 ;
      RECT  0.305000  4.865000  0.625000  5.185000 ;
      RECT  0.305000  5.265000  0.625000  5.585000 ;
      RECT  0.305000  5.665000  0.625000  5.985000 ;
      RECT  0.305000  6.065000  0.625000  6.385000 ;
      RECT  0.305000  6.465000  0.625000  6.785000 ;
      RECT  0.305000  6.865000  0.625000  7.185000 ;
      RECT  0.305000  7.265000  0.625000  7.585000 ;
      RECT  0.305000  7.665000  0.625000  7.985000 ;
      RECT  0.305000  8.065000  0.625000  8.385000 ;
      RECT  0.305000  8.465000  0.625000  8.785000 ;
      RECT  0.305000  8.865000  0.625000  9.185000 ;
      RECT  0.305000  9.265000  0.625000  9.585000 ;
      RECT  0.305000  9.665000  0.625000  9.985000 ;
      RECT  0.305000 10.065000  0.625000 10.385000 ;
      RECT  0.305000 10.465000  0.625000 10.785000 ;
      RECT  0.305000 10.865000  0.625000 11.185000 ;
      RECT  0.305000 11.265000  0.625000 11.585000 ;
      RECT  0.305000 12.005000  0.625000 12.325000 ;
      RECT  0.305000 12.405000  0.625000 12.725000 ;
      RECT  0.305000 12.805000  0.625000 13.125000 ;
      RECT  0.305000 13.205000  0.625000 13.525000 ;
      RECT  0.305000 13.605000  0.625000 13.925000 ;
      RECT  0.305000 14.005000  0.625000 14.325000 ;
      RECT  0.305000 14.405000  0.625000 14.725000 ;
      RECT  0.305000 14.805000  0.625000 15.125000 ;
      RECT  0.305000 15.205000  0.625000 15.525000 ;
      RECT  0.305000 15.605000  0.625000 15.925000 ;
      RECT  0.305000 16.005000  0.625000 16.325000 ;
      RECT  0.305000 16.405000  0.625000 16.725000 ;
      RECT  0.305000 16.805000  0.625000 17.125000 ;
      RECT  0.305000 17.205000  0.625000 17.525000 ;
      RECT  0.305000 17.605000  0.625000 17.925000 ;
      RECT  0.305000 18.005000  0.625000 18.325000 ;
      RECT  0.305000 18.405000  0.625000 18.725000 ;
      RECT  0.305000 18.805000  0.625000 19.125000 ;
      RECT  0.305000 19.205000  0.625000 19.525000 ;
      RECT  0.305000 19.605000  0.625000 19.925000 ;
      RECT  0.305000 20.005000  0.625000 20.325000 ;
      RECT  0.305000 20.405000  0.625000 20.725000 ;
      RECT  0.305000 20.805000  0.625000 21.125000 ;
      RECT  0.305000 21.205000  0.625000 21.525000 ;
      RECT  0.305000 21.605000  0.625000 21.925000 ;
      RECT  0.305000 22.005000  0.625000 22.325000 ;
      RECT  0.305000 22.405000  0.625000 22.725000 ;
      RECT  0.305000 22.805000  0.625000 23.125000 ;
      RECT  0.970000  0.670000  1.290000  0.990000 ;
      RECT  0.970000  1.070000  1.290000  1.390000 ;
      RECT  0.970000  1.470000  1.290000  1.790000 ;
      RECT  0.970000  1.870000  1.290000  2.190000 ;
      RECT  0.970000  2.270000  1.290000  2.590000 ;
      RECT  0.970000  2.670000  1.290000  2.990000 ;
      RECT  0.970000  3.070000  1.290000  3.390000 ;
      RECT  0.970000  3.470000  1.290000  3.790000 ;
      RECT  0.970000  3.870000  1.290000  4.190000 ;
      RECT  0.970000  4.270000  1.290000  4.590000 ;
      RECT  0.970000  4.670000  1.290000  4.990000 ;
      RECT  0.970000  5.070000  1.290000  5.390000 ;
      RECT  0.970000  5.470000  1.290000  5.790000 ;
      RECT  0.970000  5.870000  1.290000  6.190000 ;
      RECT  0.970000  6.270000  1.290000  6.590000 ;
      RECT  0.970000  6.670000  1.290000  6.990000 ;
      RECT  0.970000  7.070000  1.290000  7.390000 ;
      RECT  0.970000  7.470000  1.290000  7.790000 ;
      RECT  0.970000  7.870000  1.290000  8.190000 ;
      RECT  0.970000  8.270000  1.290000  8.590000 ;
      RECT  0.970000  8.670000  1.290000  8.990000 ;
      RECT  0.970000  9.070000  1.290000  9.390000 ;
      RECT  0.970000  9.470000  1.290000  9.790000 ;
      RECT  0.970000  9.870000  1.290000 10.190000 ;
      RECT  0.970000 10.270000  1.290000 10.590000 ;
      RECT  0.970000 10.670000  1.290000 10.990000 ;
      RECT  0.970000 12.210000  1.290000 12.530000 ;
      RECT  0.970000 12.610000  1.290000 12.930000 ;
      RECT  0.970000 13.010000  1.290000 13.330000 ;
      RECT  0.970000 13.410000  1.290000 13.730000 ;
      RECT  0.970000 13.810000  1.290000 14.130000 ;
      RECT  0.970000 14.210000  1.290000 14.530000 ;
      RECT  0.970000 14.610000  1.290000 14.930000 ;
      RECT  0.970000 15.010000  1.290000 15.330000 ;
      RECT  0.970000 15.410000  1.290000 15.730000 ;
      RECT  0.970000 15.810000  1.290000 16.130000 ;
      RECT  0.970000 16.210000  1.290000 16.530000 ;
      RECT  0.970000 16.610000  1.290000 16.930000 ;
      RECT  0.970000 17.010000  1.290000 17.330000 ;
      RECT  0.970000 17.410000  1.290000 17.730000 ;
      RECT  0.970000 17.810000  1.290000 18.130000 ;
      RECT  0.970000 18.210000  1.290000 18.530000 ;
      RECT  0.970000 18.610000  1.290000 18.930000 ;
      RECT  0.970000 19.010000  1.290000 19.330000 ;
      RECT  0.970000 19.410000  1.290000 19.730000 ;
      RECT  0.970000 19.810000  1.290000 20.130000 ;
      RECT  0.970000 20.210000  1.290000 20.530000 ;
      RECT  0.970000 20.610000  1.290000 20.930000 ;
      RECT  0.970000 21.010000  1.290000 21.330000 ;
      RECT  0.970000 21.410000  1.290000 21.730000 ;
      RECT  0.970000 21.810000  1.290000 22.130000 ;
      RECT  0.970000 22.210000  1.290000 22.530000 ;
      RECT  1.310000  0.240000  1.630000  0.560000 ;
      RECT  1.310000 11.100000  1.630000 11.420000 ;
      RECT  1.310000 11.780000  1.630000 12.100000 ;
      RECT  1.310000 22.640000  1.630000 22.960000 ;
      RECT  1.625000  5.670000  1.945000  5.990000 ;
      RECT  1.625000 17.210000  1.945000 17.530000 ;
      RECT  1.710000  0.240000  2.030000  0.560000 ;
      RECT  1.710000 11.100000  2.030000 11.420000 ;
      RECT  1.710000 11.780000  2.030000 12.100000 ;
      RECT  1.710000 22.640000  2.030000 22.960000 ;
      RECT  2.025000  5.670000  2.345000  5.990000 ;
      RECT  2.025000 17.210000  2.345000 17.530000 ;
      RECT  2.110000  0.240000  2.430000  0.560000 ;
      RECT  2.110000 11.100000  2.430000 11.420000 ;
      RECT  2.110000 11.780000  2.430000 12.100000 ;
      RECT  2.110000 22.640000  2.430000 22.960000 ;
      RECT  2.425000  5.670000  2.745000  5.990000 ;
      RECT  2.425000 17.210000  2.745000 17.530000 ;
      RECT  2.510000  0.240000  2.830000  0.560000 ;
      RECT  2.510000 11.100000  2.830000 11.420000 ;
      RECT  2.510000 11.780000  2.830000 12.100000 ;
      RECT  2.510000 22.640000  2.830000 22.960000 ;
      RECT  2.825000  5.670000  3.145000  5.990000 ;
      RECT  2.825000 17.210000  3.145000 17.530000 ;
      RECT  2.910000  0.240000  3.230000  0.560000 ;
      RECT  2.910000 11.100000  3.230000 11.420000 ;
      RECT  2.910000 11.780000  3.230000 12.100000 ;
      RECT  2.910000 22.640000  3.230000 22.960000 ;
      RECT  3.225000  5.670000  3.545000  5.990000 ;
      RECT  3.225000 17.210000  3.545000 17.530000 ;
      RECT  3.310000  0.240000  3.630000  0.560000 ;
      RECT  3.310000 11.100000  3.630000 11.420000 ;
      RECT  3.310000 11.780000  3.630000 12.100000 ;
      RECT  3.310000 22.640000  3.630000 22.960000 ;
      RECT  3.625000  5.670000  3.945000  5.990000 ;
      RECT  3.625000 17.210000  3.945000 17.530000 ;
      RECT  3.710000  0.240000  4.030000  0.560000 ;
      RECT  3.710000 11.100000  4.030000 11.420000 ;
      RECT  3.710000 11.780000  4.030000 12.100000 ;
      RECT  3.710000 22.640000  4.030000 22.960000 ;
      RECT  4.025000  5.670000  4.345000  5.990000 ;
      RECT  4.025000 17.210000  4.345000 17.530000 ;
      RECT  4.110000  0.240000  4.430000  0.560000 ;
      RECT  4.110000 11.100000  4.430000 11.420000 ;
      RECT  4.110000 11.780000  4.430000 12.100000 ;
      RECT  4.110000 22.640000  4.430000 22.960000 ;
      RECT  4.425000  5.670000  4.745000  5.990000 ;
      RECT  4.425000 17.210000  4.745000 17.530000 ;
      RECT  4.510000  0.240000  4.830000  0.560000 ;
      RECT  4.510000 11.100000  4.830000 11.420000 ;
      RECT  4.510000 11.780000  4.830000 12.100000 ;
      RECT  4.510000 22.640000  4.830000 22.960000 ;
      RECT  4.825000  5.670000  5.145000  5.990000 ;
      RECT  4.825000 17.210000  5.145000 17.530000 ;
      RECT  4.910000  0.240000  5.230000  0.560000 ;
      RECT  4.910000 11.100000  5.230000 11.420000 ;
      RECT  4.910000 11.780000  5.230000 12.100000 ;
      RECT  4.910000 22.640000  5.230000 22.960000 ;
      RECT  5.310000  0.240000  5.630000  0.560000 ;
      RECT  5.310000 11.100000  5.630000 11.420000 ;
      RECT  5.310000 11.780000  5.630000 12.100000 ;
      RECT  5.310000 22.640000  5.630000 22.960000 ;
      RECT  5.510000  0.870000  5.830000  1.190000 ;
      RECT  5.510000  1.270000  5.830000  1.590000 ;
      RECT  5.510000  1.670000  5.830000  1.990000 ;
      RECT  5.510000  2.070000  5.830000  2.390000 ;
      RECT  5.510000  2.470000  5.830000  2.790000 ;
      RECT  5.510000  2.870000  5.830000  3.190000 ;
      RECT  5.510000  3.270000  5.830000  3.590000 ;
      RECT  5.510000  3.670000  5.830000  3.990000 ;
      RECT  5.510000  4.070000  5.830000  4.390000 ;
      RECT  5.510000  4.470000  5.830000  4.790000 ;
      RECT  5.510000  4.870000  5.830000  5.190000 ;
      RECT  5.510000  5.270000  5.830000  5.590000 ;
      RECT  5.510000  5.670000  5.830000  5.990000 ;
      RECT  5.510000  6.070000  5.830000  6.390000 ;
      RECT  5.510000  6.470000  5.830000  6.790000 ;
      RECT  5.510000  6.870000  5.830000  7.190000 ;
      RECT  5.510000  7.270000  5.830000  7.590000 ;
      RECT  5.510000  7.670000  5.830000  7.990000 ;
      RECT  5.510000  8.070000  5.830000  8.390000 ;
      RECT  5.510000  8.470000  5.830000  8.790000 ;
      RECT  5.510000  8.870000  5.830000  9.190000 ;
      RECT  5.510000  9.270000  5.830000  9.590000 ;
      RECT  5.510000  9.670000  5.830000  9.990000 ;
      RECT  5.510000 10.070000  5.830000 10.390000 ;
      RECT  5.510000 10.470000  5.830000 10.790000 ;
      RECT  5.510000 12.410000  5.830000 12.730000 ;
      RECT  5.510000 12.810000  5.830000 13.130000 ;
      RECT  5.510000 13.210000  5.830000 13.530000 ;
      RECT  5.510000 13.610000  5.830000 13.930000 ;
      RECT  5.510000 14.010000  5.830000 14.330000 ;
      RECT  5.510000 14.410000  5.830000 14.730000 ;
      RECT  5.510000 14.810000  5.830000 15.130000 ;
      RECT  5.510000 15.210000  5.830000 15.530000 ;
      RECT  5.510000 15.610000  5.830000 15.930000 ;
      RECT  5.510000 16.010000  5.830000 16.330000 ;
      RECT  5.510000 16.410000  5.830000 16.730000 ;
      RECT  5.510000 16.810000  5.830000 17.130000 ;
      RECT  5.510000 17.210000  5.830000 17.530000 ;
      RECT  5.510000 17.610000  5.830000 17.930000 ;
      RECT  5.510000 18.010000  5.830000 18.330000 ;
      RECT  5.510000 18.410000  5.830000 18.730000 ;
      RECT  5.510000 18.810000  5.830000 19.130000 ;
      RECT  5.510000 19.210000  5.830000 19.530000 ;
      RECT  5.510000 19.610000  5.830000 19.930000 ;
      RECT  5.510000 20.010000  5.830000 20.330000 ;
      RECT  5.510000 20.410000  5.830000 20.730000 ;
      RECT  5.510000 20.810000  5.830000 21.130000 ;
      RECT  5.510000 21.210000  5.830000 21.530000 ;
      RECT  5.510000 21.610000  5.830000 21.930000 ;
      RECT  5.510000 22.010000  5.830000 22.330000 ;
      RECT  5.710000  0.240000  6.030000  0.560000 ;
      RECT  5.710000 11.100000  6.030000 11.420000 ;
      RECT  5.710000 11.780000  6.030000 12.100000 ;
      RECT  5.710000 22.640000  6.030000 22.960000 ;
      RECT  6.110000  0.240000  6.430000  0.560000 ;
      RECT  6.110000 11.100000  6.430000 11.420000 ;
      RECT  6.110000 11.780000  6.430000 12.100000 ;
      RECT  6.110000 22.640000  6.430000 22.960000 ;
      RECT  6.195000  5.670000  6.515000  5.990000 ;
      RECT  6.195000 17.210000  6.515000 17.530000 ;
      RECT  6.510000  0.240000  6.830000  0.560000 ;
      RECT  6.510000 11.100000  6.830000 11.420000 ;
      RECT  6.510000 11.780000  6.830000 12.100000 ;
      RECT  6.510000 22.640000  6.830000 22.960000 ;
      RECT  6.595000  5.670000  6.915000  5.990000 ;
      RECT  6.595000 17.210000  6.915000 17.530000 ;
      RECT  6.910000  0.240000  7.230000  0.560000 ;
      RECT  6.910000 11.100000  7.230000 11.420000 ;
      RECT  6.910000 11.780000  7.230000 12.100000 ;
      RECT  6.910000 22.640000  7.230000 22.960000 ;
      RECT  6.995000  5.670000  7.315000  5.990000 ;
      RECT  6.995000 17.210000  7.315000 17.530000 ;
      RECT  7.310000  0.240000  7.630000  0.560000 ;
      RECT  7.310000 11.100000  7.630000 11.420000 ;
      RECT  7.310000 11.780000  7.630000 12.100000 ;
      RECT  7.310000 22.640000  7.630000 22.960000 ;
      RECT  7.395000  5.670000  7.715000  5.990000 ;
      RECT  7.395000 17.210000  7.715000 17.530000 ;
      RECT  7.710000  0.240000  8.030000  0.560000 ;
      RECT  7.710000 11.100000  8.030000 11.420000 ;
      RECT  7.710000 11.780000  8.030000 12.100000 ;
      RECT  7.710000 22.640000  8.030000 22.960000 ;
      RECT  7.795000  5.670000  8.115000  5.990000 ;
      RECT  7.795000 17.210000  8.115000 17.530000 ;
      RECT  8.110000  0.240000  8.430000  0.560000 ;
      RECT  8.110000 11.100000  8.430000 11.420000 ;
      RECT  8.110000 11.780000  8.430000 12.100000 ;
      RECT  8.110000 22.640000  8.430000 22.960000 ;
      RECT  8.195000  5.670000  8.515000  5.990000 ;
      RECT  8.195000 17.210000  8.515000 17.530000 ;
      RECT  8.510000  0.240000  8.830000  0.560000 ;
      RECT  8.510000 11.100000  8.830000 11.420000 ;
      RECT  8.510000 11.780000  8.830000 12.100000 ;
      RECT  8.510000 22.640000  8.830000 22.960000 ;
      RECT  8.595000  5.670000  8.915000  5.990000 ;
      RECT  8.595000 17.210000  8.915000 17.530000 ;
      RECT  8.910000  0.240000  9.230000  0.560000 ;
      RECT  8.910000 11.100000  9.230000 11.420000 ;
      RECT  8.910000 11.780000  9.230000 12.100000 ;
      RECT  8.910000 22.640000  9.230000 22.960000 ;
      RECT  8.995000  5.670000  9.315000  5.990000 ;
      RECT  8.995000 17.210000  9.315000 17.530000 ;
      RECT  9.310000  0.240000  9.630000  0.560000 ;
      RECT  9.310000 11.100000  9.630000 11.420000 ;
      RECT  9.310000 11.780000  9.630000 12.100000 ;
      RECT  9.310000 22.640000  9.630000 22.960000 ;
      RECT  9.395000  5.670000  9.715000  5.990000 ;
      RECT  9.395000 17.210000  9.715000 17.530000 ;
      RECT  9.710000  0.240000 10.030000  0.560000 ;
      RECT  9.710000 11.100000 10.030000 11.420000 ;
      RECT  9.710000 11.780000 10.030000 12.100000 ;
      RECT  9.710000 22.640000 10.030000 22.960000 ;
      RECT 10.050000  0.670000 10.370000  0.990000 ;
      RECT 10.050000  1.070000 10.370000  1.390000 ;
      RECT 10.050000  1.470000 10.370000  1.790000 ;
      RECT 10.050000  1.870000 10.370000  2.190000 ;
      RECT 10.050000  2.270000 10.370000  2.590000 ;
      RECT 10.050000  2.670000 10.370000  2.990000 ;
      RECT 10.050000  3.070000 10.370000  3.390000 ;
      RECT 10.050000  3.470000 10.370000  3.790000 ;
      RECT 10.050000  3.870000 10.370000  4.190000 ;
      RECT 10.050000  4.270000 10.370000  4.590000 ;
      RECT 10.050000  4.670000 10.370000  4.990000 ;
      RECT 10.050000  5.070000 10.370000  5.390000 ;
      RECT 10.050000  5.470000 10.370000  5.790000 ;
      RECT 10.050000  5.870000 10.370000  6.190000 ;
      RECT 10.050000  6.270000 10.370000  6.590000 ;
      RECT 10.050000  6.670000 10.370000  6.990000 ;
      RECT 10.050000  7.070000 10.370000  7.390000 ;
      RECT 10.050000  7.470000 10.370000  7.790000 ;
      RECT 10.050000  7.870000 10.370000  8.190000 ;
      RECT 10.050000  8.270000 10.370000  8.590000 ;
      RECT 10.050000  8.670000 10.370000  8.990000 ;
      RECT 10.050000  9.070000 10.370000  9.390000 ;
      RECT 10.050000  9.470000 10.370000  9.790000 ;
      RECT 10.050000  9.870000 10.370000 10.190000 ;
      RECT 10.050000 10.270000 10.370000 10.590000 ;
      RECT 10.050000 10.670000 10.370000 10.990000 ;
      RECT 10.050000 12.210000 10.370000 12.530000 ;
      RECT 10.050000 12.610000 10.370000 12.930000 ;
      RECT 10.050000 13.010000 10.370000 13.330000 ;
      RECT 10.050000 13.410000 10.370000 13.730000 ;
      RECT 10.050000 13.810000 10.370000 14.130000 ;
      RECT 10.050000 14.210000 10.370000 14.530000 ;
      RECT 10.050000 14.610000 10.370000 14.930000 ;
      RECT 10.050000 15.010000 10.370000 15.330000 ;
      RECT 10.050000 15.410000 10.370000 15.730000 ;
      RECT 10.050000 15.810000 10.370000 16.130000 ;
      RECT 10.050000 16.210000 10.370000 16.530000 ;
      RECT 10.050000 16.610000 10.370000 16.930000 ;
      RECT 10.050000 17.010000 10.370000 17.330000 ;
      RECT 10.050000 17.410000 10.370000 17.730000 ;
      RECT 10.050000 17.810000 10.370000 18.130000 ;
      RECT 10.050000 18.210000 10.370000 18.530000 ;
      RECT 10.050000 18.610000 10.370000 18.930000 ;
      RECT 10.050000 19.010000 10.370000 19.330000 ;
      RECT 10.050000 19.410000 10.370000 19.730000 ;
      RECT 10.050000 19.810000 10.370000 20.130000 ;
      RECT 10.050000 20.210000 10.370000 20.530000 ;
      RECT 10.050000 20.610000 10.370000 20.930000 ;
      RECT 10.050000 21.010000 10.370000 21.330000 ;
      RECT 10.050000 21.410000 10.370000 21.730000 ;
      RECT 10.050000 21.810000 10.370000 22.130000 ;
      RECT 10.050000 22.210000 10.370000 22.530000 ;
      RECT 10.715000  0.465000 11.035000  0.785000 ;
      RECT 10.715000  0.865000 11.035000  1.185000 ;
      RECT 10.715000  1.265000 11.035000  1.585000 ;
      RECT 10.715000  1.665000 11.035000  1.985000 ;
      RECT 10.715000  2.065000 11.035000  2.385000 ;
      RECT 10.715000  2.465000 11.035000  2.785000 ;
      RECT 10.715000  2.865000 11.035000  3.185000 ;
      RECT 10.715000  3.265000 11.035000  3.585000 ;
      RECT 10.715000  3.665000 11.035000  3.985000 ;
      RECT 10.715000  4.065000 11.035000  4.385000 ;
      RECT 10.715000  4.465000 11.035000  4.785000 ;
      RECT 10.715000  4.865000 11.035000  5.185000 ;
      RECT 10.715000  5.265000 11.035000  5.585000 ;
      RECT 10.715000  5.665000 11.035000  5.985000 ;
      RECT 10.715000  6.065000 11.035000  6.385000 ;
      RECT 10.715000  6.465000 11.035000  6.785000 ;
      RECT 10.715000  6.865000 11.035000  7.185000 ;
      RECT 10.715000  7.265000 11.035000  7.585000 ;
      RECT 10.715000  7.665000 11.035000  7.985000 ;
      RECT 10.715000  8.065000 11.035000  8.385000 ;
      RECT 10.715000  8.465000 11.035000  8.785000 ;
      RECT 10.715000  8.865000 11.035000  9.185000 ;
      RECT 10.715000  9.265000 11.035000  9.585000 ;
      RECT 10.715000  9.665000 11.035000  9.985000 ;
      RECT 10.715000 10.065000 11.035000 10.385000 ;
      RECT 10.715000 10.465000 11.035000 10.785000 ;
      RECT 10.715000 10.865000 11.035000 11.185000 ;
      RECT 10.715000 11.265000 11.035000 11.585000 ;
      RECT 10.715000 12.005000 11.035000 12.325000 ;
      RECT 10.715000 12.405000 11.035000 12.725000 ;
      RECT 10.715000 12.805000 11.035000 13.125000 ;
      RECT 10.715000 13.205000 11.035000 13.525000 ;
      RECT 10.715000 13.605000 11.035000 13.925000 ;
      RECT 10.715000 14.005000 11.035000 14.325000 ;
      RECT 10.715000 14.405000 11.035000 14.725000 ;
      RECT 10.715000 14.805000 11.035000 15.125000 ;
      RECT 10.715000 15.205000 11.035000 15.525000 ;
      RECT 10.715000 15.605000 11.035000 15.925000 ;
      RECT 10.715000 16.005000 11.035000 16.325000 ;
      RECT 10.715000 16.405000 11.035000 16.725000 ;
      RECT 10.715000 16.805000 11.035000 17.125000 ;
      RECT 10.715000 17.205000 11.035000 17.525000 ;
      RECT 10.715000 17.605000 11.035000 17.925000 ;
      RECT 10.715000 18.005000 11.035000 18.325000 ;
      RECT 10.715000 18.405000 11.035000 18.725000 ;
      RECT 10.715000 18.805000 11.035000 19.125000 ;
      RECT 10.715000 19.205000 11.035000 19.525000 ;
      RECT 10.715000 19.605000 11.035000 19.925000 ;
      RECT 10.715000 20.005000 11.035000 20.325000 ;
      RECT 10.715000 20.405000 11.035000 20.725000 ;
      RECT 10.715000 20.805000 11.035000 21.125000 ;
      RECT 10.715000 21.205000 11.035000 21.525000 ;
      RECT 10.715000 21.605000 11.035000 21.925000 ;
      RECT 10.715000 22.005000 11.035000 22.325000 ;
      RECT 10.715000 22.405000 11.035000 22.725000 ;
      RECT 10.715000 22.805000 11.035000 23.125000 ;
      RECT 11.380000  0.670000 11.700000  0.990000 ;
      RECT 11.380000  1.070000 11.700000  1.390000 ;
      RECT 11.380000  1.470000 11.700000  1.790000 ;
      RECT 11.380000  1.870000 11.700000  2.190000 ;
      RECT 11.380000  2.270000 11.700000  2.590000 ;
      RECT 11.380000  2.670000 11.700000  2.990000 ;
      RECT 11.380000  3.070000 11.700000  3.390000 ;
      RECT 11.380000  3.470000 11.700000  3.790000 ;
      RECT 11.380000  3.870000 11.700000  4.190000 ;
      RECT 11.380000  4.270000 11.700000  4.590000 ;
      RECT 11.380000  4.670000 11.700000  4.990000 ;
      RECT 11.380000  5.070000 11.700000  5.390000 ;
      RECT 11.380000  5.470000 11.700000  5.790000 ;
      RECT 11.380000  5.870000 11.700000  6.190000 ;
      RECT 11.380000  6.270000 11.700000  6.590000 ;
      RECT 11.380000  6.670000 11.700000  6.990000 ;
      RECT 11.380000  7.070000 11.700000  7.390000 ;
      RECT 11.380000  7.470000 11.700000  7.790000 ;
      RECT 11.380000  7.870000 11.700000  8.190000 ;
      RECT 11.380000  8.270000 11.700000  8.590000 ;
      RECT 11.380000  8.670000 11.700000  8.990000 ;
      RECT 11.380000  9.070000 11.700000  9.390000 ;
      RECT 11.380000  9.470000 11.700000  9.790000 ;
      RECT 11.380000  9.870000 11.700000 10.190000 ;
      RECT 11.380000 10.270000 11.700000 10.590000 ;
      RECT 11.380000 10.670000 11.700000 10.990000 ;
      RECT 11.380000 12.210000 11.700000 12.530000 ;
      RECT 11.380000 12.610000 11.700000 12.930000 ;
      RECT 11.380000 13.010000 11.700000 13.330000 ;
      RECT 11.380000 13.410000 11.700000 13.730000 ;
      RECT 11.380000 13.810000 11.700000 14.130000 ;
      RECT 11.380000 14.210000 11.700000 14.530000 ;
      RECT 11.380000 14.610000 11.700000 14.930000 ;
      RECT 11.380000 15.010000 11.700000 15.330000 ;
      RECT 11.380000 15.410000 11.700000 15.730000 ;
      RECT 11.380000 15.810000 11.700000 16.130000 ;
      RECT 11.380000 16.210000 11.700000 16.530000 ;
      RECT 11.380000 16.610000 11.700000 16.930000 ;
      RECT 11.380000 17.010000 11.700000 17.330000 ;
      RECT 11.380000 17.410000 11.700000 17.730000 ;
      RECT 11.380000 17.810000 11.700000 18.130000 ;
      RECT 11.380000 18.210000 11.700000 18.530000 ;
      RECT 11.380000 18.610000 11.700000 18.930000 ;
      RECT 11.380000 19.010000 11.700000 19.330000 ;
      RECT 11.380000 19.410000 11.700000 19.730000 ;
      RECT 11.380000 19.810000 11.700000 20.130000 ;
      RECT 11.380000 20.210000 11.700000 20.530000 ;
      RECT 11.380000 20.610000 11.700000 20.930000 ;
      RECT 11.380000 21.010000 11.700000 21.330000 ;
      RECT 11.380000 21.410000 11.700000 21.730000 ;
      RECT 11.380000 21.810000 11.700000 22.130000 ;
      RECT 11.380000 22.210000 11.700000 22.530000 ;
      RECT 11.720000  0.240000 12.040000  0.560000 ;
      RECT 11.720000 11.100000 12.040000 11.420000 ;
      RECT 11.720000 11.780000 12.040000 12.100000 ;
      RECT 11.720000 22.640000 12.040000 22.960000 ;
      RECT 12.035000  5.670000 12.355000  5.990000 ;
      RECT 12.035000 17.210000 12.355000 17.530000 ;
      RECT 12.120000  0.240000 12.440000  0.560000 ;
      RECT 12.120000 11.100000 12.440000 11.420000 ;
      RECT 12.120000 11.780000 12.440000 12.100000 ;
      RECT 12.120000 22.640000 12.440000 22.960000 ;
      RECT 12.435000  5.670000 12.755000  5.990000 ;
      RECT 12.435000 17.210000 12.755000 17.530000 ;
      RECT 12.520000  0.240000 12.840000  0.560000 ;
      RECT 12.520000 11.100000 12.840000 11.420000 ;
      RECT 12.520000 11.780000 12.840000 12.100000 ;
      RECT 12.520000 22.640000 12.840000 22.960000 ;
      RECT 12.835000  5.670000 13.155000  5.990000 ;
      RECT 12.835000 17.210000 13.155000 17.530000 ;
      RECT 12.920000  0.240000 13.240000  0.560000 ;
      RECT 12.920000 11.100000 13.240000 11.420000 ;
      RECT 12.920000 11.780000 13.240000 12.100000 ;
      RECT 12.920000 22.640000 13.240000 22.960000 ;
      RECT 13.235000  5.670000 13.555000  5.990000 ;
      RECT 13.235000 17.210000 13.555000 17.530000 ;
      RECT 13.320000  0.240000 13.640000  0.560000 ;
      RECT 13.320000 11.100000 13.640000 11.420000 ;
      RECT 13.320000 11.780000 13.640000 12.100000 ;
      RECT 13.320000 22.640000 13.640000 22.960000 ;
      RECT 13.635000  5.670000 13.955000  5.990000 ;
      RECT 13.635000 17.210000 13.955000 17.530000 ;
      RECT 13.720000  0.240000 14.040000  0.560000 ;
      RECT 13.720000 11.100000 14.040000 11.420000 ;
      RECT 13.720000 11.780000 14.040000 12.100000 ;
      RECT 13.720000 22.640000 14.040000 22.960000 ;
      RECT 14.035000  5.670000 14.355000  5.990000 ;
      RECT 14.035000 17.210000 14.355000 17.530000 ;
      RECT 14.120000  0.240000 14.440000  0.560000 ;
      RECT 14.120000 11.100000 14.440000 11.420000 ;
      RECT 14.120000 11.780000 14.440000 12.100000 ;
      RECT 14.120000 22.640000 14.440000 22.960000 ;
      RECT 14.435000  5.670000 14.755000  5.990000 ;
      RECT 14.435000 17.210000 14.755000 17.530000 ;
      RECT 14.520000  0.240000 14.840000  0.560000 ;
      RECT 14.520000 11.100000 14.840000 11.420000 ;
      RECT 14.520000 11.780000 14.840000 12.100000 ;
      RECT 14.520000 22.640000 14.840000 22.960000 ;
      RECT 14.835000  5.670000 15.155000  5.990000 ;
      RECT 14.835000 17.210000 15.155000 17.530000 ;
      RECT 14.920000  0.240000 15.240000  0.560000 ;
      RECT 14.920000 11.100000 15.240000 11.420000 ;
      RECT 14.920000 11.780000 15.240000 12.100000 ;
      RECT 14.920000 22.640000 15.240000 22.960000 ;
      RECT 15.235000  5.670000 15.555000  5.990000 ;
      RECT 15.235000 17.210000 15.555000 17.530000 ;
      RECT 15.320000  0.240000 15.640000  0.560000 ;
      RECT 15.320000 11.100000 15.640000 11.420000 ;
      RECT 15.320000 11.780000 15.640000 12.100000 ;
      RECT 15.320000 22.640000 15.640000 22.960000 ;
      RECT 15.720000  0.240000 16.040000  0.560000 ;
      RECT 15.720000 11.100000 16.040000 11.420000 ;
      RECT 15.720000 11.780000 16.040000 12.100000 ;
      RECT 15.720000 22.640000 16.040000 22.960000 ;
      RECT 15.920000  0.870000 16.240000  1.190000 ;
      RECT 15.920000  1.270000 16.240000  1.590000 ;
      RECT 15.920000  1.670000 16.240000  1.990000 ;
      RECT 15.920000  2.070000 16.240000  2.390000 ;
      RECT 15.920000  2.470000 16.240000  2.790000 ;
      RECT 15.920000  2.870000 16.240000  3.190000 ;
      RECT 15.920000  3.270000 16.240000  3.590000 ;
      RECT 15.920000  3.670000 16.240000  3.990000 ;
      RECT 15.920000  4.070000 16.240000  4.390000 ;
      RECT 15.920000  4.470000 16.240000  4.790000 ;
      RECT 15.920000  4.870000 16.240000  5.190000 ;
      RECT 15.920000  5.270000 16.240000  5.590000 ;
      RECT 15.920000  5.670000 16.240000  5.990000 ;
      RECT 15.920000  6.070000 16.240000  6.390000 ;
      RECT 15.920000  6.470000 16.240000  6.790000 ;
      RECT 15.920000  6.870000 16.240000  7.190000 ;
      RECT 15.920000  7.270000 16.240000  7.590000 ;
      RECT 15.920000  7.670000 16.240000  7.990000 ;
      RECT 15.920000  8.070000 16.240000  8.390000 ;
      RECT 15.920000  8.470000 16.240000  8.790000 ;
      RECT 15.920000  8.870000 16.240000  9.190000 ;
      RECT 15.920000  9.270000 16.240000  9.590000 ;
      RECT 15.920000  9.670000 16.240000  9.990000 ;
      RECT 15.920000 10.070000 16.240000 10.390000 ;
      RECT 15.920000 10.470000 16.240000 10.790000 ;
      RECT 15.920000 12.410000 16.240000 12.730000 ;
      RECT 15.920000 12.810000 16.240000 13.130000 ;
      RECT 15.920000 13.210000 16.240000 13.530000 ;
      RECT 15.920000 13.610000 16.240000 13.930000 ;
      RECT 15.920000 14.010000 16.240000 14.330000 ;
      RECT 15.920000 14.410000 16.240000 14.730000 ;
      RECT 15.920000 14.810000 16.240000 15.130000 ;
      RECT 15.920000 15.210000 16.240000 15.530000 ;
      RECT 15.920000 15.610000 16.240000 15.930000 ;
      RECT 15.920000 16.010000 16.240000 16.330000 ;
      RECT 15.920000 16.410000 16.240000 16.730000 ;
      RECT 15.920000 16.810000 16.240000 17.130000 ;
      RECT 15.920000 17.210000 16.240000 17.530000 ;
      RECT 15.920000 17.610000 16.240000 17.930000 ;
      RECT 15.920000 18.010000 16.240000 18.330000 ;
      RECT 15.920000 18.410000 16.240000 18.730000 ;
      RECT 15.920000 18.810000 16.240000 19.130000 ;
      RECT 15.920000 19.210000 16.240000 19.530000 ;
      RECT 15.920000 19.610000 16.240000 19.930000 ;
      RECT 15.920000 20.010000 16.240000 20.330000 ;
      RECT 15.920000 20.410000 16.240000 20.730000 ;
      RECT 15.920000 20.810000 16.240000 21.130000 ;
      RECT 15.920000 21.210000 16.240000 21.530000 ;
      RECT 15.920000 21.610000 16.240000 21.930000 ;
      RECT 15.920000 22.010000 16.240000 22.330000 ;
      RECT 16.120000  0.240000 16.440000  0.560000 ;
      RECT 16.120000 11.100000 16.440000 11.420000 ;
      RECT 16.120000 11.780000 16.440000 12.100000 ;
      RECT 16.120000 22.640000 16.440000 22.960000 ;
      RECT 16.520000  0.240000 16.840000  0.560000 ;
      RECT 16.520000 11.100000 16.840000 11.420000 ;
      RECT 16.520000 11.780000 16.840000 12.100000 ;
      RECT 16.520000 22.640000 16.840000 22.960000 ;
      RECT 16.605000  5.670000 16.925000  5.990000 ;
      RECT 16.605000 17.210000 16.925000 17.530000 ;
      RECT 16.920000  0.240000 17.240000  0.560000 ;
      RECT 16.920000 11.100000 17.240000 11.420000 ;
      RECT 16.920000 11.780000 17.240000 12.100000 ;
      RECT 16.920000 22.640000 17.240000 22.960000 ;
      RECT 17.005000  5.670000 17.325000  5.990000 ;
      RECT 17.005000 17.210000 17.325000 17.530000 ;
      RECT 17.320000  0.240000 17.640000  0.560000 ;
      RECT 17.320000 11.100000 17.640000 11.420000 ;
      RECT 17.320000 11.780000 17.640000 12.100000 ;
      RECT 17.320000 22.640000 17.640000 22.960000 ;
      RECT 17.405000  5.670000 17.725000  5.990000 ;
      RECT 17.405000 17.210000 17.725000 17.530000 ;
      RECT 17.720000  0.240000 18.040000  0.560000 ;
      RECT 17.720000 11.100000 18.040000 11.420000 ;
      RECT 17.720000 11.780000 18.040000 12.100000 ;
      RECT 17.720000 22.640000 18.040000 22.960000 ;
      RECT 17.805000  5.670000 18.125000  5.990000 ;
      RECT 17.805000 17.210000 18.125000 17.530000 ;
      RECT 18.120000  0.240000 18.440000  0.560000 ;
      RECT 18.120000 11.100000 18.440000 11.420000 ;
      RECT 18.120000 11.780000 18.440000 12.100000 ;
      RECT 18.120000 22.640000 18.440000 22.960000 ;
      RECT 18.205000  5.670000 18.525000  5.990000 ;
      RECT 18.205000 17.210000 18.525000 17.530000 ;
      RECT 18.520000  0.240000 18.840000  0.560000 ;
      RECT 18.520000 11.100000 18.840000 11.420000 ;
      RECT 18.520000 11.780000 18.840000 12.100000 ;
      RECT 18.520000 22.640000 18.840000 22.960000 ;
      RECT 18.605000  5.670000 18.925000  5.990000 ;
      RECT 18.605000 17.210000 18.925000 17.530000 ;
      RECT 18.920000  0.240000 19.240000  0.560000 ;
      RECT 18.920000 11.100000 19.240000 11.420000 ;
      RECT 18.920000 11.780000 19.240000 12.100000 ;
      RECT 18.920000 22.640000 19.240000 22.960000 ;
      RECT 19.005000  5.670000 19.325000  5.990000 ;
      RECT 19.005000 17.210000 19.325000 17.530000 ;
      RECT 19.320000  0.240000 19.640000  0.560000 ;
      RECT 19.320000 11.100000 19.640000 11.420000 ;
      RECT 19.320000 11.780000 19.640000 12.100000 ;
      RECT 19.320000 22.640000 19.640000 22.960000 ;
      RECT 19.405000  5.670000 19.725000  5.990000 ;
      RECT 19.405000 17.210000 19.725000 17.530000 ;
      RECT 19.720000  0.240000 20.040000  0.560000 ;
      RECT 19.720000 11.100000 20.040000 11.420000 ;
      RECT 19.720000 11.780000 20.040000 12.100000 ;
      RECT 19.720000 22.640000 20.040000 22.960000 ;
      RECT 19.805000  5.670000 20.125000  5.990000 ;
      RECT 19.805000 17.210000 20.125000 17.530000 ;
      RECT 20.120000  0.240000 20.440000  0.560000 ;
      RECT 20.120000 11.100000 20.440000 11.420000 ;
      RECT 20.120000 11.780000 20.440000 12.100000 ;
      RECT 20.120000 22.640000 20.440000 22.960000 ;
      RECT 20.460000  0.670000 20.780000  0.990000 ;
      RECT 20.460000  1.070000 20.780000  1.390000 ;
      RECT 20.460000  1.470000 20.780000  1.790000 ;
      RECT 20.460000  1.870000 20.780000  2.190000 ;
      RECT 20.460000  2.270000 20.780000  2.590000 ;
      RECT 20.460000  2.670000 20.780000  2.990000 ;
      RECT 20.460000  3.070000 20.780000  3.390000 ;
      RECT 20.460000  3.470000 20.780000  3.790000 ;
      RECT 20.460000  3.870000 20.780000  4.190000 ;
      RECT 20.460000  4.270000 20.780000  4.590000 ;
      RECT 20.460000  4.670000 20.780000  4.990000 ;
      RECT 20.460000  5.070000 20.780000  5.390000 ;
      RECT 20.460000  5.470000 20.780000  5.790000 ;
      RECT 20.460000  5.870000 20.780000  6.190000 ;
      RECT 20.460000  6.270000 20.780000  6.590000 ;
      RECT 20.460000  6.670000 20.780000  6.990000 ;
      RECT 20.460000  7.070000 20.780000  7.390000 ;
      RECT 20.460000  7.470000 20.780000  7.790000 ;
      RECT 20.460000  7.870000 20.780000  8.190000 ;
      RECT 20.460000  8.270000 20.780000  8.590000 ;
      RECT 20.460000  8.670000 20.780000  8.990000 ;
      RECT 20.460000  9.070000 20.780000  9.390000 ;
      RECT 20.460000  9.470000 20.780000  9.790000 ;
      RECT 20.460000  9.870000 20.780000 10.190000 ;
      RECT 20.460000 10.270000 20.780000 10.590000 ;
      RECT 20.460000 10.670000 20.780000 10.990000 ;
      RECT 20.460000 12.210000 20.780000 12.530000 ;
      RECT 20.460000 12.610000 20.780000 12.930000 ;
      RECT 20.460000 13.010000 20.780000 13.330000 ;
      RECT 20.460000 13.410000 20.780000 13.730000 ;
      RECT 20.460000 13.810000 20.780000 14.130000 ;
      RECT 20.460000 14.210000 20.780000 14.530000 ;
      RECT 20.460000 14.610000 20.780000 14.930000 ;
      RECT 20.460000 15.010000 20.780000 15.330000 ;
      RECT 20.460000 15.410000 20.780000 15.730000 ;
      RECT 20.460000 15.810000 20.780000 16.130000 ;
      RECT 20.460000 16.210000 20.780000 16.530000 ;
      RECT 20.460000 16.610000 20.780000 16.930000 ;
      RECT 20.460000 17.010000 20.780000 17.330000 ;
      RECT 20.460000 17.410000 20.780000 17.730000 ;
      RECT 20.460000 17.810000 20.780000 18.130000 ;
      RECT 20.460000 18.210000 20.780000 18.530000 ;
      RECT 20.460000 18.610000 20.780000 18.930000 ;
      RECT 20.460000 19.010000 20.780000 19.330000 ;
      RECT 20.460000 19.410000 20.780000 19.730000 ;
      RECT 20.460000 19.810000 20.780000 20.130000 ;
      RECT 20.460000 20.210000 20.780000 20.530000 ;
      RECT 20.460000 20.610000 20.780000 20.930000 ;
      RECT 20.460000 21.010000 20.780000 21.330000 ;
      RECT 20.460000 21.410000 20.780000 21.730000 ;
      RECT 20.460000 21.810000 20.780000 22.130000 ;
      RECT 20.460000 22.210000 20.780000 22.530000 ;
      RECT 21.125000  0.465000 21.445000  0.785000 ;
      RECT 21.125000  0.865000 21.445000  1.185000 ;
      RECT 21.125000  1.265000 21.445000  1.585000 ;
      RECT 21.125000  1.665000 21.445000  1.985000 ;
      RECT 21.125000  2.065000 21.445000  2.385000 ;
      RECT 21.125000  2.465000 21.445000  2.785000 ;
      RECT 21.125000  2.865000 21.445000  3.185000 ;
      RECT 21.125000  3.265000 21.445000  3.585000 ;
      RECT 21.125000  3.665000 21.445000  3.985000 ;
      RECT 21.125000  4.065000 21.445000  4.385000 ;
      RECT 21.125000  4.465000 21.445000  4.785000 ;
      RECT 21.125000  4.865000 21.445000  5.185000 ;
      RECT 21.125000  5.265000 21.445000  5.585000 ;
      RECT 21.125000  5.665000 21.445000  5.985000 ;
      RECT 21.125000  6.065000 21.445000  6.385000 ;
      RECT 21.125000  6.465000 21.445000  6.785000 ;
      RECT 21.125000  6.865000 21.445000  7.185000 ;
      RECT 21.125000  7.265000 21.445000  7.585000 ;
      RECT 21.125000  7.665000 21.445000  7.985000 ;
      RECT 21.125000  8.065000 21.445000  8.385000 ;
      RECT 21.125000  8.465000 21.445000  8.785000 ;
      RECT 21.125000  8.865000 21.445000  9.185000 ;
      RECT 21.125000  9.265000 21.445000  9.585000 ;
      RECT 21.125000  9.665000 21.445000  9.985000 ;
      RECT 21.125000 10.065000 21.445000 10.385000 ;
      RECT 21.125000 10.465000 21.445000 10.785000 ;
      RECT 21.125000 10.865000 21.445000 11.185000 ;
      RECT 21.125000 11.265000 21.445000 11.585000 ;
      RECT 21.125000 12.005000 21.445000 12.325000 ;
      RECT 21.125000 12.405000 21.445000 12.725000 ;
      RECT 21.125000 12.805000 21.445000 13.125000 ;
      RECT 21.125000 13.205000 21.445000 13.525000 ;
      RECT 21.125000 13.605000 21.445000 13.925000 ;
      RECT 21.125000 14.005000 21.445000 14.325000 ;
      RECT 21.125000 14.405000 21.445000 14.725000 ;
      RECT 21.125000 14.805000 21.445000 15.125000 ;
      RECT 21.125000 15.205000 21.445000 15.525000 ;
      RECT 21.125000 15.605000 21.445000 15.925000 ;
      RECT 21.125000 16.005000 21.445000 16.325000 ;
      RECT 21.125000 16.405000 21.445000 16.725000 ;
      RECT 21.125000 16.805000 21.445000 17.125000 ;
      RECT 21.125000 17.205000 21.445000 17.525000 ;
      RECT 21.125000 17.605000 21.445000 17.925000 ;
      RECT 21.125000 18.005000 21.445000 18.325000 ;
      RECT 21.125000 18.405000 21.445000 18.725000 ;
      RECT 21.125000 18.805000 21.445000 19.125000 ;
      RECT 21.125000 19.205000 21.445000 19.525000 ;
      RECT 21.125000 19.605000 21.445000 19.925000 ;
      RECT 21.125000 20.005000 21.445000 20.325000 ;
      RECT 21.125000 20.405000 21.445000 20.725000 ;
      RECT 21.125000 20.805000 21.445000 21.125000 ;
      RECT 21.125000 21.205000 21.445000 21.525000 ;
      RECT 21.125000 21.605000 21.445000 21.925000 ;
      RECT 21.125000 22.005000 21.445000 22.325000 ;
      RECT 21.125000 22.405000 21.445000 22.725000 ;
      RECT 21.125000 22.805000 21.445000 23.125000 ;
  END
END sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhvtop
END LIBRARY
