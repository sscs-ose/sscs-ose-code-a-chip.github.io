* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 9
.param
+ sky130_fd_pr__nfet_03v3_nvt__toxe_mult = 0.948
+ sky130_fd_pr__nfet_03v3_nvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_03v3_nvt__overlap_mult = 0.40927
+ sky130_fd_pr__nfet_03v3_nvt__ajunction_mult = 0.56418
+ sky130_fd_pr__nfet_03v3_nvt__pjunction_mult = 0.84099
+ sky130_fd_pr__nfet_03v3_nvt__lint_diff = 1.7325e-8
+ sky130_fd_pr__nfet_03v3_nvt__wint_diff = -3.2175e-8
+ sky130_fd_pr__nfet_03v3_nvt__dlc_diff = 3.0000e-8
+ sky130_fd_pr__nfet_03v3_nvt__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 000, W = 10.0, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_0 = -0.0010542
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_0 = -0.026492
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0 = -1.0339
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0 = -0.047264
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_0 = 0.00016819
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0 = -3949.2
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_0 = 4.2013e-19
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_0 = 5.9282e-11
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 001, W = 1.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_1 = 8.318e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_1 = -0.020875
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_1 = -0.0056301
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1 = -1.707
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1 = -0.060897
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_1 = -0.0028636
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1 = -14012.0
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_1 = 4.2893e-19
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 002, W = 1.0, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_2 = 1.0603e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_2 = 4.1221e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_2 = -0.00080074
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2 = -0.47778
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2 = -0.050539
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_2 = -0.00039963
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2 = -12436.0
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_2 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 003, W = 4.0, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_3 = 7.9696e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_3 = 5.7902e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_3 = -0.0026756
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_3 = -0.023644
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3 = -0.95532
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3 = -0.048464
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_3 = 0.0011558
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3 = -6147.9
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_3 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 004, W = 0.42, L = 0.5
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_4 = 1.7046e-19
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_4 = 3.9478e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_4 = 0.032977
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_4 = 0.0069451
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4 = -1.6941
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4 = -0.083671
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_4 = -0.0011543
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4 = -12626.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 005, W = 0.42, L = 0.6
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_5 = 0.0089834
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5 = -11481.0
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_5 = 1.7135e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_5 = 4.1927e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_5 = 0.0029293
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5 = -1.5761
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5 = -0.0016017
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 006, W = 0.42, L = 0.8
* -------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6 = -0.73851
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6 = -0.014966
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_6 = 0.0066129
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6 = -9425.6
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_6 = 1.5395e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_6 = 6.8955e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_6 = 0.0030242
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 007, W = 0.7, L = 0.5
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_7 = -0.0078507
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_7 = -0.0030712
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7 = -1.5397
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7 = -0.053605
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_7 = -0.000432
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7 = -14226.0
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_7 = 1.2313e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_7 = 6.9284e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_7 = 0.0
*
* sky130_fd_pr__nfet_03v3_nvt, Bin 008, W = 0.7, L = 0.6
* ------------------------------------
+ sky130_fd_pr__nfet_03v3_nvt__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_8 = 0.0019101
+ sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8 = -0.52333
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8 = -0.057025
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_8 = 0.00086474
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8 = -12780.0
+ sky130_fd_pr__nfet_03v3_nvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_8 = 1.3078e-18
+ sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_8 = 4.5353e-11
+ sky130_fd_pr__nfet_03v3_nvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8 = 0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"
