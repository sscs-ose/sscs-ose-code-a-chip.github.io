magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< nwell >>
rect -246 -973 246 973
<< pmos >>
rect -50 554 50 754
rect -50 118 50 318
rect -50 -318 50 -118
rect -50 -754 50 -554
<< pdiff >>
rect -108 742 -50 754
rect -108 566 -96 742
rect -62 566 -50 742
rect -108 554 -50 566
rect 50 742 108 754
rect 50 566 62 742
rect 96 566 108 742
rect 50 554 108 566
rect -108 306 -50 318
rect -108 130 -96 306
rect -62 130 -50 306
rect -108 118 -50 130
rect 50 306 108 318
rect 50 130 62 306
rect 96 130 108 306
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -306 -96 -130
rect -62 -306 -50 -130
rect -108 -318 -50 -306
rect 50 -130 108 -118
rect 50 -306 62 -130
rect 96 -306 108 -130
rect 50 -318 108 -306
rect -108 -566 -50 -554
rect -108 -742 -96 -566
rect -62 -742 -50 -566
rect -108 -754 -50 -742
rect 50 -566 108 -554
rect 50 -742 62 -566
rect 96 -742 108 -566
rect 50 -754 108 -742
<< pdiffc >>
rect -96 566 -62 742
rect 62 566 96 742
rect -96 130 -62 306
rect 62 130 96 306
rect -96 -306 -62 -130
rect 62 -306 96 -130
rect -96 -742 -62 -566
rect 62 -742 96 -566
<< nsubdiff >>
rect -210 903 -114 937
rect 114 903 210 937
rect -210 841 -176 903
rect 176 841 210 903
rect -210 -903 -176 -841
rect 176 -903 210 -841
rect -210 -937 -114 -903
rect 114 -937 210 -903
<< nsubdiffcont >>
rect -114 903 114 937
rect -210 -841 -176 841
rect 176 -841 210 841
rect -114 -937 114 -903
<< poly >>
rect -50 835 50 851
rect -50 801 -34 835
rect 34 801 50 835
rect -50 754 50 801
rect -50 507 50 554
rect -50 473 -34 507
rect 34 473 50 507
rect -50 457 50 473
rect -50 399 50 415
rect -50 365 -34 399
rect 34 365 50 399
rect -50 318 50 365
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -365 50 -318
rect -50 -399 -34 -365
rect 34 -399 50 -365
rect -50 -415 50 -399
rect -50 -473 50 -457
rect -50 -507 -34 -473
rect 34 -507 50 -473
rect -50 -554 50 -507
rect -50 -801 50 -754
rect -50 -835 -34 -801
rect 34 -835 50 -801
rect -50 -851 50 -835
<< polycont >>
rect -34 801 34 835
rect -34 473 34 507
rect -34 365 34 399
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -399 34 -365
rect -34 -507 34 -473
rect -34 -835 34 -801
<< locali >>
rect -210 903 -114 937
rect 114 903 210 937
rect -210 841 -176 903
rect 176 841 210 903
rect -50 801 -34 835
rect 34 801 50 835
rect -96 742 -62 758
rect -96 550 -62 566
rect 62 742 96 758
rect 62 550 96 566
rect -50 473 -34 507
rect 34 473 50 507
rect -50 365 -34 399
rect 34 365 50 399
rect -96 306 -62 322
rect -96 114 -62 130
rect 62 306 96 322
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -322 -62 -306
rect 62 -130 96 -114
rect 62 -322 96 -306
rect -50 -399 -34 -365
rect 34 -399 50 -365
rect -50 -507 -34 -473
rect 34 -507 50 -473
rect -96 -566 -62 -550
rect -96 -758 -62 -742
rect 62 -566 96 -550
rect 62 -758 96 -742
rect -50 -835 -34 -801
rect 34 -835 50 -801
rect -210 -903 -176 -841
rect 176 -903 210 -841
rect -210 -937 -114 -903
rect 114 -937 210 -903
<< viali >>
rect -34 801 34 835
rect -96 566 -62 742
rect 62 566 96 742
rect -34 473 34 507
rect -34 365 34 399
rect -96 130 -62 306
rect 62 130 96 306
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -306 -62 -130
rect 62 -306 96 -130
rect -34 -399 34 -365
rect -34 -507 34 -473
rect -96 -742 -62 -566
rect 62 -742 96 -566
rect -34 -835 34 -801
<< metal1 >>
rect -46 835 46 841
rect -46 801 -34 835
rect 34 801 46 835
rect -46 795 46 801
rect -102 742 -56 754
rect -102 566 -96 742
rect -62 566 -56 742
rect -102 554 -56 566
rect 56 742 102 754
rect 56 566 62 742
rect 96 566 102 742
rect 56 554 102 566
rect -46 507 46 513
rect -46 473 -34 507
rect 34 473 46 507
rect -46 467 46 473
rect -46 399 46 405
rect -46 365 -34 399
rect 34 365 46 399
rect -46 359 46 365
rect -102 306 -56 318
rect -102 130 -96 306
rect -62 130 -56 306
rect -102 118 -56 130
rect 56 306 102 318
rect 56 130 62 306
rect 96 130 102 306
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -306 -96 -130
rect -62 -306 -56 -130
rect -102 -318 -56 -306
rect 56 -130 102 -118
rect 56 -306 62 -130
rect 96 -306 102 -130
rect 56 -318 102 -306
rect -46 -365 46 -359
rect -46 -399 -34 -365
rect 34 -399 46 -365
rect -46 -405 46 -399
rect -46 -473 46 -467
rect -46 -507 -34 -473
rect 34 -507 46 -473
rect -46 -513 46 -507
rect -102 -566 -56 -554
rect -102 -742 -96 -566
rect -62 -742 -56 -566
rect -102 -754 -56 -742
rect 56 -566 102 -554
rect 56 -742 62 -566
rect 96 -742 102 -566
rect 56 -754 102 -742
rect -46 -801 46 -795
rect -46 -835 -34 -801
rect 34 -835 46 -801
rect -46 -841 46 -835
<< labels >>
rlabel nsubdiffcont 0 -920 0 -920 0 B
port 14 nsew
rlabel pdiffc -79 -654 -79 -654 0 D0
port 15 nsew
rlabel pdiffc 79 -654 79 -654 0 S0
port 16 nsew
rlabel polycont 0 -490 0 -490 0 G0
port 17 nsew
rlabel pdiffc -79 -218 -79 -218 0 D1
port 18 nsew
rlabel pdiffc 79 -218 79 -218 0 S1
port 19 nsew
rlabel polycont 0 -54 0 -54 0 G1
port 20 nsew
rlabel pdiffc -79 218 -79 218 0 D2
port 21 nsew
rlabel pdiffc 79 218 79 218 0 S2
port 22 nsew
rlabel polycont 0 382 0 382 0 G2
port 23 nsew
rlabel pdiffc -79 654 -79 654 0 D3
port 24 nsew
rlabel pdiffc 79 654 79 654 0 S3
port 25 nsew
rlabel polycont 0 818 0 818 0 G3
port 26 nsew
<< properties >>
string FIXED_BBOX -193 -920 193 920
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.5 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 4
<< end >>
