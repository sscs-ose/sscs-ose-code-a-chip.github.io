magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -307 -4782 307 4782
<< psubdiff >>
rect -271 4712 -175 4746
rect 175 4712 271 4746
rect -271 4650 -237 4712
rect 237 4650 271 4712
rect -271 -4712 -237 -4650
rect 237 -4712 271 -4650
rect -271 -4746 -175 -4712
rect 175 -4746 271 -4712
<< psubdiffcont >>
rect -175 4712 175 4746
rect -271 -4650 -237 4650
rect 237 -4650 271 4650
rect -175 -4746 175 -4712
<< xpolycontact >>
rect -141 4184 141 4616
rect -141 -4616 141 -4184
<< ppolyres >>
rect -141 -4184 141 4184
<< locali >>
rect -271 4712 -175 4746
rect 175 4712 271 4746
rect -271 4650 -237 4712
rect 237 4650 271 4712
rect -271 -4712 -237 -4650
rect 237 -4712 271 -4650
rect -271 -4746 -175 -4712
rect 175 -4746 271 -4712
<< viali >>
rect -125 4201 125 4598
rect -125 -4598 125 -4201
<< metal1 >>
rect -131 4598 131 4610
rect -131 4201 -125 4598
rect 125 4201 131 4598
rect -131 4189 131 4201
rect -131 -4201 131 -4189
rect -131 -4598 -125 -4201
rect 125 -4598 131 -4201
rect -131 -4610 131 -4598
<< labels >>
rlabel psubdiffcont 0 -4729 0 -4729 0 B
port 7 nsew
rlabel xpolycontact 0 4581 0 4581 0 R1
port 8 nsew
rlabel xpolycontact 0 -4581 0 -4581 0 R2
port 9 nsew
<< properties >>
string FIXED_BBOX -254 -4729 254 4729
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 42.0 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 319.8 val 9.802k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1 mult 1
<< end >>
