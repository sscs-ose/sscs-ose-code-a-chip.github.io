* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
*
* model corner
* , Bin 000, W = 30.0, L = 1.0
* ----------------------------
.param
+ sky130_fd_pr__nfet_20v0_zvt__rdrift_mult = 0.694573191726037
+ sky130_fd_pr__nfet_20v0_zvt__hvvsat_mult = 1.0
+ sky130_fd_pr__nfet_20v0_zvt__vth0_diff = -0.37085
+ sky130_fd_pr__nfet_20v0_zvt__k2_diff = 0.0
+ sky130_fd_pr__nfet_20v0_zvt__lint_diff= 0.0
+ sky130_fd_pr__nfet_20v0_zvt__u0_diff = 1.5631e-1
+ sky130_fd_pr__nfet_20v0_zvt__agidl_diff = 1.4e-14
+ sky130_fd_pr__nfet_20v0_zvt__vsat_diff = 0.0
+ sky130_fd_pr__nfet_20v0_zvt__ags_diff = 0.0
+ sky130_fd_pr__nfet_20v0_zvt__keta_diff = 0.0
+ n20zvtvh1defet_js_mult_pmc = 10.0
.include "sky130_fd_pr__nfet_20v0_zvt__subcircuit.pm3.spice"
