# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_npn_05v5_W1p00L1p00
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_npn_05v5_W1p00L1p00 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.620000 BY  8.620000 ;
  OBS
    LAYER li1 ;
      RECT 0.630000 0.630000 7.990000 0.960000 ;
      RECT 0.630000 0.960000 0.960000 7.660000 ;
      RECT 0.630000 7.660000 7.990000 7.990000 ;
      RECT 2.640000 2.640000 5.980000 2.970000 ;
      RECT 2.640000 2.970000 2.970000 5.650000 ;
      RECT 2.640000 5.650000 5.980000 5.980000 ;
      RECT 3.805000 3.805000 4.815000 4.815000 ;
      RECT 5.650000 2.970000 5.980000 5.650000 ;
      RECT 7.660000 0.960000 7.990000 7.660000 ;
    LAYER mcon ;
      RECT 0.710000 0.710000 0.880000 0.880000 ;
      RECT 0.710000 1.165000 0.880000 1.335000 ;
      RECT 0.710000 1.525000 0.880000 1.695000 ;
      RECT 0.710000 1.885000 0.880000 2.055000 ;
      RECT 0.710000 2.245000 0.880000 2.415000 ;
      RECT 0.710000 2.605000 0.880000 2.775000 ;
      RECT 0.710000 2.965000 0.880000 3.135000 ;
      RECT 0.710000 3.325000 0.880000 3.495000 ;
      RECT 0.710000 3.685000 0.880000 3.855000 ;
      RECT 0.710000 4.045000 0.880000 4.215000 ;
      RECT 0.710000 4.405000 0.880000 4.575000 ;
      RECT 0.710000 4.765000 0.880000 4.935000 ;
      RECT 0.710000 5.125000 0.880000 5.295000 ;
      RECT 0.710000 5.485000 0.880000 5.655000 ;
      RECT 0.710000 5.845000 0.880000 6.015000 ;
      RECT 0.710000 6.205000 0.880000 6.375000 ;
      RECT 0.710000 6.565000 0.880000 6.735000 ;
      RECT 0.710000 6.925000 0.880000 7.095000 ;
      RECT 0.710000 7.285000 0.880000 7.455000 ;
      RECT 0.710000 7.740000 0.880000 7.910000 ;
      RECT 1.165000 0.710000 1.335000 0.880000 ;
      RECT 1.165000 7.740000 1.335000 7.910000 ;
      RECT 1.525000 0.710000 1.695000 0.880000 ;
      RECT 1.525000 7.740000 1.695000 7.910000 ;
      RECT 1.885000 0.710000 2.055000 0.880000 ;
      RECT 1.885000 7.740000 2.055000 7.910000 ;
      RECT 2.245000 0.710000 2.415000 0.880000 ;
      RECT 2.245000 7.740000 2.415000 7.910000 ;
      RECT 2.605000 0.710000 2.775000 0.880000 ;
      RECT 2.605000 7.740000 2.775000 7.910000 ;
      RECT 2.720000 2.720000 2.890000 2.890000 ;
      RECT 2.720000 3.145000 2.890000 3.315000 ;
      RECT 2.720000 3.505000 2.890000 3.675000 ;
      RECT 2.720000 3.865000 2.890000 4.035000 ;
      RECT 2.720000 4.225000 2.890000 4.395000 ;
      RECT 2.720000 4.585000 2.890000 4.755000 ;
      RECT 2.720000 4.945000 2.890000 5.115000 ;
      RECT 2.720000 5.305000 2.890000 5.475000 ;
      RECT 2.720000 5.730000 2.890000 5.900000 ;
      RECT 2.965000 0.710000 3.135000 0.880000 ;
      RECT 2.965000 7.740000 3.135000 7.910000 ;
      RECT 3.145000 2.720000 3.315000 2.890000 ;
      RECT 3.145000 5.730000 3.315000 5.900000 ;
      RECT 3.325000 0.710000 3.495000 0.880000 ;
      RECT 3.325000 7.740000 3.495000 7.910000 ;
      RECT 3.505000 2.720000 3.675000 2.890000 ;
      RECT 3.505000 5.730000 3.675000 5.900000 ;
      RECT 3.685000 0.710000 3.855000 0.880000 ;
      RECT 3.685000 7.740000 3.855000 7.910000 ;
      RECT 3.865000 2.720000 4.035000 2.890000 ;
      RECT 3.865000 3.865000 4.755000 4.755000 ;
      RECT 3.865000 5.730000 4.035000 5.900000 ;
      RECT 4.045000 0.710000 4.215000 0.880000 ;
      RECT 4.045000 7.740000 4.215000 7.910000 ;
      RECT 4.225000 2.720000 4.395000 2.890000 ;
      RECT 4.225000 5.730000 4.395000 5.900000 ;
      RECT 4.405000 0.710000 4.575000 0.880000 ;
      RECT 4.405000 7.740000 4.575000 7.910000 ;
      RECT 4.585000 2.720000 4.755000 2.890000 ;
      RECT 4.585000 5.730000 4.755000 5.900000 ;
      RECT 4.765000 0.710000 4.935000 0.880000 ;
      RECT 4.765000 7.740000 4.935000 7.910000 ;
      RECT 4.945000 2.720000 5.115000 2.890000 ;
      RECT 4.945000 5.730000 5.115000 5.900000 ;
      RECT 5.125000 0.710000 5.295000 0.880000 ;
      RECT 5.125000 7.740000 5.295000 7.910000 ;
      RECT 5.305000 2.720000 5.475000 2.890000 ;
      RECT 5.305000 5.730000 5.475000 5.900000 ;
      RECT 5.485000 0.710000 5.655000 0.880000 ;
      RECT 5.485000 7.740000 5.655000 7.910000 ;
      RECT 5.730000 2.720000 5.900000 2.890000 ;
      RECT 5.730000 3.145000 5.900000 3.315000 ;
      RECT 5.730000 3.505000 5.900000 3.675000 ;
      RECT 5.730000 3.865000 5.900000 4.035000 ;
      RECT 5.730000 4.225000 5.900000 4.395000 ;
      RECT 5.730000 4.585000 5.900000 4.755000 ;
      RECT 5.730000 4.945000 5.900000 5.115000 ;
      RECT 5.730000 5.305000 5.900000 5.475000 ;
      RECT 5.730000 5.730000 5.900000 5.900000 ;
      RECT 5.845000 0.710000 6.015000 0.880000 ;
      RECT 5.845000 7.740000 6.015000 7.910000 ;
      RECT 6.205000 0.710000 6.375000 0.880000 ;
      RECT 6.205000 7.740000 6.375000 7.910000 ;
      RECT 6.565000 0.710000 6.735000 0.880000 ;
      RECT 6.565000 7.740000 6.735000 7.910000 ;
      RECT 6.925000 0.710000 7.095000 0.880000 ;
      RECT 6.925000 7.740000 7.095000 7.910000 ;
      RECT 7.285000 0.710000 7.455000 0.880000 ;
      RECT 7.285000 7.740000 7.455000 7.910000 ;
      RECT 7.740000 0.710000 7.910000 0.880000 ;
      RECT 7.740000 1.165000 7.910000 1.335000 ;
      RECT 7.740000 1.525000 7.910000 1.695000 ;
      RECT 7.740000 1.885000 7.910000 2.055000 ;
      RECT 7.740000 2.245000 7.910000 2.415000 ;
      RECT 7.740000 2.605000 7.910000 2.775000 ;
      RECT 7.740000 2.965000 7.910000 3.135000 ;
      RECT 7.740000 3.325000 7.910000 3.495000 ;
      RECT 7.740000 3.685000 7.910000 3.855000 ;
      RECT 7.740000 4.045000 7.910000 4.215000 ;
      RECT 7.740000 4.405000 7.910000 4.575000 ;
      RECT 7.740000 4.765000 7.910000 4.935000 ;
      RECT 7.740000 5.125000 7.910000 5.295000 ;
      RECT 7.740000 5.485000 7.910000 5.655000 ;
      RECT 7.740000 5.845000 7.910000 6.015000 ;
      RECT 7.740000 6.205000 7.910000 6.375000 ;
      RECT 7.740000 6.565000 7.910000 6.735000 ;
      RECT 7.740000 6.925000 7.910000 7.095000 ;
      RECT 7.740000 7.285000 7.910000 7.455000 ;
      RECT 7.740000 7.740000 7.910000 7.910000 ;
    LAYER met1 ;
      RECT 0.650000 0.650000 7.970000 0.940000 ;
      RECT 0.650000 0.940000 0.940000 7.680000 ;
      RECT 0.650000 7.680000 7.970000 7.970000 ;
      RECT 2.660000 2.660000 5.960000 2.950000 ;
      RECT 2.660000 2.950000 2.950000 5.670000 ;
      RECT 2.660000 5.670000 5.960000 5.960000 ;
      RECT 3.805000 3.805000 4.815000 4.815000 ;
      RECT 5.670000 2.950000 5.960000 5.670000 ;
      RECT 7.680000 0.940000 7.970000 7.680000 ;
  END
END sky130_fd_pr__rf_npn_05v5_W1p00L1p00
END LIBRARY
