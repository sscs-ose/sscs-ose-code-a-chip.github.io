# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.880000 BY  6.070000 ;
  PIN BULK
    ANTENNADIFFAREA  2.929000 ;
    PORT
      LAYER li1 ;
        RECT 0.240000 0.610000 0.410000 5.460000 ;
        RECT 4.470000 0.610000 4.640000 5.460000 ;
      LAYER mcon ;
        RECT 0.240000 0.970000 0.410000 1.140000 ;
        RECT 0.240000 1.330000 0.410000 1.500000 ;
        RECT 0.240000 1.690000 0.410000 1.860000 ;
        RECT 0.240000 2.050000 0.410000 2.220000 ;
        RECT 0.240000 2.410000 0.410000 2.580000 ;
        RECT 0.240000 2.770000 0.410000 2.940000 ;
        RECT 0.240000 3.130000 0.410000 3.300000 ;
        RECT 0.240000 3.490000 0.410000 3.660000 ;
        RECT 0.240000 3.850000 0.410000 4.020000 ;
        RECT 0.240000 4.210000 0.410000 4.380000 ;
        RECT 0.240000 4.570000 0.410000 4.740000 ;
        RECT 0.240000 4.930000 0.410000 5.100000 ;
        RECT 0.240000 5.290000 0.410000 5.460000 ;
        RECT 4.470000 0.970000 4.640000 1.140000 ;
        RECT 4.470000 1.330000 4.640000 1.500000 ;
        RECT 4.470000 1.690000 4.640000 1.860000 ;
        RECT 4.470000 2.050000 4.640000 2.220000 ;
        RECT 4.470000 2.410000 4.640000 2.580000 ;
        RECT 4.470000 2.770000 4.640000 2.940000 ;
        RECT 4.470000 3.130000 4.640000 3.300000 ;
        RECT 4.470000 3.490000 4.640000 3.660000 ;
        RECT 4.470000 3.850000 4.640000 4.020000 ;
        RECT 4.470000 4.210000 4.640000 4.380000 ;
        RECT 4.470000 4.570000 4.640000 4.740000 ;
        RECT 4.470000 4.930000 4.640000 5.100000 ;
        RECT 4.470000 5.290000 4.640000 5.460000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.180000 0.550000 0.470000 5.520000 ;
        RECT 4.410000 0.550000 4.700000 5.520000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 3.160000 4.830000 5.520000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  10.099999 ;
    PORT
      LAYER li1 ;
        RECT 0.915000 0.100000 3.965000 0.270000 ;
        RECT 0.915000 5.800000 3.965000 5.970000 ;
      LAYER mcon ;
        RECT 0.915000 0.100000 1.085000 0.270000 ;
        RECT 0.915000 5.800000 1.085000 5.970000 ;
        RECT 1.275000 0.100000 1.445000 0.270000 ;
        RECT 1.275000 5.800000 1.445000 5.970000 ;
        RECT 1.635000 0.100000 1.805000 0.270000 ;
        RECT 1.635000 5.800000 1.805000 5.970000 ;
        RECT 1.995000 0.100000 2.165000 0.270000 ;
        RECT 1.995000 5.800000 2.165000 5.970000 ;
        RECT 2.355000 0.100000 2.525000 0.270000 ;
        RECT 2.355000 5.800000 2.525000 5.970000 ;
        RECT 2.715000 0.100000 2.885000 0.270000 ;
        RECT 2.715000 5.800000 2.885000 5.970000 ;
        RECT 3.075000 0.100000 3.245000 0.270000 ;
        RECT 3.075000 5.800000 3.245000 5.970000 ;
        RECT 3.435000 0.100000 3.605000 0.270000 ;
        RECT 3.435000 5.800000 3.605000 5.970000 ;
        RECT 3.795000 0.100000 3.965000 0.270000 ;
        RECT 3.795000 5.800000 3.965000 5.970000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.855000 0.000000 4.025000 0.330000 ;
        RECT 0.855000 5.740000 4.025000 6.070000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.550000 4.830000 2.910000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.795000 0.490000 0.965000 5.580000 ;
      RECT 1.575000 0.490000 1.745000 5.580000 ;
      RECT 2.355000 0.490000 2.525000 5.580000 ;
      RECT 3.135000 0.490000 3.305000 5.580000 ;
      RECT 3.915000 0.490000 4.085000 5.580000 ;
    LAYER mcon ;
      RECT 0.795000 0.610000 0.965000 0.780000 ;
      RECT 0.795000 0.970000 0.965000 1.140000 ;
      RECT 0.795000 1.330000 0.965000 1.500000 ;
      RECT 0.795000 1.690000 0.965000 1.860000 ;
      RECT 0.795000 2.050000 0.965000 2.220000 ;
      RECT 0.795000 2.410000 0.965000 2.580000 ;
      RECT 0.795000 2.770000 0.965000 2.940000 ;
      RECT 0.795000 3.130000 0.965000 3.300000 ;
      RECT 0.795000 3.490000 0.965000 3.660000 ;
      RECT 0.795000 3.850000 0.965000 4.020000 ;
      RECT 0.795000 4.210000 0.965000 4.380000 ;
      RECT 0.795000 4.570000 0.965000 4.740000 ;
      RECT 0.795000 4.930000 0.965000 5.100000 ;
      RECT 0.795000 5.290000 0.965000 5.460000 ;
      RECT 1.575000 0.610000 1.745000 0.780000 ;
      RECT 1.575000 0.970000 1.745000 1.140000 ;
      RECT 1.575000 1.330000 1.745000 1.500000 ;
      RECT 1.575000 1.690000 1.745000 1.860000 ;
      RECT 1.575000 2.050000 1.745000 2.220000 ;
      RECT 1.575000 2.410000 1.745000 2.580000 ;
      RECT 1.575000 2.770000 1.745000 2.940000 ;
      RECT 1.575000 3.130000 1.745000 3.300000 ;
      RECT 1.575000 3.490000 1.745000 3.660000 ;
      RECT 1.575000 3.850000 1.745000 4.020000 ;
      RECT 1.575000 4.210000 1.745000 4.380000 ;
      RECT 1.575000 4.570000 1.745000 4.740000 ;
      RECT 1.575000 4.930000 1.745000 5.100000 ;
      RECT 1.575000 5.290000 1.745000 5.460000 ;
      RECT 2.355000 0.610000 2.525000 0.780000 ;
      RECT 2.355000 0.970000 2.525000 1.140000 ;
      RECT 2.355000 1.330000 2.525000 1.500000 ;
      RECT 2.355000 1.690000 2.525000 1.860000 ;
      RECT 2.355000 2.050000 2.525000 2.220000 ;
      RECT 2.355000 2.410000 2.525000 2.580000 ;
      RECT 2.355000 2.770000 2.525000 2.940000 ;
      RECT 2.355000 3.130000 2.525000 3.300000 ;
      RECT 2.355000 3.490000 2.525000 3.660000 ;
      RECT 2.355000 3.850000 2.525000 4.020000 ;
      RECT 2.355000 4.210000 2.525000 4.380000 ;
      RECT 2.355000 4.570000 2.525000 4.740000 ;
      RECT 2.355000 4.930000 2.525000 5.100000 ;
      RECT 2.355000 5.290000 2.525000 5.460000 ;
      RECT 3.135000 0.610000 3.305000 0.780000 ;
      RECT 3.135000 0.970000 3.305000 1.140000 ;
      RECT 3.135000 1.330000 3.305000 1.500000 ;
      RECT 3.135000 1.690000 3.305000 1.860000 ;
      RECT 3.135000 2.050000 3.305000 2.220000 ;
      RECT 3.135000 2.410000 3.305000 2.580000 ;
      RECT 3.135000 2.770000 3.305000 2.940000 ;
      RECT 3.135000 3.130000 3.305000 3.300000 ;
      RECT 3.135000 3.490000 3.305000 3.660000 ;
      RECT 3.135000 3.850000 3.305000 4.020000 ;
      RECT 3.135000 4.210000 3.305000 4.380000 ;
      RECT 3.135000 4.570000 3.305000 4.740000 ;
      RECT 3.135000 4.930000 3.305000 5.100000 ;
      RECT 3.135000 5.290000 3.305000 5.460000 ;
      RECT 3.915000 0.610000 4.085000 0.780000 ;
      RECT 3.915000 0.970000 4.085000 1.140000 ;
      RECT 3.915000 1.330000 4.085000 1.500000 ;
      RECT 3.915000 1.690000 4.085000 1.860000 ;
      RECT 3.915000 2.050000 4.085000 2.220000 ;
      RECT 3.915000 2.410000 4.085000 2.580000 ;
      RECT 3.915000 2.770000 4.085000 2.940000 ;
      RECT 3.915000 3.130000 4.085000 3.300000 ;
      RECT 3.915000 3.490000 4.085000 3.660000 ;
      RECT 3.915000 3.850000 4.085000 4.020000 ;
      RECT 3.915000 4.210000 4.085000 4.380000 ;
      RECT 3.915000 4.570000 4.085000 4.740000 ;
      RECT 3.915000 4.930000 4.085000 5.100000 ;
      RECT 3.915000 5.290000 4.085000 5.460000 ;
    LAYER met1 ;
      RECT 0.750000 0.550000 1.010000 5.520000 ;
      RECT 1.530000 0.550000 1.790000 5.520000 ;
      RECT 2.310000 0.550000 2.570000 5.520000 ;
      RECT 3.090000 0.550000 3.350000 5.520000 ;
      RECT 3.870000 0.550000 4.130000 5.520000 ;
    LAYER via ;
      RECT 0.750000 0.580000 1.010000 0.840000 ;
      RECT 0.750000 0.900000 1.010000 1.160000 ;
      RECT 0.750000 1.220000 1.010000 1.480000 ;
      RECT 0.750000 1.540000 1.010000 1.800000 ;
      RECT 0.750000 1.860000 1.010000 2.120000 ;
      RECT 0.750000 2.180000 1.010000 2.440000 ;
      RECT 0.750000 2.500000 1.010000 2.760000 ;
      RECT 1.530000 3.310000 1.790000 3.570000 ;
      RECT 1.530000 3.630000 1.790000 3.890000 ;
      RECT 1.530000 3.950000 1.790000 4.210000 ;
      RECT 1.530000 4.270000 1.790000 4.530000 ;
      RECT 1.530000 4.590000 1.790000 4.850000 ;
      RECT 1.530000 4.910000 1.790000 5.170000 ;
      RECT 1.530000 5.230000 1.790000 5.490000 ;
      RECT 2.310000 0.580000 2.570000 0.840000 ;
      RECT 2.310000 0.900000 2.570000 1.160000 ;
      RECT 2.310000 1.220000 2.570000 1.480000 ;
      RECT 2.310000 1.540000 2.570000 1.800000 ;
      RECT 2.310000 1.860000 2.570000 2.120000 ;
      RECT 2.310000 2.180000 2.570000 2.440000 ;
      RECT 2.310000 2.500000 2.570000 2.760000 ;
      RECT 3.090000 3.310000 3.350000 3.570000 ;
      RECT 3.090000 3.630000 3.350000 3.890000 ;
      RECT 3.090000 3.950000 3.350000 4.210000 ;
      RECT 3.090000 4.270000 3.350000 4.530000 ;
      RECT 3.090000 4.590000 3.350000 4.850000 ;
      RECT 3.090000 4.910000 3.350000 5.170000 ;
      RECT 3.090000 5.230000 3.350000 5.490000 ;
      RECT 3.870000 0.580000 4.130000 0.840000 ;
      RECT 3.870000 0.900000 4.130000 1.160000 ;
      RECT 3.870000 1.220000 4.130000 1.480000 ;
      RECT 3.870000 1.540000 4.130000 1.800000 ;
      RECT 3.870000 1.860000 4.130000 2.120000 ;
      RECT 3.870000 2.180000 4.130000 2.440000 ;
      RECT 3.870000 2.500000 4.130000 2.760000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50
END LIBRARY
