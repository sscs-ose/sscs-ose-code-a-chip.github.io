MACRO NMOS_S_33976710_X10_Y5
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_33976710_X10_Y5 0 0 ;
  SIZE 10320 BY 31080 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4590 260 4870 24100 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5020 4460 5300 28300 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5450 680 5730 30400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 30745 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 30745 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 30745 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 30745 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 30745 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 21505 ;
    LAYER M1 ;
      RECT 5465 21755 5715 22765 ;
    LAYER M1 ;
      RECT 5465 23855 5715 27385 ;
    LAYER M1 ;
      RECT 5465 27635 5715 28645 ;
    LAYER M1 ;
      RECT 5465 29735 5715 30745 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 5895 23855 6145 27385 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 21505 ;
    LAYER M1 ;
      RECT 6325 21755 6575 22765 ;
    LAYER M1 ;
      RECT 6325 23855 6575 27385 ;
    LAYER M1 ;
      RECT 6325 27635 6575 28645 ;
    LAYER M1 ;
      RECT 6325 29735 6575 30745 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 6755 17975 7005 21505 ;
    LAYER M1 ;
      RECT 6755 23855 7005 27385 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 21505 ;
    LAYER M1 ;
      RECT 7185 21755 7435 22765 ;
    LAYER M1 ;
      RECT 7185 23855 7435 27385 ;
    LAYER M1 ;
      RECT 7185 27635 7435 28645 ;
    LAYER M1 ;
      RECT 7185 29735 7435 30745 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 7615 17975 7865 21505 ;
    LAYER M1 ;
      RECT 7615 23855 7865 27385 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 15625 ;
    LAYER M1 ;
      RECT 8045 15875 8295 16885 ;
    LAYER M1 ;
      RECT 8045 17975 8295 21505 ;
    LAYER M1 ;
      RECT 8045 21755 8295 22765 ;
    LAYER M1 ;
      RECT 8045 23855 8295 27385 ;
    LAYER M1 ;
      RECT 8045 27635 8295 28645 ;
    LAYER M1 ;
      RECT 8045 29735 8295 30745 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8475 12095 8725 15625 ;
    LAYER M1 ;
      RECT 8475 17975 8725 21505 ;
    LAYER M1 ;
      RECT 8475 23855 8725 27385 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 15625 ;
    LAYER M1 ;
      RECT 8905 15875 9155 16885 ;
    LAYER M1 ;
      RECT 8905 17975 9155 21505 ;
    LAYER M1 ;
      RECT 8905 21755 9155 22765 ;
    LAYER M1 ;
      RECT 8905 23855 9155 27385 ;
    LAYER M1 ;
      RECT 8905 27635 9155 28645 ;
    LAYER M1 ;
      RECT 8905 29735 9155 30745 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9335 12095 9585 15625 ;
    LAYER M1 ;
      RECT 9335 17975 9585 21505 ;
    LAYER M1 ;
      RECT 9335 23855 9585 27385 ;
    LAYER M2 ;
      RECT 1120 280 9200 560 ;
    LAYER M2 ;
      RECT 1120 4480 9200 4760 ;
    LAYER M2 ;
      RECT 690 700 9630 980 ;
    LAYER M2 ;
      RECT 1120 6160 9200 6440 ;
    LAYER M2 ;
      RECT 1120 10360 9200 10640 ;
    LAYER M2 ;
      RECT 690 6580 9630 6860 ;
    LAYER M2 ;
      RECT 1120 12040 9200 12320 ;
    LAYER M2 ;
      RECT 1120 16240 9200 16520 ;
    LAYER M2 ;
      RECT 690 12460 9630 12740 ;
    LAYER M2 ;
      RECT 1120 17920 9200 18200 ;
    LAYER M2 ;
      RECT 1120 22120 9200 22400 ;
    LAYER M2 ;
      RECT 690 18340 9630 18620 ;
    LAYER M2 ;
      RECT 1120 23800 9200 24080 ;
    LAYER M2 ;
      RECT 1120 28000 9200 28280 ;
    LAYER M2 ;
      RECT 1120 30100 9200 30380 ;
    LAYER M2 ;
      RECT 690 24220 9630 24500 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 30155 1375 30325 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 30155 2235 30325 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 30155 3095 30325 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 30155 3955 30325 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 30155 4815 30325 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 17975 5675 18145 ;
    LAYER V1 ;
      RECT 5505 22175 5675 22345 ;
    LAYER V1 ;
      RECT 5505 23855 5675 24025 ;
    LAYER V1 ;
      RECT 5505 28055 5675 28225 ;
    LAYER V1 ;
      RECT 5505 30155 5675 30325 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 17975 6535 18145 ;
    LAYER V1 ;
      RECT 6365 22175 6535 22345 ;
    LAYER V1 ;
      RECT 6365 23855 6535 24025 ;
    LAYER V1 ;
      RECT 6365 28055 6535 28225 ;
    LAYER V1 ;
      RECT 6365 30155 6535 30325 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 17975 7395 18145 ;
    LAYER V1 ;
      RECT 7225 22175 7395 22345 ;
    LAYER V1 ;
      RECT 7225 23855 7395 24025 ;
    LAYER V1 ;
      RECT 7225 28055 7395 28225 ;
    LAYER V1 ;
      RECT 7225 30155 7395 30325 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12095 8255 12265 ;
    LAYER V1 ;
      RECT 8085 16295 8255 16465 ;
    LAYER V1 ;
      RECT 8085 17975 8255 18145 ;
    LAYER V1 ;
      RECT 8085 22175 8255 22345 ;
    LAYER V1 ;
      RECT 8085 23855 8255 24025 ;
    LAYER V1 ;
      RECT 8085 28055 8255 28225 ;
    LAYER V1 ;
      RECT 8085 30155 8255 30325 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12095 9115 12265 ;
    LAYER V1 ;
      RECT 8945 16295 9115 16465 ;
    LAYER V1 ;
      RECT 8945 17975 9115 18145 ;
    LAYER V1 ;
      RECT 8945 22175 9115 22345 ;
    LAYER V1 ;
      RECT 8945 23855 9115 24025 ;
    LAYER V1 ;
      RECT 8945 28055 9115 28225 ;
    LAYER V1 ;
      RECT 8945 30155 9115 30325 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 5935 18395 6105 18565 ;
    LAYER V1 ;
      RECT 5935 24275 6105 24445 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 6795 18395 6965 18565 ;
    LAYER V1 ;
      RECT 6795 24275 6965 24445 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V1 ;
      RECT 7655 18395 7825 18565 ;
    LAYER V1 ;
      RECT 7655 24275 7825 24445 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 8515 12515 8685 12685 ;
    LAYER V1 ;
      RECT 8515 18395 8685 18565 ;
    LAYER V1 ;
      RECT 8515 24275 8685 24445 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 9375 6635 9545 6805 ;
    LAYER V1 ;
      RECT 9375 12515 9545 12685 ;
    LAYER V1 ;
      RECT 9375 18395 9545 18565 ;
    LAYER V1 ;
      RECT 9375 24275 9545 24445 ;
    LAYER V2 ;
      RECT 4655 345 4805 495 ;
    LAYER V2 ;
      RECT 4655 6225 4805 6375 ;
    LAYER V2 ;
      RECT 4655 12105 4805 12255 ;
    LAYER V2 ;
      RECT 4655 17985 4805 18135 ;
    LAYER V2 ;
      RECT 4655 23865 4805 24015 ;
    LAYER V2 ;
      RECT 5085 4545 5235 4695 ;
    LAYER V2 ;
      RECT 5085 10425 5235 10575 ;
    LAYER V2 ;
      RECT 5085 16305 5235 16455 ;
    LAYER V2 ;
      RECT 5085 22185 5235 22335 ;
    LAYER V2 ;
      RECT 5085 28065 5235 28215 ;
    LAYER V2 ;
      RECT 5515 765 5665 915 ;
    LAYER V2 ;
      RECT 5515 6645 5665 6795 ;
    LAYER V2 ;
      RECT 5515 12525 5665 12675 ;
    LAYER V2 ;
      RECT 5515 18405 5665 18555 ;
    LAYER V2 ;
      RECT 5515 24285 5665 24435 ;
    LAYER V2 ;
      RECT 5515 30165 5665 30315 ;
  END
END NMOS_S_33976710_X10_Y5
