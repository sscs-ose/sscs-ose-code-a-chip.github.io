* Transient simulation

.lib "../skywater_pdk/sky130_fd_pr/models/sky130.lib.spice" tt

* Pulsegen ckt
.include pulsegen.cir

v1 vdd gnd dc 3.3
v2 vss gnd dc 0
v3 in gnd pulse(0 3.3 0 30n 15n 1u 2u)

X1 vdd vss in outp outm pulsegen

C1 outp gnd 50ff 
C2 outm gnd 50ff

*Simulation Command
.tran 0.05u 4u

* ngspice control statements
.control

run
* print v(in) v(outp) v(outm) > plot_data_v.txt
* print alli > plot_data_i.txt
plot v(in) v(outp) v(outm)

*For Transient Analysis
*hardcopy file.svg v(inAC1) v(inAC2) v(out2) ; diff amplifier
*hardcopy file plotargs v(out2) v(out3) v(out4) ; high-pass filter and buffer
*hardcopy file plotargs v(inOff) v(out4) v(out5) ; non-inv amplifier
*hardcopy file plotargs v(out5) v(inOff) v(out6) ; comparator

.endc

.end
