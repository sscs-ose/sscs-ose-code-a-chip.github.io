# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_test_coil3
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_test_coil3 ;
  ORIGIN  182.5400  182.5400 ;
  SIZE  370.0800 BY  365.0800 ;
  OBS
    LAYER met2 ;
      POLYGON -10.115000  125.010000   4.895000  125.010000   4.895000  110.000000 ;
      POLYGON -10.115000  155.030000   4.895000  155.030000   4.895000  140.020000 ;
      POLYGON  -4.935000 -170.040000   7.565000 -170.040000  -4.935000 -182.540000 ;
      POLYGON  -4.935000 -140.020000   7.565000 -140.020000  -4.935000 -152.520000 ;
      POLYGON  -4.935000  137.510000   7.565000  125.010000  -4.935000  125.010000 ;
      POLYGON  -4.935000  167.530000   7.565000  155.030000  -4.935000  155.030000 ;
      POLYGON   4.895000 -155.030000   4.895000 -170.040000 -10.115000 -170.040000 ;
      POLYGON   4.895000 -125.010000   4.895000 -140.020000 -10.115000 -140.020000 ;
      POLYGON   7.565000 -167.530000  10.075000 -167.530000   7.565000 -170.040000 ;
      POLYGON   7.565000 -137.510000  10.075000 -137.510000   7.565000 -140.020000 ;
      POLYGON   7.565000  125.010000  10.075000  122.500000   7.565000  122.500000 ;
      POLYGON   7.565000  155.030000  10.075000  152.520000   7.565000  152.520000 ;
      RECT -37.720000 -182.540000  -4.935000 -170.040000 ;
      RECT -37.720000 -152.520000  -4.935000 -140.020000 ;
      RECT -37.160000  125.010000  -4.935000  137.510000 ;
      RECT -37.160000  155.030000  -4.935000  167.530000 ;
      RECT   4.895000 -170.040000   7.565000 -167.530000 ;
      RECT   4.895000 -167.530000  38.375000 -155.030000 ;
      RECT   4.895000 -140.020000   7.565000 -137.510000 ;
      RECT   4.895000 -137.510000  38.375000 -125.010000 ;
      RECT   4.895000  110.000000  38.935000  122.500000 ;
      RECT   4.895000  122.500000   7.565000  125.010000 ;
      RECT   4.895000  140.020000  38.935000  152.520000 ;
      RECT   4.895000  152.520000   7.565000  155.030000 ;
      RECT  97.040000   -6.250000 187.540000    6.250000 ;
    LAYER met3 ;
      POLYGON -182.540000  -75.620000 -171.075000  -75.620000 -171.075000  -87.085000 ;
      POLYGON -171.075000  -87.085000 -153.395000  -87.085000 -153.395000 -104.765000 ;
      POLYGON -170.040000  -70.440000 -167.530000  -72.950000 -170.040000  -72.950000 ;
      POLYGON -170.040000   72.950000 -167.530000   72.950000 -170.040000   70.440000 ;
      POLYGON -167.530000  -72.950000 -164.020000  -76.460000 -167.530000  -76.460000 ;
      POLYGON -167.530000  -69.405000 -166.495000  -69.405000 -166.495000  -70.440000 ;
      POLYGON -167.530000   75.620000 -164.860000   75.620000 -167.530000   72.950000 ;
      POLYGON -166.495000  -70.440000 -163.985000  -70.440000 -163.985000  -72.950000 ;
      POLYGON -166.495000   70.440000 -166.495000   69.405000 -167.530000   69.405000 ;
      POLYGON -164.860000   79.130000 -161.350000   79.130000 -164.860000   75.620000 ;
      POLYGON -164.860000   93.300000 -164.860000   75.620000 -182.540000   75.620000 ;
      POLYGON -164.020000  -76.460000 -160.475000  -80.005000 -164.020000  -80.005000 ;
      POLYGON -163.985000  -72.950000 -160.475000  -72.950000 -160.475000  -76.460000 ;
      POLYGON -163.985000   72.950000 -163.985000   70.440000 -166.495000   70.440000 ;
      POLYGON -161.350000   82.675000 -157.805000   82.675000 -161.350000   79.130000 ;
      POLYGON -161.315000   75.620000 -161.315000   72.950000 -163.985000   72.950000 ;
      POLYGON -160.475000  -80.005000 -156.940000  -83.540000 -160.475000  -83.540000 ;
      POLYGON -160.475000  -76.460000 -156.930000  -76.460000 -156.930000  -80.005000 ;
      POLYGON -157.805000   79.130000 -157.805000   75.620000 -161.315000   75.620000 ;
      POLYGON -157.805000   86.220000 -154.260000   86.220000 -157.805000   82.675000 ;
      POLYGON -156.940000  -83.540000 -153.395000  -87.085000 -156.940000  -87.085000 ;
      POLYGON -156.930000  -80.005000 -153.395000  -80.005000 -153.395000  -83.540000 ;
      POLYGON -155.030000  -64.225000 -152.520000  -66.735000 -155.030000  -66.735000 ;
      POLYGON -155.030000   67.670000 -151.585000   67.670000 -155.030000   64.225000 ;
      POLYGON -154.260000   82.675000 -154.260000   79.130000 -157.805000   79.130000 ;
      POLYGON -154.260000   89.755000 -150.725000   89.755000 -154.260000   86.220000 ;
      POLYGON -153.395000 -104.765000 -135.715000 -104.765000 -135.715000 -122.445000 ;
      POLYGON -153.395000  -87.085000 -149.850000  -90.630000 -153.395000  -90.630000 ;
      POLYGON -153.395000  -83.540000 -149.850000  -83.540000 -149.850000  -87.085000 ;
      POLYGON -152.520000  -66.735000 -149.850000  -69.405000 -152.520000  -69.405000 ;
      POLYGON -152.520000  -63.185000 -151.480000  -63.185000 -151.480000  -64.225000 ;
      POLYGON -151.585000   64.120000 -151.585000   63.185000 -152.520000   63.185000 ;
      POLYGON -151.585000   69.405000 -149.850000   69.405000 -151.585000   67.670000 ;
      POLYGON -151.480000  -64.225000 -148.970000  -64.225000 -148.970000  -66.735000 ;
      POLYGON -151.480000   64.225000 -151.480000   64.120000 -151.585000   64.120000 ;
      POLYGON -150.725000   93.300000 -147.180000   93.300000 -150.725000   89.755000 ;
      POLYGON -150.715000   86.220000 -150.715000   82.675000 -154.260000   82.675000 ;
      POLYGON -149.850000  -90.630000 -146.340000  -94.140000 -149.850000  -94.140000 ;
      POLYGON -149.850000  -87.085000 -146.305000  -87.085000 -146.305000  -90.630000 ;
      POLYGON -149.850000  -69.405000 -147.185000  -72.070000 -149.850000  -72.070000 ;
      POLYGON -149.850000   72.070000 -147.185000   72.070000 -149.850000   69.405000 ;
      POLYGON -148.970000  -66.735000 -146.300000  -66.735000 -146.300000  -69.405000 ;
      POLYGON -148.035000   67.670000 -148.035000   64.225000 -151.480000   64.225000 ;
      POLYGON -147.185000  -72.070000 -143.635000  -75.620000 -147.185000  -75.620000 ;
      POLYGON -147.185000   75.620000 -143.635000   75.620000 -147.185000   72.070000 ;
      POLYGON -147.180000   89.755000 -147.180000   86.220000 -150.715000   86.220000 ;
      POLYGON -147.180000   96.810000 -143.670000   96.810000 -147.180000   93.300000 ;
      POLYGON -147.180000  110.980000 -147.180000   93.300000 -164.860000   93.300000 ;
      POLYGON -146.340000  -94.140000 -142.795000  -97.685000 -146.340000  -97.685000 ;
      POLYGON -146.305000  -90.630000 -142.795000  -90.630000 -142.795000  -94.140000 ;
      POLYGON -146.300000  -69.405000 -143.635000  -69.405000 -143.635000  -72.070000 ;
      POLYGON -146.300000   69.405000 -146.300000   67.670000 -148.035000   67.670000 ;
      POLYGON -145.265000   70.440000 -145.265000   69.405000 -146.300000   69.405000 ;
      POLYGON -143.670000  100.355000 -140.125000  100.355000 -143.670000   96.810000 ;
      POLYGON -143.635000  -75.620000 -140.125000  -79.130000 -143.635000  -79.130000 ;
      POLYGON -143.635000  -72.070000 -140.085000  -72.070000 -140.085000  -75.620000 ;
      POLYGON -143.635000   72.070000 -143.635000   70.440000 -145.265000   70.440000 ;
      POLYGON -143.635000   79.130000 -140.125000   79.130000 -143.635000   75.620000 ;
      POLYGON -143.635000   93.300000 -143.635000   89.755000 -147.180000   89.755000 ;
      POLYGON -142.795000  -97.685000 -139.260000 -101.220000 -142.795000 -101.220000 ;
      POLYGON -142.795000  -94.140000 -139.250000  -94.140000 -139.250000  -97.685000 ;
      POLYGON -140.125000  -79.130000 -138.390000  -80.865000 -140.125000  -80.865000 ;
      POLYGON -140.125000   81.800000 -137.455000   81.800000 -140.125000   79.130000 ;
      POLYGON -140.125000   96.810000 -140.125000   93.300000 -143.635000   93.300000 ;
      POLYGON -140.125000  103.900000 -136.580000  103.900000 -140.125000  100.355000 ;
      POLYGON -140.085000  -75.620000 -136.575000  -75.620000 -136.575000  -79.130000 ;
      POLYGON -140.085000   75.620000 -140.085000   72.070000 -143.635000   72.070000 ;
      POLYGON -140.020000  -58.005000 -137.510000  -60.515000 -140.020000  -60.515000 ;
      POLYGON -140.020000   60.515000 -137.510000   60.515000 -140.020000   58.005000 ;
      POLYGON -139.735000  118.425000 -139.735000  110.980000 -147.180000  110.980000 ;
      POLYGON -139.260000 -101.220000 -135.715000 -104.765000 -139.260000 -104.765000 ;
      POLYGON -139.250000  -97.685000 -135.715000  -97.685000 -135.715000 -101.220000 ;
      POLYGON -138.390000  -80.865000 -134.840000  -84.415000 -138.390000  -84.415000 ;
      POLYGON -137.510000  -60.515000 -134.840000  -63.185000 -137.510000  -63.185000 ;
      POLYGON -137.510000  -56.970000 -136.475000  -56.970000 -136.475000  -58.005000 ;
      POLYGON -137.510000   63.185000 -134.840000   63.185000 -137.510000   60.515000 ;
      POLYGON -137.455000   85.350000 -133.905000   85.350000 -137.455000   81.800000 ;
      POLYGON -136.580000  100.355000 -136.580000   96.810000 -140.125000   96.810000 ;
      POLYGON -136.580000  107.435000 -133.045000  107.435000 -136.580000  103.900000 ;
      POLYGON -136.575000  -79.130000 -134.840000  -79.130000 -134.840000  -80.865000 ;
      POLYGON -136.575000   79.130000 -136.575000   75.620000 -140.085000   75.620000 ;
      POLYGON -136.475000  -58.005000 -133.965000  -58.005000 -133.965000  -60.515000 ;
      POLYGON -136.475000   58.005000 -136.475000   56.970000 -137.510000   56.970000 ;
      POLYGON -135.715000 -122.445000 -118.035000 -122.445000 -118.035000 -140.125000 ;
      POLYGON -135.715000 -104.765000 -132.170000 -108.310000 -135.715000 -108.310000 ;
      POLYGON -135.715000 -101.220000 -132.170000 -101.220000 -132.170000 -104.765000 ;
      POLYGON -134.840000  -84.415000 -132.170000  -87.085000 -134.840000  -87.085000 ;
      POLYGON -134.840000  -80.865000 -131.290000  -80.865000 -131.290000  -84.415000 ;
      POLYGON -134.840000  -63.185000 -132.165000  -65.860000 -134.840000  -65.860000 ;
      POLYGON -134.840000   64.120000 -133.905000   64.120000 -134.840000   63.185000 ;
      POLYGON -133.965000  -60.515000 -131.295000  -60.515000 -131.295000  -63.185000 ;
      POLYGON -133.965000   60.515000 -133.965000   58.005000 -136.475000   58.005000 ;
      POLYGON -133.905000   66.790000 -131.235000   66.790000 -133.905000   64.120000 ;
      POLYGON -133.905000   81.800000 -133.905000   79.130000 -136.575000   79.130000 ;
      POLYGON -133.905000   87.085000 -132.170000   87.085000 -133.905000   85.350000 ;
      POLYGON -133.045000  110.980000 -129.500000  110.980000 -133.045000  107.435000 ;
      POLYGON -133.035000  103.900000 -133.035000  100.355000 -136.580000  100.355000 ;
      POLYGON -132.170000 -108.310000 -128.660000 -111.820000 -132.170000 -111.820000 ;
      POLYGON -132.170000 -104.765000 -128.625000 -104.765000 -128.625000 -108.310000 ;
      POLYGON -132.170000  -87.085000 -129.505000  -89.750000 -132.170000  -89.750000 ;
      POLYGON -132.170000   89.750000 -129.505000   89.750000 -132.170000   87.085000 ;
      POLYGON -132.165000  -65.860000 -128.620000  -69.405000 -132.165000  -69.405000 ;
      POLYGON -131.545000  126.615000 -131.545000  118.425000 -139.735000  118.425000 ;
      POLYGON -131.295000  -63.185000 -128.620000  -63.185000 -128.620000  -65.860000 ;
      POLYGON -131.295000   63.185000 -131.295000   60.515000 -133.965000   60.515000 ;
      POLYGON -131.290000  -84.415000 -128.620000  -84.415000 -128.620000  -87.085000 ;
      POLYGON -131.235000   69.405000 -128.620000   69.405000 -131.235000   66.790000 ;
      POLYGON -130.360000   64.120000 -130.360000   63.185000 -131.295000   63.185000 ;
      POLYGON -130.355000   85.350000 -130.355000   81.800000 -133.905000   81.800000 ;
      POLYGON -129.505000  -89.750000 -125.955000  -93.300000 -129.505000  -93.300000 ;
      POLYGON -129.505000   93.300000 -125.955000   93.300000 -129.505000   89.750000 ;
      POLYGON -129.500000  107.435000 -129.500000  103.900000 -133.035000  103.900000 ;
      POLYGON -129.500000  114.490000 -125.990000  114.490000 -129.500000  110.980000 ;
      POLYGON -128.660000 -111.820000 -125.115000 -115.365000 -128.660000 -115.365000 ;
      POLYGON -128.625000 -108.310000 -125.115000 -108.310000 -125.115000 -111.820000 ;
      POLYGON -128.620000  -87.085000 -125.955000  -87.085000 -125.955000  -89.750000 ;
      POLYGON -128.620000  -69.405000 -126.920000  -71.105000 -128.620000  -71.105000 ;
      POLYGON -128.620000  -65.860000 -125.075000  -65.860000 -125.075000  -69.405000 ;
      POLYGON -128.620000   72.075000 -125.950000   72.075000 -128.620000   69.405000 ;
      POLYGON -128.620000   87.085000 -128.620000   85.350000 -130.355000   85.350000 ;
      POLYGON -127.690000   66.790000 -127.690000   64.120000 -130.360000   64.120000 ;
      POLYGON -126.920000  -71.105000 -123.375000  -74.650000 -126.920000  -74.650000 ;
      POLYGON -125.990000  118.035000 -122.445000  118.035000 -125.990000  114.490000 ;
      POLYGON -125.955000  -93.300000 -122.445000  -96.810000 -125.955000  -96.810000 ;
      POLYGON -125.955000  -89.750000 -122.405000  -89.750000 -122.405000  -93.300000 ;
      POLYGON -125.955000   89.750000 -125.955000   87.085000 -128.620000   87.085000 ;
      POLYGON -125.955000   96.810000 -122.445000   96.810000 -125.955000   93.300000 ;
      POLYGON -125.955000  110.980000 -125.955000  107.435000 -129.500000  107.435000 ;
      POLYGON -125.950000   75.620000 -122.405000   75.620000 -125.950000   72.075000 ;
      POLYGON -125.115000 -115.365000 -121.580000 -118.900000 -125.115000 -118.900000 ;
      POLYGON -125.115000 -111.820000 -121.570000 -111.820000 -121.570000 -115.365000 ;
      POLYGON -125.075000  -69.405000 -123.375000  -69.405000 -123.375000  -71.105000 ;
      POLYGON -125.075000   69.405000 -125.075000   66.790000 -127.690000   66.790000 ;
      POLYGON -125.010000  -51.790000 -122.500000  -54.300000 -125.010000  -54.300000 ;
      POLYGON -125.010000   55.330000 -121.470000   55.330000 -125.010000   51.790000 ;
      POLYGON -124.145000   70.335000 -124.145000   69.405000 -125.075000   69.405000 ;
      POLYGON -123.375000  -74.650000 -119.830000  -78.195000 -123.375000  -78.195000 ;
      POLYGON -123.375000  -71.105000 -119.830000  -71.105000 -119.830000  -74.650000 ;
      POLYGON -122.500000  -54.300000 -119.830000  -56.970000 -122.500000  -56.970000 ;
      POLYGON -122.500000  -50.750000 -121.460000  -50.750000 -121.460000  -51.790000 ;
      POLYGON -122.445000  -96.810000 -120.710000  -98.545000 -122.445000  -98.545000 ;
      POLYGON -122.445000   99.480000 -119.775000   99.480000 -122.445000   96.810000 ;
      POLYGON -122.445000  114.490000 -122.445000  110.980000 -125.955000  110.980000 ;
      POLYGON -122.445000  121.580000 -118.900000  121.580000 -122.445000  118.035000 ;
      POLYGON -122.405000  -93.300000 -118.895000  -93.300000 -118.895000  -96.810000 ;
      POLYGON -122.405000   72.075000 -122.405000   70.335000 -124.145000   70.335000 ;
      POLYGON -122.405000   79.130000 -118.895000   79.130000 -122.405000   75.620000 ;
      POLYGON -122.405000   93.300000 -122.405000   89.750000 -125.955000   89.750000 ;
      POLYGON -122.255000  135.905000 -122.255000  126.615000 -131.545000  126.615000 ;
      POLYGON -121.580000 -118.900000 -118.035000 -122.445000 -121.580000 -122.445000 ;
      POLYGON -121.570000 -115.365000 -118.035000 -115.365000 -118.035000 -118.900000 ;
      POLYGON -121.470000   51.780000 -121.470000   50.750000 -122.500000   50.750000 ;
      POLYGON -121.470000   56.970000 -119.830000   56.970000 -121.470000   55.330000 ;
      POLYGON -121.460000  -51.790000 -118.950000  -51.790000 -118.950000  -54.300000 ;
      POLYGON -121.460000   51.790000 -121.460000   51.780000 -121.470000   51.780000 ;
      POLYGON -120.710000  -98.545000 -117.160000 -102.095000 -120.710000 -102.095000 ;
      POLYGON -119.830000  -78.195000 -117.160000  -80.865000 -119.830000  -80.865000 ;
      POLYGON -119.830000  -74.650000 -116.285000  -74.650000 -116.285000  -78.195000 ;
      POLYGON -119.830000  -56.970000 -117.165000  -59.635000 -119.830000  -59.635000 ;
      POLYGON -119.830000   59.635000 -117.165000   59.635000 -119.830000   56.970000 ;
      POLYGON -119.830000   74.650000 -119.830000   72.075000 -122.405000   72.075000 ;
      POLYGON -119.775000  103.030000 -116.225000  103.030000 -119.775000   99.480000 ;
      POLYGON -118.950000  -54.300000 -116.280000  -54.300000 -116.280000  -56.970000 ;
      POLYGON -118.900000  118.035000 -118.900000  114.490000 -122.445000  114.490000 ;
      POLYGON -118.900000  125.115000 -115.365000  125.115000 -118.900000  121.580000 ;
      POLYGON -118.895000  -96.810000 -117.160000  -96.810000 -117.160000  -98.545000 ;
      POLYGON -118.895000   81.800000 -116.225000   81.800000 -118.895000   79.130000 ;
      POLYGON -118.895000   96.810000 -118.895000   93.300000 -122.405000   93.300000 ;
      POLYGON -118.860000   75.620000 -118.860000   74.650000 -119.830000   74.650000 ;
      POLYGON -118.035000 -140.125000 -100.355000 -140.125000 -100.355000 -157.805000 ;
      POLYGON -118.035000 -122.445000 -114.490000 -125.990000 -118.035000 -125.990000 ;
      POLYGON -118.035000 -118.900000 -114.490000 -118.900000 -114.490000 -122.445000 ;
      POLYGON -117.920000   55.330000 -117.920000   51.790000 -121.460000   51.790000 ;
      POLYGON -117.165000  -59.635000 -113.615000  -63.185000 -117.165000  -63.185000 ;
      POLYGON -117.165000   63.185000 -113.615000   63.185000 -117.165000   59.635000 ;
      POLYGON -117.160000 -102.095000 -114.490000 -104.765000 -117.160000 -104.765000 ;
      POLYGON -117.160000  -98.545000 -113.610000  -98.545000 -113.610000 -102.095000 ;
      POLYGON -117.160000  -80.865000 -114.485000  -83.540000 -117.160000  -83.540000 ;
      POLYGON -116.535000  141.625000 -116.535000  135.905000 -122.255000  135.905000 ;
      POLYGON -116.285000  -78.195000 -113.615000  -78.195000 -113.615000  -80.865000 ;
      POLYGON -116.280000  -56.970000 -113.615000  -56.970000 -113.615000  -59.635000 ;
      POLYGON -116.280000   56.970000 -116.280000   55.330000 -117.920000   55.330000 ;
      POLYGON -116.225000   84.470000 -113.555000   84.470000 -116.225000   81.800000 ;
      POLYGON -116.225000   99.480000 -116.225000   96.810000 -118.895000   96.810000 ;
      POLYGON -116.225000  104.765000 -114.490000  104.765000 -116.225000  103.030000 ;
      POLYGON -116.040000  120.895000 -116.040000  118.035000 -118.900000  118.035000 ;
      POLYGON -115.365000  128.660000 -111.820000  128.660000 -115.365000  125.115000 ;
      POLYGON -115.355000  121.580000 -115.355000  120.895000 -116.040000  120.895000 ;
      POLYGON -115.350000   79.130000 -115.350000   75.620000 -118.860000   75.620000 ;
      POLYGON -115.255000  142.905000 -115.255000  141.625000 -116.535000  141.625000 ;
      POLYGON -114.490000 -125.990000 -110.980000 -129.500000 -114.490000 -129.500000 ;
      POLYGON -114.490000 -122.445000 -110.945000 -122.445000 -110.945000 -125.990000 ;
      POLYGON -114.490000 -104.765000 -111.825000 -107.430000 -114.490000 -107.430000 ;
      POLYGON -114.490000  107.430000 -111.825000  107.430000 -114.490000  104.765000 ;
      POLYGON -114.485000  -83.540000 -110.940000  -87.085000 -114.485000  -87.085000 ;
      POLYGON -113.615000  -80.865000 -110.940000  -80.865000 -110.940000  -83.540000 ;
      POLYGON -113.615000  -63.185000 -112.575000  -64.225000 -113.615000  -64.225000 ;
      POLYGON -113.615000  -59.635000 -110.065000  -59.635000 -110.065000  -63.185000 ;
      POLYGON -113.615000   59.635000 -113.615000   56.970000 -116.280000   56.970000 ;
      POLYGON -113.615000   64.120000 -112.680000   64.120000 -113.615000   63.185000 ;
      POLYGON -113.610000 -102.095000 -110.940000 -102.095000 -110.940000 -104.765000 ;
      POLYGON -113.555000   87.085000 -110.940000   87.085000 -113.555000   84.470000 ;
      POLYGON -112.680000   66.790000 -110.010000   66.790000 -112.680000   64.120000 ;
      POLYGON -112.680000   81.800000 -112.680000   79.130000 -115.350000   79.130000 ;
      POLYGON -112.675000  103.030000 -112.675000   99.480000 -116.225000   99.480000 ;
      POLYGON -112.575000  -64.225000 -110.010000  -66.790000 -112.575000  -66.790000 ;
      POLYGON -111.825000 -107.430000 -108.275000 -110.980000 -111.825000 -110.980000 ;
      POLYGON -111.825000  110.980000 -108.275000  110.980000 -111.825000  107.430000 ;
      POLYGON -111.820000  125.115000 -111.820000  121.580000 -115.355000  121.580000 ;
      POLYGON -111.820000  132.170000 -108.310000  132.170000 -111.820000  128.660000 ;
      POLYGON -110.980000 -129.500000 -107.435000 -133.045000 -110.980000 -133.045000 ;
      POLYGON -110.945000 -125.990000 -107.435000 -125.990000 -107.435000 -129.500000 ;
      POLYGON -110.940000 -104.765000 -108.275000 -104.765000 -108.275000 -107.430000 ;
      POLYGON -110.940000  -87.085000 -109.240000  -88.785000 -110.940000  -88.785000 ;
      POLYGON -110.940000  -83.540000 -107.395000  -83.540000 -107.395000  -87.085000 ;
      POLYGON -110.940000   89.755000 -108.270000   89.755000 -110.940000   87.085000 ;
      POLYGON -110.940000  104.765000 -110.940000  103.030000 -112.675000  103.030000 ;
      POLYGON -110.065000  -63.185000 -109.025000  -63.185000 -109.025000  -64.225000 ;
      POLYGON -110.065000   63.185000 -110.065000   59.635000 -113.615000   59.635000 ;
      POLYGON -110.010000  -66.790000 -107.395000  -69.405000 -110.010000  -69.405000 ;
      POLYGON -110.010000   69.460000 -107.340000   69.460000 -110.010000   66.790000 ;
      POLYGON -110.010000   84.470000 -110.010000   81.800000 -112.680000   81.800000 ;
      POLYGON -110.000000  -45.570000  -92.385000  -63.185000 -110.000000  -63.185000 ;
      POLYGON -110.000000   58.005000  -97.565000   58.005000 -110.000000   45.570000 ;
      POLYGON -109.240000  -88.785000 -105.695000  -92.330000 -109.240000  -92.330000 ;
      POLYGON -109.130000   64.120000 -109.130000   63.185000 -110.065000   63.185000 ;
      POLYGON -109.025000  -64.225000 -106.460000  -64.225000 -106.460000  -66.790000 ;
      POLYGON -108.310000  135.715000 -104.765000  135.715000 -108.310000  132.170000 ;
      POLYGON -108.275000 -110.980000 -104.765000 -114.490000 -108.275000 -114.490000 ;
      POLYGON -108.275000 -107.430000 -104.725000 -107.430000 -104.725000 -110.980000 ;
      POLYGON -108.275000  107.430000 -108.275000  104.765000 -110.940000  104.765000 ;
      POLYGON -108.275000  112.885000 -106.370000  112.885000 -108.275000  110.980000 ;
      POLYGON -108.275000  128.660000 -108.275000  125.115000 -111.820000  125.115000 ;
      POLYGON -108.270000   93.300000 -104.725000   93.300000 -108.270000   89.755000 ;
      POLYGON -107.435000 -133.045000 -103.900000 -136.580000 -107.435000 -136.580000 ;
      POLYGON -107.435000 -129.500000 -103.890000 -129.500000 -103.890000 -133.045000 ;
      POLYGON -107.395000  -87.085000 -105.695000  -87.085000 -105.695000  -88.785000 ;
      POLYGON -107.395000  -69.405000 -104.820000  -71.980000 -107.395000  -71.980000 ;
      POLYGON -107.395000   87.085000 -107.395000   84.470000 -110.010000   84.470000 ;
      POLYGON -107.340000   73.010000 -103.790000   73.010000 -107.340000   69.460000 ;
      POLYGON -106.465000   88.015000 -106.465000   87.085000 -107.395000   87.085000 ;
      POLYGON -106.460000  -66.790000 -103.845000  -66.790000 -103.845000  -69.405000 ;
      POLYGON -106.460000   66.790000 -106.460000   64.120000 -109.130000   64.120000 ;
      POLYGON -106.370000  116.225000 -103.030000  116.225000 -106.370000  112.885000 ;
      POLYGON -105.695000  -92.330000 -102.150000  -95.875000 -105.695000  -95.875000 ;
      POLYGON -105.695000  -88.785000 -102.150000  -88.785000 -102.150000  -92.330000 ;
      POLYGON -104.820000  -71.980000 -102.150000  -74.650000 -104.820000  -74.650000 ;
      POLYGON -104.765000 -114.490000 -103.030000 -116.225000 -104.765000 -116.225000 ;
      POLYGON -104.765000  132.170000 -104.765000  128.660000 -108.275000  128.660000 ;
      POLYGON -104.765000  139.260000 -101.220000  139.260000 -104.765000  135.715000 ;
      POLYGON -104.725000 -110.980000 -101.215000 -110.980000 -101.215000 -114.490000 ;
      POLYGON -104.725000   89.755000 -104.725000   88.015000 -106.465000   88.015000 ;
      POLYGON -104.725000   96.810000 -101.215000   96.810000 -104.725000   93.300000 ;
      POLYGON -104.725000  110.980000 -104.725000  107.430000 -108.275000  107.430000 ;
      POLYGON -103.900000 -136.580000 -100.355000 -140.125000 -103.900000 -140.125000 ;
      POLYGON -103.890000 -133.045000 -100.355000 -133.045000 -100.355000 -136.580000 ;
      POLYGON -103.845000  -69.405000 -101.270000  -69.405000 -101.270000  -71.980000 ;
      POLYGON -103.790000   69.460000 -103.790000   66.790000 -106.460000   66.790000 ;
      POLYGON -103.790000   75.620000 -101.180000   75.620000 -103.790000   73.010000 ;
      POLYGON -103.030000 -116.225000  -99.480000 -119.775000 -103.030000 -119.775000 ;
      POLYGON -103.030000  119.615000  -99.640000  119.615000 -103.030000  116.225000 ;
      POLYGON -102.820000  112.885000 -102.820000  110.980000 -104.725000  110.980000 ;
      POLYGON -102.150000  -95.875000  -99.480000  -98.545000 -102.150000  -98.545000 ;
      POLYGON -102.150000  -92.330000  -98.605000  -92.330000  -98.605000  -95.875000 ;
      POLYGON -102.150000  -74.650000 -100.340000  -76.460000 -102.150000  -76.460000 ;
      POLYGON -102.150000   92.330000 -102.150000   89.755000 -104.725000   89.755000 ;
      POLYGON -101.525000  156.635000 -101.525000  142.905000 -115.255000  142.905000 ;
      POLYGON -101.270000  -71.980000  -98.600000  -71.980000  -98.600000  -74.650000 ;
      POLYGON -101.220000  135.715000 -101.220000  132.170000 -104.765000  132.170000 ;
      POLYGON -101.220000  142.795000  -97.685000  142.795000 -101.220000  139.260000 ;
      POLYGON -101.215000 -114.490000  -99.480000 -114.490000  -99.480000 -116.225000 ;
      POLYGON -101.215000   99.480000  -98.545000   99.480000 -101.215000   96.810000 ;
      POLYGON -101.180000   79.130000  -97.670000   79.130000 -101.180000   75.620000 ;
      POLYGON -101.180000   93.300000 -101.180000   92.330000 -102.150000   92.330000 ;
      POLYGON -100.355000 -157.805000  -82.765000 -157.805000  -82.765000 -175.395000 ;
      POLYGON -100.355000 -140.125000  -96.810000 -143.670000 -100.355000 -143.670000 ;
      POLYGON -100.355000 -136.580000  -96.810000 -136.580000  -96.810000 -140.125000 ;
      POLYGON -100.340000  -76.460000  -97.670000  -79.130000 -100.340000  -79.130000 ;
      POLYGON -100.245000  157.915000 -100.245000  156.635000 -101.525000  156.635000 ;
      POLYGON -100.240000   73.010000 -100.240000   69.460000 -103.790000   69.460000 ;
      POLYGON  -99.640000  122.445000  -96.810000  122.445000  -99.640000  119.615000 ;
      POLYGON  -99.480000 -119.775000  -96.810000 -122.445000  -99.480000 -122.445000 ;
      POLYGON  -99.480000 -116.225000  -95.930000 -116.225000  -95.930000 -119.775000 ;
      POLYGON  -99.480000  -98.545000  -96.805000 -101.220000  -99.480000 -101.220000 ;
      POLYGON  -99.480000  116.225000  -99.480000  112.885000 -102.820000  112.885000 ;
      POLYGON  -98.605000  -95.875000  -95.935000  -95.875000  -95.935000  -98.545000 ;
      POLYGON  -98.600000  -74.650000  -96.790000  -74.650000  -96.790000  -76.460000 ;
      POLYGON  -98.545000  102.150000  -95.875000  102.150000  -98.545000   99.480000 ;
      POLYGON  -97.685000  146.340000  -94.140000  146.340000  -97.685000  142.795000 ;
      POLYGON  -97.675000  139.260000  -97.675000  135.715000 -101.220000  135.715000 ;
      POLYGON  -97.670000  -79.130000  -95.000000  -81.800000  -97.670000  -81.800000 ;
      POLYGON  -97.670000   81.800000  -95.000000   81.800000  -97.670000   79.130000 ;
      POLYGON  -97.670000   96.810000  -97.670000   93.300000 -101.180000   93.300000 ;
      POLYGON  -97.630000   75.620000  -97.630000   73.010000 -100.240000   73.010000 ;
      POLYGON  -97.565000   75.620000  -79.950000   75.620000  -97.565000   58.005000 ;
      POLYGON  -96.810000 -143.670000  -93.300000 -147.180000  -96.810000 -147.180000 ;
      POLYGON  -96.810000 -140.125000  -93.265000 -140.125000  -93.265000 -143.670000 ;
      POLYGON  -96.810000 -122.445000  -94.145000 -125.110000  -96.810000 -125.110000 ;
      POLYGON  -96.810000  125.110000  -94.145000  125.110000  -96.810000  122.445000 ;
      POLYGON  -96.805000 -101.220000  -93.260000 -104.765000  -96.805000 -104.765000 ;
      POLYGON  -96.790000  -76.460000  -94.120000  -76.460000  -94.120000  -79.130000 ;
      POLYGON  -96.090000  119.615000  -96.090000  116.225000  -99.480000  116.225000 ;
      POLYGON  -95.985000  162.175000  -95.985000  157.915000 -100.245000  157.915000 ;
      POLYGON  -95.935000  -98.545000  -93.260000  -98.545000  -93.260000 -101.220000 ;
      POLYGON  -95.930000 -119.775000  -93.260000 -119.775000  -93.260000 -122.445000 ;
      POLYGON  -95.875000  104.765000  -93.260000  104.765000  -95.875000  102.150000 ;
      POLYGON  -95.310000  141.625000  -95.310000  139.260000  -97.675000  139.260000 ;
      POLYGON  -95.000000  -81.800000  -92.330000  -84.470000  -95.000000  -84.470000 ;
      POLYGON  -95.000000   84.470000  -92.330000   84.470000  -95.000000   81.800000 ;
      POLYGON  -95.000000   99.480000  -95.000000   96.810000  -97.670000   96.810000 ;
      POLYGON  -94.995000  120.710000  -94.995000  119.615000  -96.090000  119.615000 ;
      POLYGON  -94.145000 -125.110000  -90.595000 -128.660000  -94.145000 -128.660000 ;
      POLYGON  -94.145000  128.660000  -90.595000  128.660000  -94.145000  125.110000 ;
      POLYGON  -94.140000  142.795000  -94.140000  141.625000  -95.310000  141.625000 ;
      POLYGON  -94.140000  149.850000  -90.630000  149.850000  -94.140000  146.340000 ;
      POLYGON  -94.120000  -79.130000  -92.385000  -79.130000  -92.385000  -80.865000 ;
      POLYGON  -94.120000   79.130000  -94.120000   75.620000  -97.630000   75.620000 ;
      POLYGON  -93.300000 -147.180000  -89.755000 -150.725000  -93.300000 -150.725000 ;
      POLYGON  -93.265000 -143.670000  -89.755000 -143.670000  -89.755000 -147.180000 ;
      POLYGON  -93.260000 -122.445000  -90.595000 -122.445000  -90.595000 -125.110000 ;
      POLYGON  -93.260000 -104.765000  -91.560000 -106.465000  -93.260000 -106.465000 ;
      POLYGON  -93.260000 -101.220000  -89.715000 -101.220000  -89.715000 -104.765000 ;
      POLYGON  -93.260000  107.435000  -90.590000  107.435000  -93.260000  104.765000 ;
      POLYGON  -93.260000  122.445000  -93.260000  120.710000  -94.995000  120.710000 ;
      POLYGON  -92.385000  -80.865000  -91.450000  -80.865000  -91.450000  -81.800000 ;
      POLYGON  -92.385000  -63.185000  -74.705000  -80.865000  -92.385000  -80.865000 ;
      POLYGON  -92.330000  -84.470000  -89.715000  -87.085000  -92.330000  -87.085000 ;
      POLYGON  -92.330000   87.140000  -89.660000   87.140000  -92.330000   84.470000 ;
      POLYGON  -92.330000  102.150000  -92.330000   99.480000  -95.000000   99.480000 ;
      POLYGON  -91.560000 -106.465000  -88.015000 -110.010000  -91.560000 -110.010000 ;
      POLYGON  -91.450000  -81.800000  -88.780000  -81.800000  -88.780000  -84.470000 ;
      POLYGON  -91.450000   81.800000  -91.450000   79.130000  -94.120000   79.130000 ;
      POLYGON  -90.630000  153.395000  -87.085000  153.395000  -90.630000  149.850000 ;
      POLYGON  -90.595000 -128.660000  -87.085000 -132.170000  -90.595000 -132.170000 ;
      POLYGON  -90.595000 -125.110000  -87.045000 -125.110000  -87.045000 -128.660000 ;
      POLYGON  -90.595000  125.110000  -90.595000  122.445000  -93.260000  122.445000 ;
      POLYGON  -90.595000  132.155000  -87.100000  132.155000  -90.595000  128.660000 ;
      POLYGON  -90.595000  146.340000  -90.595000  142.795000  -94.140000  142.795000 ;
      POLYGON  -90.590000  110.010000  -88.015000  110.010000  -90.590000  107.435000 ;
      POLYGON  -89.755000 -150.725000  -86.220000 -154.260000  -89.755000 -154.260000 ;
      POLYGON  -89.755000 -147.180000  -86.210000 -147.180000  -86.210000 -150.725000 ;
      POLYGON  -89.715000 -104.765000  -88.015000 -104.765000  -88.015000 -106.465000 ;
      POLYGON  -89.715000  -87.085000  -87.140000  -89.660000  -89.715000  -89.660000 ;
      POLYGON  -89.715000  104.765000  -89.715000  102.150000  -92.330000  102.150000 ;
      POLYGON  -89.660000   90.690000  -86.110000   90.690000  -89.660000   87.140000 ;
      POLYGON  -89.090000  126.615000  -89.090000  125.110000  -90.595000  125.110000 ;
      POLYGON  -88.785000  105.695000  -88.785000  104.765000  -89.715000  104.765000 ;
      POLYGON  -88.780000  -84.470000  -86.165000  -84.470000  -86.165000  -87.085000 ;
      POLYGON  -88.780000   84.470000  -88.780000   81.800000  -91.450000   81.800000 ;
      POLYGON  -88.120000  170.040000  -88.120000  162.175000  -95.985000  162.175000 ;
      POLYGON  -88.015000 -110.010000  -84.470000 -113.555000  -88.015000 -113.555000 ;
      POLYGON  -88.015000 -106.465000  -84.470000 -106.465000  -84.470000 -110.010000 ;
      POLYGON  -88.015000  112.885000  -85.140000  112.885000  -88.015000  110.010000 ;
      POLYGON  -87.140000  -89.660000  -84.470000  -92.330000  -87.140000  -92.330000 ;
      POLYGON  -87.100000  134.840000  -84.415000  134.840000  -87.100000  132.155000 ;
      POLYGON  -87.085000 -132.170000  -84.625000 -134.630000  -87.085000 -134.630000 ;
      POLYGON  -87.085000  149.850000  -87.085000  146.340000  -90.595000  146.340000 ;
      POLYGON  -87.085000  156.940000  -83.540000  156.940000  -87.085000  153.395000 ;
      POLYGON  -87.045000 -128.660000  -83.535000 -128.660000  -83.535000 -132.170000 ;
      POLYGON  -87.045000  107.435000  -87.045000  105.695000  -88.785000  105.695000 ;
      POLYGON  -87.045000  128.660000  -87.045000  126.615000  -89.090000  126.615000 ;
      POLYGON  -86.220000 -154.260000  -82.675000 -157.805000  -86.220000 -157.805000 ;
      POLYGON  -86.210000 -150.725000  -82.675000 -150.725000  -82.675000 -154.260000 ;
      POLYGON  -86.165000  -87.085000  -83.590000  -87.085000  -83.590000  -89.660000 ;
      POLYGON  -86.110000   87.140000  -86.110000   84.470000  -88.780000   84.470000 ;
      POLYGON  -86.110000   93.300000  -83.500000   93.300000  -86.110000   90.690000 ;
      POLYGON  -85.140000  116.225000  -81.800000  116.225000  -85.140000  112.885000 ;
      POLYGON  -84.625000 -134.630000  -81.800000 -137.455000  -84.625000 -137.455000 ;
      POLYGON  -84.470000 -113.555000  -81.800000 -116.225000  -84.470000 -116.225000 ;
      POLYGON  -84.470000 -110.010000  -80.925000 -110.010000  -80.925000 -113.555000 ;
      POLYGON  -84.470000  -92.330000  -82.660000  -94.140000  -84.470000  -94.140000 ;
      POLYGON  -84.470000  110.010000  -84.470000  107.435000  -87.045000  107.435000 ;
      POLYGON  -84.415000  138.390000  -80.865000  138.390000  -84.415000  134.840000 ;
      POLYGON  -83.590000  -89.660000  -80.920000  -89.660000  -80.920000  -92.330000 ;
      POLYGON  -83.550000  132.155000  -83.550000  128.660000  -87.045000  128.660000 ;
      POLYGON  -83.540000  153.395000  -83.540000  149.850000  -87.085000  149.850000 ;
      POLYGON  -83.540000  160.475000  -80.005000  160.475000  -83.540000  156.940000 ;
      POLYGON  -83.535000 -132.170000  -81.075000 -132.170000  -81.075000 -134.630000 ;
      POLYGON  -83.500000   96.810000  -79.990000   96.810000  -83.500000   93.300000 ;
      POLYGON  -82.765000 -175.395000  -75.620000 -175.395000  -75.620000 -182.540000 ;
      POLYGON  -82.675000 -157.805000  -79.130000 -161.350000  -82.675000 -161.350000 ;
      POLYGON  -82.675000 -154.260000  -79.130000 -154.260000  -79.130000 -157.805000 ;
      POLYGON  -82.660000  -94.140000  -79.990000  -96.810000  -82.660000  -96.810000 ;
      POLYGON  -82.560000   90.690000  -82.560000   87.140000  -86.110000   87.140000 ;
      POLYGON  -81.800000 -137.455000  -79.130000 -140.125000  -81.800000 -140.125000 ;
      POLYGON  -81.800000 -116.225000  -79.125000 -118.900000  -81.800000 -118.900000 ;
      POLYGON  -81.800000  119.615000  -78.410000  119.615000  -81.800000  116.225000 ;
      POLYGON  -81.595000  112.885000  -81.595000  110.010000  -84.470000  110.010000 ;
      POLYGON  -81.075000 -134.630000  -78.250000 -134.630000  -78.250000 -137.455000 ;
      POLYGON  -80.925000 -113.555000  -78.255000 -113.555000  -78.255000 -116.225000 ;
      POLYGON  -80.920000  -92.330000  -79.110000  -92.330000  -79.110000  -94.140000 ;
      POLYGON  -80.865000  134.840000  -80.865000  132.155000  -83.550000  132.155000 ;
      POLYGON  -80.865000  140.125000  -79.130000  140.125000  -80.865000  138.390000 ;
      POLYGON  -80.300000  156.635000  -80.300000  153.395000  -83.540000  153.395000 ;
      POLYGON  -80.005000  164.020000  -76.460000  164.020000  -80.005000  160.475000 ;
      POLYGON  -79.995000  156.940000  -79.995000  156.635000  -80.300000  156.635000 ;
      POLYGON  -79.990000  -96.810000  -77.320000  -99.480000  -79.990000  -99.480000 ;
      POLYGON  -79.990000   99.480000  -77.320000   99.480000  -79.990000   96.810000 ;
      POLYGON  -79.950000   92.330000  -63.240000   92.330000  -79.950000   75.620000 ;
      POLYGON  -79.950000   93.300000  -79.950000   90.690000  -82.560000   90.690000 ;
      POLYGON  -79.130000 -161.350000  -75.620000 -164.860000  -79.130000 -164.860000 ;
      POLYGON  -79.130000 -157.805000  -75.585000 -157.805000  -75.585000 -161.350000 ;
      POLYGON  -79.130000 -140.125000  -76.350000 -142.905000  -79.130000 -142.905000 ;
      POLYGON  -79.130000  142.790000  -76.465000  142.790000  -79.130000  140.125000 ;
      POLYGON  -79.125000 -118.900000  -75.580000 -122.445000  -79.125000 -122.445000 ;
      POLYGON  -79.110000  -94.140000  -76.440000  -94.140000  -76.440000  -96.810000 ;
      POLYGON  -78.410000  122.445000  -75.580000  122.445000  -78.410000  119.615000 ;
      POLYGON  -78.255000 -116.225000  -75.580000 -116.225000  -75.580000 -118.900000 ;
      POLYGON  -78.255000  116.225000  -78.255000  112.885000  -81.595000  112.885000 ;
      POLYGON  -78.250000 -137.455000  -75.580000 -137.455000  -75.580000 -140.125000 ;
      POLYGON  -77.320000  -99.480000  -74.650000 -102.150000  -77.320000 -102.150000 ;
      POLYGON  -77.320000  102.150000  -74.650000  102.150000  -77.320000   99.480000 ;
      POLYGON  -77.315000  138.390000  -77.315000  134.840000  -80.865000  134.840000 ;
      POLYGON  -76.465000  145.375000  -73.880000  145.375000  -76.465000  142.790000 ;
      POLYGON  -76.460000  160.475000  -76.460000  156.940000  -79.995000  156.940000 ;
      POLYGON  -76.460000  167.530000  -72.950000  167.530000  -76.460000  164.020000 ;
      POLYGON  -76.440000  -96.810000  -74.705000  -96.810000  -74.705000  -98.545000 ;
      POLYGON  -76.440000   96.810000  -76.440000   93.300000  -79.950000   93.300000 ;
      POLYGON  -76.350000 -142.905000  -72.915000 -146.340000  -76.350000 -146.340000 ;
      POLYGON  -75.620000 -164.860000  -72.950000 -167.530000  -75.620000 -167.530000 ;
      POLYGON  -75.620000  182.540000  -75.620000  170.040000  -88.120000  170.040000 ;
      POLYGON  -75.585000 -161.350000  -72.075000 -161.350000  -72.075000 -164.860000 ;
      POLYGON  -75.580000 -140.125000  -72.800000 -140.125000  -72.800000 -142.905000 ;
      POLYGON  -75.580000 -122.445000  -73.015000 -125.010000  -75.580000 -125.010000 ;
      POLYGON  -75.580000 -118.900000  -72.035000 -118.900000  -72.035000 -122.445000 ;
      POLYGON  -75.580000  125.115000  -72.910000  125.115000  -75.580000  122.445000 ;
      POLYGON  -75.580000  140.125000  -75.580000  138.390000  -77.315000  138.390000 ;
      POLYGON  -74.865000  119.615000  -74.865000  116.225000  -78.255000  116.225000 ;
      POLYGON  -74.705000  -98.545000  -73.770000  -98.545000  -73.770000  -99.480000 ;
      POLYGON  -74.705000  -80.865000  -57.025000  -98.545000  -74.705000  -98.545000 ;
      POLYGON  -74.650000 -102.150000  -72.035000 -104.765000  -74.650000 -104.765000 ;
      POLYGON  -74.650000  104.820000  -71.980000  104.820000  -74.650000  102.150000 ;
      POLYGON  -73.880000  148.445000  -70.810000  148.445000  -73.880000  145.375000 ;
      POLYGON  -73.770000  -99.480000  -71.100000  -99.480000  -71.100000 -102.150000 ;
      POLYGON  -73.770000   99.480000  -73.770000   96.810000  -76.440000   96.810000 ;
      POLYGON  -73.015000 -125.010000  -70.125000 -127.900000  -73.015000 -127.900000 ;
      POLYGON  -72.950000 -167.530000  -70.440000 -170.040000  -72.950000 -170.040000 ;
      POLYGON  -72.950000  170.040000  -70.440000  170.040000  -72.950000  167.530000 ;
      POLYGON  -72.915000 -146.340000  -69.405000 -149.850000  -72.915000 -149.850000 ;
      POLYGON  -72.915000  142.790000  -72.915000  140.125000  -75.580000  140.125000 ;
      POLYGON  -72.915000  164.020000  -72.915000  160.475000  -76.460000  160.475000 ;
      POLYGON  -72.910000  128.660000  -69.365000  128.660000  -72.910000  125.115000 ;
      POLYGON  -72.800000 -142.905000  -69.365000 -142.905000  -69.365000 -146.340000 ;
      POLYGON  -72.075000 -164.860000  -69.405000 -164.860000  -69.405000 -167.530000 ;
      POLYGON  -72.035000 -122.445000  -69.470000 -122.445000  -69.470000 -125.010000 ;
      POLYGON  -72.035000 -104.765000  -69.460000 -107.340000  -72.035000 -107.340000 ;
      POLYGON  -72.035000  122.445000  -72.035000  119.615000  -74.865000  119.615000 ;
      POLYGON  -71.980000  108.370000  -68.430000  108.370000  -71.980000  104.820000 ;
      POLYGON  -71.105000  123.375000  -71.105000  122.445000  -72.035000  122.445000 ;
      POLYGON  -71.100000 -102.150000  -68.485000 -102.150000  -68.485000 -104.765000 ;
      POLYGON  -71.100000  102.150000  -71.100000   99.480000  -73.770000   99.480000 ;
      POLYGON  -70.810000  151.585000  -67.670000  151.585000  -70.810000  148.445000 ;
      POLYGON  -70.330000  145.375000  -70.330000  142.790000  -72.915000  142.790000 ;
      POLYGON  -70.125000 -127.900000  -66.790000 -131.235000  -70.125000 -131.235000 ;
      POLYGON  -69.470000 -125.010000  -66.580000 -125.010000  -66.580000 -127.900000 ;
      POLYGON  -69.460000 -107.340000  -66.790000 -110.010000  -69.460000 -110.010000 ;
      POLYGON  -69.405000 -149.850000  -67.670000 -151.585000  -69.405000 -151.585000 ;
      POLYGON  -69.405000  167.530000  -69.405000  164.020000  -72.915000  164.020000 ;
      POLYGON  -69.365000 -146.340000  -65.855000 -146.340000  -65.855000 -149.850000 ;
      POLYGON  -69.365000  125.115000  -69.365000  123.375000  -71.105000  123.375000 ;
      POLYGON  -69.365000  132.155000  -65.870000  132.155000  -69.365000  128.660000 ;
      POLYGON  -68.485000 -104.765000  -65.910000 -104.765000  -65.910000 -107.340000 ;
      POLYGON  -68.430000  104.820000  -68.430000  102.150000  -71.100000  102.150000 ;
      POLYGON  -68.430000  111.820000  -64.980000  111.820000  -68.430000  108.370000 ;
      POLYGON  -67.865000  126.615000  -67.865000  125.115000  -69.365000  125.115000 ;
      POLYGON  -67.670000 -151.585000  -64.225000 -155.030000  -67.670000 -155.030000 ;
      POLYGON  -67.670000  155.030000  -64.225000  155.030000  -67.670000  151.585000 ;
      POLYGON  -67.260000  148.445000  -67.260000  145.375000  -70.330000  145.375000 ;
      POLYGON  -66.790000 -131.235000  -63.395000 -134.630000  -66.790000 -134.630000 ;
      POLYGON  -66.790000 -110.010000  -64.980000 -111.820000  -66.790000 -111.820000 ;
      POLYGON  -66.580000 -127.900000  -63.245000 -127.900000  -63.245000 -131.235000 ;
      POLYGON  -65.910000 -107.340000  -63.240000 -107.340000  -63.240000 -110.010000 ;
      POLYGON  -65.870000  134.625000  -63.400000  134.625000  -65.870000  132.155000 ;
      POLYGON  -65.855000 -149.850000  -64.120000 -149.850000  -64.120000 -151.585000 ;
      POLYGON  -65.820000  128.660000  -65.820000  126.615000  -67.865000  126.615000 ;
      POLYGON  -64.980000 -111.820000  -62.310000 -114.490000  -64.980000 -114.490000 ;
      POLYGON  -64.980000  115.355000  -61.445000  115.355000  -64.980000  111.820000 ;
      POLYGON  -64.880000  108.370000  -64.880000  104.820000  -68.430000  104.820000 ;
      POLYGON  -64.120000 -151.585000  -63.185000 -151.585000  -63.185000 -152.520000 ;
      POLYGON  -64.120000  151.585000  -64.120000  148.445000  -67.260000  148.445000 ;
      POLYGON  -63.400000  137.510000  -60.515000  137.510000  -63.400000  134.625000 ;
      POLYGON  -63.395000 -134.630000  -60.515000 -137.510000  -63.395000 -137.510000 ;
      POLYGON  -63.245000 -131.235000  -59.850000 -131.235000  -59.850000 -134.630000 ;
      POLYGON  -63.240000 -110.010000  -61.430000 -110.010000  -61.430000 -111.820000 ;
      POLYGON  -63.240000  110.000000  -45.570000  110.000000  -63.240000   92.330000 ;
      POLYGON  -63.240000  110.010000  -63.240000  108.370000  -64.880000  108.370000 ;
      POLYGON  -63.185000  152.520000  -63.185000  151.585000  -64.120000  151.585000 ;
      POLYGON  -62.325000  132.155000  -62.325000  128.660000  -65.820000  128.660000 ;
      POLYGON  -62.310000 -114.490000  -59.640000 -117.160000  -62.310000 -117.160000 ;
      POLYGON  -61.445000  118.425000  -58.375000  118.425000  -61.445000  115.355000 ;
      POLYGON  -61.430000 -111.820000  -58.760000 -111.820000  -58.760000 -114.490000 ;
      POLYGON  -61.430000  111.820000  -61.430000  110.010000  -63.240000  110.010000 ;
      POLYGON  -60.515000 -137.510000  -58.005000 -140.020000  -60.515000 -140.020000 ;
      POLYGON  -60.515000  140.020000  -58.005000  140.020000  -60.515000  137.510000 ;
      POLYGON  -59.855000  134.625000  -59.855000  132.155000  -62.325000  132.155000 ;
      POLYGON  -59.850000 -134.630000  -56.970000 -134.630000  -56.970000 -137.510000 ;
      POLYGON  -59.640000 -117.160000  -56.970000 -119.830000  -59.640000 -119.830000 ;
      POLYGON  -58.760000 -114.490000  -56.090000 -114.490000  -56.090000 -117.160000 ;
      POLYGON  -58.375000  121.470000  -55.330000  121.470000  -58.375000  118.425000 ;
      POLYGON  -57.895000  115.355000  -57.895000  111.820000  -61.430000  111.820000 ;
      POLYGON  -57.025000  -98.545000  -45.570000 -110.000000  -57.025000 -110.000000 ;
      POLYGON  -56.970000 -119.830000  -54.355000 -122.445000  -56.970000 -122.445000 ;
      POLYGON  -56.970000  137.510000  -56.970000  134.625000  -59.855000  134.625000 ;
      POLYGON  -56.090000 -117.160000  -53.420000 -117.160000  -53.420000 -119.830000 ;
      POLYGON  -55.330000  125.010000  -51.790000  125.010000  -55.330000  121.470000 ;
      POLYGON  -54.825000  118.425000  -54.825000  115.355000  -57.895000  115.355000 ;
      POLYGON  -54.355000 -122.445000  -51.790000 -125.010000  -54.355000 -125.010000 ;
      POLYGON  -53.420000 -119.830000  -50.805000 -119.830000  -50.805000 -122.445000 ;
      POLYGON  -51.780000  121.470000  -51.780000  118.425000  -54.825000  118.425000 ;
      POLYGON  -50.805000 -122.445000  -50.750000 -122.445000  -50.750000 -122.500000 ;
      POLYGON  -50.750000  122.500000  -50.750000  121.470000  -51.780000  121.470000 ;
      POLYGON  -11.900000 -181.440000  -10.800000 -181.440000  -11.900000 -182.540000 ;
      POLYGON  -11.900000 -170.040000  -10.800000 -171.140000  -11.900000 -171.140000 ;
      POLYGON  -11.900000 -151.420000  -10.800000 -151.420000  -11.900000 -152.520000 ;
      POLYGON  -11.900000 -140.020000  -10.800000 -141.120000  -11.900000 -141.120000 ;
      POLYGON  -11.340000  126.110000  -10.240000  126.110000  -11.340000  125.010000 ;
      POLYGON  -11.340000  137.510000  -10.240000  136.410000  -11.340000  136.410000 ;
      POLYGON  -11.340000  156.130000  -10.240000  156.130000  -11.340000  155.030000 ;
      POLYGON  -11.340000  167.530000  -10.240000  166.430000  -11.340000  166.430000 ;
      POLYGON  -10.075000 -167.530000   -7.565000 -167.530000   -7.565000 -170.040000 ;
      POLYGON  -10.075000 -137.510000   -7.565000 -137.510000   -7.565000 -140.020000 ;
      POLYGON   -7.565000 -170.040000    4.935000 -170.040000    4.935000 -182.540000 ;
      POLYGON   -7.565000 -140.020000   -7.460000 -140.020000   -7.460000 -140.125000 ;
      POLYGON   -7.565000  125.010000   -7.565000  122.500000  -10.075000  122.500000 ;
      POLYGON   -7.565000  155.030000   -7.565000  152.520000  -10.075000  152.520000 ;
      POLYGON   -7.460000 -140.125000    4.935000 -140.125000    4.935000 -152.520000 ;
      POLYGON   -4.895000 -155.030000   10.115000 -170.040000   -4.895000 -170.040000 ;
      POLYGON   -4.895000 -125.010000   10.115000 -140.020000   -4.895000 -140.020000 ;
      POLYGON   -4.895000  114.490000   -0.405000  114.490000   -4.895000  110.000000 ;
      POLYGON   -4.895000  146.340000    1.425000  146.340000   -4.895000  140.020000 ;
      POLYGON   -0.405000  125.010000   10.115000  125.010000   -0.405000  114.490000 ;
      POLYGON   -0.405000  132.170000   -0.405000  125.010000   -7.565000  125.010000 ;
      POLYGON    1.425000  155.030000   10.115000  155.030000    1.425000  146.340000 ;
      POLYGON    1.425000  164.020000    1.425000  155.030000   -7.565000  155.030000 ;
      POLYGON    2.265000  134.840000    2.265000  132.170000   -0.405000  132.170000 ;
      POLYGON    4.935000  137.510000    4.935000  134.840000    2.265000  134.840000 ;
      POLYGON    4.935000  167.530000    4.935000  164.020000    1.425000  164.020000 ;
      POLYGON   11.455000 -166.430000   12.555000 -166.430000   12.555000 -167.530000 ;
      POLYGON   11.455000 -136.410000   12.555000 -136.410000   12.555000 -137.510000 ;
      POLYGON   12.015000  111.100000   13.115000  111.100000   13.115000  110.000000 ;
      POLYGON   12.015000  141.120000   13.115000  141.120000   13.115000  140.020000 ;
      POLYGON   12.555000 -155.030000   12.555000 -156.130000   11.455000 -156.130000 ;
      POLYGON   12.555000 -125.010000   12.555000 -126.110000   11.455000 -126.110000 ;
      POLYGON   13.115000  122.500000   13.115000  121.400000   12.015000  121.400000 ;
      POLYGON   13.115000  152.520000   13.115000  151.420000   12.015000  151.420000 ;
      POLYGON   45.570000  110.000000   63.240000  110.000000   63.240000   92.330000 ;
      POLYGON   50.750000 -119.830000   53.420000 -119.830000   50.750000 -122.500000 ;
      POLYGON   50.750000 -104.820000   50.750000 -110.000000   45.570000 -110.000000 ;
      POLYGON   50.750000  122.500000   51.780000  121.470000   50.750000  121.470000 ;
      POLYGON   51.780000  121.470000   53.420000  119.830000   51.780000  119.830000 ;
      POLYGON   51.790000  125.010000   54.300000  125.010000   54.300000  122.500000 ;
      POLYGON   53.420000 -117.160000   56.090000 -117.160000   53.420000 -119.830000 ;
      POLYGON   53.420000  119.830000   56.090000  117.160000   53.420000  117.160000 ;
      POLYGON   54.300000 -122.500000   54.300000 -125.010000   51.790000 -125.010000 ;
      POLYGON   54.300000  122.500000   55.330000  122.500000   55.330000  121.470000 ;
      POLYGON   55.330000  121.470000   56.970000  121.470000   56.970000  119.830000 ;
      POLYGON   56.090000 -114.490000   58.760000 -114.490000   56.090000 -117.160000 ;
      POLYGON   56.090000  117.160000   58.760000  114.490000   56.090000  114.490000 ;
      POLYGON   56.970000 -134.840000   59.640000 -134.840000   56.970000 -137.510000 ;
      POLYGON   56.970000 -119.830000   56.970000 -122.500000   54.300000 -122.500000 ;
      POLYGON   56.970000  119.830000   59.640000  119.830000   59.640000  117.160000 ;
      POLYGON   56.970000  137.510000   60.515000  133.965000   56.970000  133.965000 ;
      POLYGON   57.025000  -98.545000   57.025000 -104.820000   50.750000 -104.820000 ;
      POLYGON   58.005000  140.020000   60.515000  140.020000   60.515000  137.510000 ;
      POLYGON   58.760000 -111.820000   61.430000 -111.820000   58.760000 -114.490000 ;
      POLYGON   58.760000  114.490000   62.270000  110.980000   58.760000  110.980000 ;
      POLYGON   59.640000 -132.170000   62.310000 -132.170000   59.640000 -134.840000 ;
      POLYGON   59.640000 -117.160000   59.640000 -119.830000   56.970000 -119.830000 ;
      POLYGON   59.640000  117.160000   62.310000  117.160000   62.310000  114.490000 ;
      POLYGON   60.515000 -137.510000   60.515000 -140.020000   58.005000 -140.020000 ;
      POLYGON   60.515000  133.965000   63.245000  131.235000   60.515000  131.235000 ;
      POLYGON   60.515000  137.510000   64.060000  137.510000   64.060000  133.965000 ;
      POLYGON   61.430000 -108.370000   64.880000 -108.370000   61.430000 -111.820000 ;
      POLYGON   62.270000  110.980000   63.240000  110.010000   62.270000  110.010000 ;
      POLYGON   62.310000 -128.660000   65.820000 -128.660000   62.310000 -132.170000 ;
      POLYGON   62.310000 -114.490000   62.310000 -117.160000   59.640000 -117.160000 ;
      POLYGON   62.310000  114.490000   65.820000  114.490000   65.820000  110.980000 ;
      POLYGON   63.185000 -149.850000   65.855000 -149.850000   63.185000 -152.520000 ;
      POLYGON   63.185000 -134.840000   63.185000 -137.510000   60.515000 -137.510000 ;
      POLYGON   63.185000  152.520000   64.120000  151.585000   63.185000  151.585000 ;
      POLYGON   63.240000   92.330000   79.950000   92.330000   79.950000   75.620000 ;
      POLYGON   63.240000  110.010000   65.910000  107.340000   63.240000  107.340000 ;
      POLYGON   63.245000  131.235000   66.790000  127.690000   63.245000  127.690000 ;
      POLYGON   64.060000  133.965000   66.790000  133.965000   66.790000  131.235000 ;
      POLYGON   64.120000  151.585000   65.855000  149.850000   64.120000  149.850000 ;
      POLYGON   64.225000  155.030000   66.735000  155.030000   66.735000  152.520000 ;
      POLYGON   64.880000 -104.820000   68.430000 -104.820000   64.880000 -108.370000 ;
      POLYGON   64.980000 -111.820000   64.980000 -114.490000   62.310000 -114.490000 ;
      POLYGON   65.820000 -125.115000   69.365000 -125.115000   65.820000 -128.660000 ;
      POLYGON   65.820000  110.980000   66.790000  110.980000   66.790000  110.010000 ;
      POLYGON   65.855000 -146.340000   69.365000 -146.340000   65.855000 -149.850000 ;
      POLYGON   65.855000 -132.170000   65.855000 -134.840000   63.185000 -134.840000 ;
      POLYGON   65.855000  149.850000   69.365000  146.340000   65.855000  146.340000 ;
      POLYGON   65.910000  107.340000   69.460000  103.790000   65.910000  103.790000 ;
      POLYGON   66.735000 -152.520000   66.735000 -155.030000   64.225000 -155.030000 ;
      POLYGON   66.735000  152.520000   67.670000  152.520000   67.670000  151.585000 ;
      POLYGON   66.790000  110.010000   69.460000  110.010000   69.460000  107.340000 ;
      POLYGON   66.790000  127.690000   70.335000  124.145000   66.790000  124.145000 ;
      POLYGON   66.790000  131.235000   70.335000  131.235000   70.335000  127.690000 ;
      POLYGON   67.670000  151.585000   69.405000  151.585000   69.405000  149.850000 ;
      POLYGON   68.430000 -108.370000   68.430000 -111.820000   64.980000 -111.820000 ;
      POLYGON   68.430000 -102.150000   71.100000 -102.150000   68.430000 -104.820000 ;
      POLYGON   68.430000  -87.140000   68.430000  -98.545000   57.025000  -98.545000 ;
      POLYGON   69.365000 -142.790000   72.915000 -142.790000   69.365000 -146.340000 ;
      POLYGON   69.365000 -128.660000   69.365000 -132.170000   65.855000 -132.170000 ;
      POLYGON   69.365000 -123.375000   71.105000 -123.375000   69.365000 -125.115000 ;
      POLYGON   69.365000  146.340000   72.915000  142.790000   69.365000  142.790000 ;
      POLYGON   69.405000 -164.860000   72.075000 -164.860000   69.405000 -167.530000 ;
      POLYGON   69.405000 -149.850000   69.405000 -152.520000   66.735000 -152.520000 ;
      POLYGON   69.405000  149.850000   72.915000  149.850000   72.915000  146.340000 ;
      POLYGON   69.405000  167.530000   72.915000  164.020000   69.405000  164.020000 ;
      POLYGON   69.460000  103.790000   73.010000  100.240000   69.460000  100.240000 ;
      POLYGON   69.460000  107.340000   73.010000  107.340000   73.010000  103.790000 ;
      POLYGON   70.335000  124.145000   72.035000  122.445000   70.335000  122.445000 ;
      POLYGON   70.335000  127.690000   73.880000  127.690000   73.880000  124.145000 ;
      POLYGON   70.440000  170.040000   72.950000  170.040000   72.950000  167.530000 ;
      POLYGON   71.100000  -99.480000   73.770000  -99.480000   71.100000 -102.150000 ;
      POLYGON   71.105000 -119.830000   74.650000 -119.830000   71.105000 -123.375000 ;
      POLYGON   71.980000 -104.820000   71.980000 -108.370000   68.430000 -108.370000 ;
      POLYGON   72.035000  122.445000   75.580000  118.900000   72.035000  118.900000 ;
      POLYGON   72.075000 -161.315000   75.620000 -161.315000   72.075000 -164.860000 ;
      POLYGON   72.910000 -125.115000   72.910000 -128.660000   69.365000 -128.660000 ;
      POLYGON   72.915000 -146.340000   72.915000 -149.850000   69.405000 -149.850000 ;
      POLYGON   72.915000 -141.940000   73.765000 -141.940000   72.915000 -142.790000 ;
      POLYGON   72.915000  142.790000   75.580000  140.125000   72.915000  140.125000 ;
      POLYGON   72.915000  146.340000   76.465000  146.340000   76.465000  142.790000 ;
      POLYGON   72.915000  164.020000   75.585000  161.350000   72.915000  161.350000 ;
      POLYGON   72.950000 -167.530000   72.950000 -170.040000   70.440000 -170.040000 ;
      POLYGON   72.950000  167.530000   76.460000  167.530000   76.460000  164.020000 ;
      POLYGON   73.010000  100.240000   76.440000   96.810000   73.010000   96.810000 ;
      POLYGON   73.010000  103.790000   76.560000  103.790000   76.560000  100.240000 ;
      POLYGON   73.015000 -125.010000   73.015000 -125.115000   72.910000 -125.115000 ;
      POLYGON   73.765000 -138.390000   77.315000 -138.390000   73.765000 -141.940000 ;
      POLYGON   73.770000  -96.810000   76.440000  -96.810000   73.770000  -99.480000 ;
      POLYGON   73.880000  124.145000   75.580000  124.145000   75.580000  122.445000 ;
      POLYGON   74.650000 -123.375000   74.650000 -125.010000   73.015000 -125.010000 ;
      POLYGON   74.650000 -117.160000   77.320000 -117.160000   74.650000 -119.830000 ;
      POLYGON   74.650000 -102.150000   74.650000 -104.820000   71.980000 -104.820000 ;
      POLYGON   74.705000  -80.865000   74.705000  -87.140000   68.430000  -87.140000 ;
      POLYGON   75.580000  118.900000   78.255000  116.225000   75.580000  116.225000 ;
      POLYGON   75.580000  122.445000   79.125000  122.445000   79.125000  118.900000 ;
      POLYGON   75.580000  140.125000   78.250000  137.455000   75.580000  137.455000 ;
      POLYGON   75.585000  161.350000   79.130000  157.805000   75.585000  157.805000 ;
      POLYGON   75.620000 -167.530000   90.630000 -167.530000   75.620000 -182.540000 ;
      POLYGON   75.620000 -164.860000   75.620000 -167.530000   72.950000 -167.530000 ;
      POLYGON   75.620000 -157.770000   79.165000 -157.770000   75.620000 -161.315000 ;
      POLYGON   75.620000  182.540000   88.120000  170.040000   75.620000  170.040000 ;
      POLYGON   76.440000  -94.140000   79.110000  -94.140000   76.440000  -96.810000 ;
      POLYGON   76.440000   96.810000   79.950000   93.300000   76.440000   93.300000 ;
      POLYGON   76.460000  164.020000   79.130000  164.020000   79.130000  161.350000 ;
      POLYGON   76.465000 -142.790000   76.465000 -146.340000   72.915000 -146.340000 ;
      POLYGON   76.465000  142.790000   79.130000  142.790000   79.130000  140.125000 ;
      POLYGON   76.560000  100.240000   79.990000  100.240000   79.990000   96.810000 ;
      POLYGON   77.315000 -141.940000   77.315000 -142.790000   76.465000 -142.790000 ;
      POLYGON   77.315000 -134.840000   80.865000 -134.840000   77.315000 -138.390000 ;
      POLYGON   77.320000 -114.490000   79.990000 -114.490000   77.320000 -117.160000 ;
      POLYGON   77.320000  -99.480000   77.320000 -102.150000   74.650000 -102.150000 ;
      POLYGON   78.195000 -119.830000   78.195000 -123.375000   74.650000 -123.375000 ;
      POLYGON   78.250000  137.455000   81.800000  133.905000   78.250000  133.905000 ;
      POLYGON   78.255000  116.225000   80.925000  113.555000   78.255000  113.555000 ;
      POLYGON   79.110000  -90.690000   82.560000  -90.690000   79.110000  -94.140000 ;
      POLYGON   79.125000  118.900000   81.800000  118.900000   81.800000  116.225000 ;
      POLYGON   79.130000  140.125000   81.800000  140.125000   81.800000  137.455000 ;
      POLYGON   79.130000  157.805000   82.675000  154.260000   79.130000  154.260000 ;
      POLYGON   79.130000  161.350000   82.675000  161.350000   82.675000  157.805000 ;
      POLYGON   79.165000 -161.315000   79.165000 -164.860000   75.620000 -164.860000 ;
      POLYGON   79.165000 -156.940000   79.995000 -156.940000   79.165000 -157.770000 ;
      POLYGON   79.235000 -140.020000   79.235000 -141.940000   77.315000 -141.940000 ;
      POLYGON   79.950000   75.620000   80.920000   75.620000   80.920000   74.650000 ;
      POLYGON   79.950000   93.300000   80.920000   92.330000   79.950000   92.330000 ;
      POLYGON   79.990000 -110.980000   83.500000 -110.980000   79.990000 -114.490000 ;
      POLYGON   79.990000  -96.810000   79.990000  -99.480000   77.320000  -99.480000 ;
      POLYGON   79.990000   96.810000   83.500000   96.810000   83.500000   93.300000 ;
      POLYGON   79.995000 -153.395000   83.540000 -153.395000   79.995000 -156.940000 ;
      POLYGON   80.865000 -138.390000   80.865000 -140.020000   79.235000 -140.020000 ;
      POLYGON   80.865000 -132.170000   83.535000 -132.170000   80.865000 -134.840000 ;
      POLYGON   80.865000 -117.160000   80.865000 -119.830000   78.195000 -119.830000 ;
      POLYGON   80.920000   74.650000   97.565000   74.650000   97.565000   58.005000 ;
      POLYGON   80.920000   92.330000   83.590000   89.660000   80.920000   89.660000 ;
      POLYGON   80.925000  113.555000   84.470000  110.010000   80.925000  110.010000 ;
      POLYGON   81.800000  116.225000   84.470000  116.225000   84.470000  113.555000 ;
      POLYGON   81.800000  133.905000   85.350000  130.355000   81.800000  130.355000 ;
      POLYGON   81.800000  137.455000   85.350000  137.455000   85.350000  133.905000 ;
      POLYGON   82.560000  -87.140000   86.110000  -87.140000   82.560000  -90.690000 ;
      POLYGON   82.660000  -94.140000   82.660000  -96.810000   79.990000  -96.810000 ;
      POLYGON   82.675000  154.260000   86.220000  150.715000   82.675000  150.715000 ;
      POLYGON   82.675000  157.805000   86.220000  157.805000   86.220000  154.260000 ;
      POLYGON   82.710000 -157.770000   82.710000 -161.315000   79.165000 -161.315000 ;
      POLYGON   83.500000 -107.435000   87.045000 -107.435000   83.500000 -110.980000 ;
      POLYGON   83.500000   93.300000   84.470000   93.300000   84.470000   92.330000 ;
      POLYGON   83.535000 -128.660000   87.045000 -128.660000   83.535000 -132.170000 ;
      POLYGON   83.535000 -114.490000   83.535000 -117.160000   80.865000 -117.160000 ;
      POLYGON   83.540000 -156.940000   83.540000 -157.770000   82.710000 -157.770000 ;
      POLYGON   83.540000 -149.850000   87.085000 -149.850000   83.540000 -153.395000 ;
      POLYGON   83.590000   89.660000   87.140000   86.110000   83.590000   86.110000 ;
      POLYGON   84.415000 -134.840000   84.415000 -138.390000   80.865000 -138.390000 ;
      POLYGON   84.470000   92.330000   87.140000   92.330000   87.140000   89.660000 ;
      POLYGON   84.470000  110.010000   88.015000  106.465000   84.470000  106.465000 ;
      POLYGON   84.470000  113.555000   88.015000  113.555000   88.015000  110.010000 ;
      POLYGON   85.130000  -70.440000   85.130000  -80.865000   74.705000  -80.865000 ;
      POLYGON   85.350000  130.355000   87.045000  128.660000   85.350000  128.660000 ;
      POLYGON   85.350000  133.905000   88.900000  133.905000   88.900000  130.355000 ;
      POLYGON   86.110000  -90.690000   86.110000  -94.140000   82.660000  -94.140000 ;
      POLYGON   86.110000  -84.470000   88.780000  -84.470000   86.110000  -87.140000 ;
      POLYGON   86.220000  150.715000   89.755000  147.180000   86.220000  147.180000 ;
      POLYGON   86.220000  154.260000   89.765000  154.260000   89.765000  150.715000 ;
      POLYGON   87.045000 -125.110000   90.595000 -125.110000   87.045000 -128.660000 ;
      POLYGON   87.045000 -110.980000   87.045000 -114.490000   83.535000 -114.490000 ;
      POLYGON   87.045000 -105.695000   88.785000 -105.695000   87.045000 -107.435000 ;
      POLYGON   87.045000  128.660000   90.595000  125.110000   87.045000  125.110000 ;
      POLYGON   87.085000 -153.395000   87.085000 -156.940000   83.540000 -156.940000 ;
      POLYGON   87.085000 -147.180000   89.755000 -147.180000   87.085000 -149.850000 ;
      POLYGON   87.085000 -132.170000   87.085000 -134.840000   84.415000 -134.840000 ;
      POLYGON   87.140000   86.110000   90.690000   82.560000   87.140000   82.560000 ;
      POLYGON   87.140000   89.660000   90.690000   89.660000   90.690000   86.110000 ;
      POLYGON   88.015000  106.465000   89.715000  104.765000   88.015000  104.765000 ;
      POLYGON   88.015000  110.010000   91.560000  110.010000   91.560000  106.465000 ;
      POLYGON   88.120000  170.040000  100.355000  157.805000   88.120000  157.805000 ;
      POLYGON   88.780000  -81.800000   91.450000  -81.800000   88.780000  -84.470000 ;
      POLYGON   88.785000 -102.150000   92.330000 -102.150000   88.785000 -105.695000 ;
      POLYGON   88.900000  130.355000   90.595000  130.355000   90.595000  128.660000 ;
      POLYGON   89.660000  -87.140000   89.660000  -90.690000   86.110000  -90.690000 ;
      POLYGON   89.715000  104.765000   93.260000  101.220000   89.715000  101.220000 ;
      POLYGON   89.755000 -143.635000   93.300000 -143.635000   89.755000 -147.180000 ;
      POLYGON   89.755000  147.180000   93.265000  143.670000   89.755000  143.670000 ;
      POLYGON   89.765000  150.715000   93.300000  150.715000   93.300000  147.180000 ;
      POLYGON   90.590000 -107.435000   90.590000 -110.980000   87.045000 -110.980000 ;
      POLYGON   90.595000 -128.660000   90.595000 -132.170000   87.085000 -132.170000 ;
      POLYGON   90.595000 -124.260000   91.445000 -124.260000   90.595000 -125.110000 ;
      POLYGON   90.595000  125.110000   93.260000  122.445000   90.595000  122.445000 ;
      POLYGON   90.595000  128.660000   94.145000  128.660000   94.145000  125.110000 ;
      POLYGON   90.630000 -149.850000   90.630000 -153.395000   87.085000 -153.395000 ;
      POLYGON   90.630000 -149.850000  108.310000 -149.850000   90.630000 -167.530000 ;
      POLYGON   90.690000   82.560000   94.120000   79.130000   90.690000   79.130000 ;
      POLYGON   90.690000   86.110000   94.240000   86.110000   94.240000   82.560000 ;
      POLYGON   91.445000 -120.710000   94.995000 -120.710000   91.445000 -124.260000 ;
      POLYGON   91.450000  -79.130000   94.120000  -79.130000   91.450000  -81.800000 ;
      POLYGON   91.560000  106.465000   93.260000  106.465000   93.260000  104.765000 ;
      POLYGON   92.330000 -105.695000   92.330000 -107.435000   90.590000 -107.435000 ;
      POLYGON   92.330000  -99.480000   95.000000  -99.480000   92.330000 -102.150000 ;
      POLYGON   92.330000  -84.470000   92.330000  -87.140000   89.660000  -87.140000 ;
      POLYGON   92.385000  -63.185000   92.385000  -70.440000   85.130000  -70.440000 ;
      POLYGON   93.260000  101.220000   95.935000   98.545000   93.260000   98.545000 ;
      POLYGON   93.260000  104.765000   96.805000  104.765000   96.805000  101.220000 ;
      POLYGON   93.260000  122.445000   95.930000  119.775000   93.260000  119.775000 ;
      POLYGON   93.265000  143.670000   96.810000  140.125000   93.265000  140.125000 ;
      POLYGON   93.300000 -147.180000   93.300000 -149.850000   90.630000 -149.850000 ;
      POLYGON   93.300000 -140.090000   96.845000 -140.090000   93.300000 -143.635000 ;
      POLYGON   93.300000  147.180000   96.810000  147.180000   96.810000  143.670000 ;
      POLYGON   94.120000  -76.460000   96.790000  -76.460000   94.120000  -79.130000 ;
      POLYGON   94.120000   79.130000   97.630000   75.620000   94.120000   75.620000 ;
      POLYGON   94.145000 -125.110000   94.145000 -128.660000   90.595000 -128.660000 ;
      POLYGON   94.145000  125.110000   96.810000  125.110000   96.810000  122.445000 ;
      POLYGON   94.240000   82.560000   97.670000   82.560000   97.670000   79.130000 ;
      POLYGON   94.995000 -124.260000   94.995000 -125.110000   94.145000 -125.110000 ;
      POLYGON   94.995000 -117.160000   98.545000 -117.160000   94.995000 -120.710000 ;
      POLYGON   95.000000  -96.810000   97.670000  -96.810000   95.000000  -99.480000 ;
      POLYGON   95.000000  -81.800000   95.000000  -84.470000   92.330000  -84.470000 ;
      POLYGON   95.875000 -102.150000   95.875000 -105.695000   92.330000 -105.695000 ;
      POLYGON   95.930000  119.775000   99.480000  116.225000   95.930000  116.225000 ;
      POLYGON   95.935000   98.545000   98.605000   95.875000   95.935000   95.875000 ;
      POLYGON   96.790000  -73.010000  100.240000  -73.010000   96.790000  -76.460000 ;
      POLYGON   96.805000  101.220000   99.480000  101.220000   99.480000   98.545000 ;
      POLYGON   96.810000  122.445000   99.480000  122.445000   99.480000  119.775000 ;
      POLYGON   96.810000  140.125000  100.355000  136.580000   96.810000  136.580000 ;
      POLYGON   96.810000  143.670000  100.355000  143.670000  100.355000  140.125000 ;
      POLYGON   96.845000 -143.635000   96.845000 -147.180000   93.300000 -147.180000 ;
      POLYGON   96.845000 -139.260000   97.675000 -139.260000   96.845000 -140.090000 ;
      POLYGON   97.565000  -58.005000   97.565000  -63.185000   92.385000  -63.185000 ;
      POLYGON   97.565000   58.005000   98.600000   58.005000   98.600000   56.970000 ;
      POLYGON   97.630000   75.620000   98.600000   74.650000   97.630000   74.650000 ;
      POLYGON   97.670000  -93.300000  101.180000  -93.300000   97.670000  -96.810000 ;
      POLYGON   97.670000  -79.130000   97.670000  -81.800000   95.000000  -81.800000 ;
      POLYGON   97.670000   79.130000  101.180000   79.130000  101.180000   75.620000 ;
      POLYGON   97.675000 -135.715000  101.220000 -135.715000   97.675000 -139.260000 ;
      POLYGON   98.545000 -120.710000   98.545000 -124.260000   94.995000 -124.260000 ;
      POLYGON   98.545000 -114.490000  101.215000 -114.490000   98.545000 -117.160000 ;
      POLYGON   98.545000  -99.480000   98.545000 -102.150000   95.875000 -102.150000 ;
      POLYGON   98.600000   56.970000  110.000000   56.970000  110.000000   45.570000 ;
      POLYGON   98.600000   74.650000  101.270000   71.980000   98.600000   71.980000 ;
      POLYGON   98.605000   95.875000  102.150000   92.330000   98.605000   92.330000 ;
      POLYGON   99.480000   98.545000  102.150000   98.545000  102.150000   95.875000 ;
      POLYGON   99.480000  116.225000  103.030000  112.675000   99.480000  112.675000 ;
      POLYGON   99.480000  119.775000  103.030000  119.775000  103.030000  116.225000 ;
      POLYGON  100.240000  -69.460000  103.790000  -69.460000  100.240000  -73.010000 ;
      POLYGON  100.340000  -76.460000  100.340000  -79.130000   97.670000  -79.130000 ;
      POLYGON  100.355000  136.580000  103.900000  133.035000  100.355000  133.035000 ;
      POLYGON  100.355000  140.125000  103.900000  140.125000  103.900000  136.580000 ;
      POLYGON  100.355000  157.805000  118.035000  140.125000  100.355000  140.125000 ;
      POLYGON  100.390000 -140.090000  100.390000 -143.635000   96.845000 -143.635000 ;
      POLYGON  101.180000  -89.755000  104.725000  -89.755000  101.180000  -93.300000 ;
      POLYGON  101.180000   75.620000  102.150000   75.620000  102.150000   74.650000 ;
      POLYGON  101.215000 -110.980000  104.725000 -110.980000  101.215000 -114.490000 ;
      POLYGON  101.215000  -96.810000  101.215000  -99.480000   98.545000  -99.480000 ;
      POLYGON  101.220000 -139.260000  101.220000 -140.090000  100.390000 -140.090000 ;
      POLYGON  101.220000 -132.170000  104.765000 -132.170000  101.220000 -135.715000 ;
      POLYGON  101.270000   71.980000  104.820000   68.430000  101.270000   68.430000 ;
      POLYGON  102.095000 -117.160000  102.095000 -120.710000   98.545000 -120.710000 ;
      POLYGON  102.150000   74.650000  104.820000   74.650000  104.820000   71.980000 ;
      POLYGON  102.150000   92.330000  105.695000   88.785000  102.150000   88.785000 ;
      POLYGON  102.150000   95.875000  105.695000   95.875000  105.695000   92.330000 ;
      POLYGON  103.030000  112.675000  104.725000  110.980000  103.030000  110.980000 ;
      POLYGON  103.030000  116.225000  106.580000  116.225000  106.580000  112.675000 ;
      POLYGON  103.780000  -51.790000  103.780000  -58.005000   97.565000  -58.005000 ;
      POLYGON  103.790000  -73.010000  103.790000  -76.460000  100.340000  -76.460000 ;
      POLYGON  103.790000  -66.790000  106.460000  -66.790000  103.790000  -69.460000 ;
      POLYGON  103.900000  133.035000  107.435000  129.500000  103.900000  129.500000 ;
      POLYGON  103.900000  136.580000  107.445000  136.580000  107.445000  133.035000 ;
      POLYGON  104.725000 -107.430000  108.275000 -107.430000  104.725000 -110.980000 ;
      POLYGON  104.725000  -93.300000  104.725000  -96.810000  101.215000  -96.810000 ;
      POLYGON  104.725000  -88.015000  106.465000  -88.015000  104.725000  -89.755000 ;
      POLYGON  104.725000  110.980000  108.275000  107.430000  104.725000  107.430000 ;
      POLYGON  104.765000 -135.715000  104.765000 -139.260000  101.220000 -139.260000 ;
      POLYGON  104.765000 -129.500000  107.435000 -129.500000  104.765000 -132.170000 ;
      POLYGON  104.765000 -114.490000  104.765000 -117.160000  102.095000 -117.160000 ;
      POLYGON  104.820000   68.430000  108.370000   64.880000  104.820000   64.880000 ;
      POLYGON  104.820000   71.980000  108.370000   71.980000  108.370000   68.430000 ;
      POLYGON  105.695000   88.785000  107.395000   87.085000  105.695000   87.085000 ;
      POLYGON  105.695000   92.330000  109.240000   92.330000  109.240000   88.785000 ;
      POLYGON  106.360000  -70.440000  106.360000  -73.010000  103.790000  -73.010000 ;
      POLYGON  106.460000  -64.225000  109.025000  -64.225000  106.460000  -66.790000 ;
      POLYGON  106.465000  -84.470000  110.010000  -84.470000  106.465000  -88.015000 ;
      POLYGON  106.580000  112.675000  108.275000  112.675000  108.275000  110.980000 ;
      POLYGON  107.340000  -69.460000  107.340000  -70.440000  106.360000  -70.440000 ;
      POLYGON  107.395000   87.085000  110.940000   83.540000  107.395000   83.540000 ;
      POLYGON  107.435000 -125.955000  110.980000 -125.955000  107.435000 -129.500000 ;
      POLYGON  107.435000  129.500000  110.945000  125.990000  107.435000  125.990000 ;
      POLYGON  107.445000  133.035000  110.980000  133.035000  110.980000  129.500000 ;
      POLYGON  108.270000  -89.755000  108.270000  -93.300000  104.725000  -93.300000 ;
      POLYGON  108.275000 -110.980000  108.275000 -114.490000  104.765000 -114.490000 ;
      POLYGON  108.275000 -106.580000  109.125000 -106.580000  108.275000 -107.430000 ;
      POLYGON  108.275000  107.430000  110.940000  104.765000  108.275000  104.765000 ;
      POLYGON  108.275000  110.980000  111.825000  110.980000  111.825000  107.430000 ;
      POLYGON  108.310000 -132.170000  108.310000 -135.715000  104.765000 -135.715000 ;
      POLYGON  108.310000 -132.170000  125.990000 -132.170000  108.310000 -149.850000 ;
      POLYGON  108.370000   64.880000  110.065000   63.185000  108.370000   63.185000 ;
      POLYGON  108.370000   68.430000  111.920000   68.430000  111.920000   64.880000 ;
      POLYGON  109.025000  -63.185000  110.065000  -63.185000  109.025000  -64.225000 ;
      POLYGON  109.125000 -103.030000  112.675000 -103.030000  109.125000 -106.580000 ;
      POLYGON  109.240000   88.785000  110.940000   88.785000  110.940000   87.085000 ;
      POLYGON  110.000000  -45.570000  110.000000  -51.790000  103.780000  -51.790000 ;
      POLYGON  110.010000  -88.015000  110.010000  -89.755000  108.270000  -89.755000 ;
      POLYGON  110.010000  -81.800000  112.680000  -81.800000  110.010000  -84.470000 ;
      POLYGON  110.010000  -66.790000  110.010000  -69.460000  107.340000  -69.460000 ;
      POLYGON  110.065000  -59.635000  113.615000  -59.635000  110.065000  -63.185000 ;
      POLYGON  110.065000   63.185000  113.615000   59.635000  110.065000   59.635000 ;
      POLYGON  110.940000   83.540000  113.615000   80.865000  110.940000   80.865000 ;
      POLYGON  110.940000   87.085000  114.485000   87.085000  114.485000   83.540000 ;
      POLYGON  110.940000  104.765000  113.610000  102.095000  110.940000  102.095000 ;
      POLYGON  110.945000  125.990000  114.490000  122.445000  110.945000  122.445000 ;
      POLYGON  110.980000 -129.500000  110.980000 -132.170000  108.310000 -132.170000 ;
      POLYGON  110.980000 -122.410000  114.525000 -122.410000  110.980000 -125.955000 ;
      POLYGON  110.980000  129.500000  114.490000  129.500000  114.490000  125.990000 ;
      POLYGON  111.825000 -107.430000  111.825000 -110.980000  108.275000 -110.980000 ;
      POLYGON  111.825000  107.430000  114.490000  107.430000  114.490000  104.765000 ;
      POLYGON  111.920000   64.880000  113.615000   64.880000  113.615000   63.185000 ;
      POLYGON  112.575000  -64.225000  112.575000  -66.790000  110.010000  -66.790000 ;
      POLYGON  112.675000 -106.580000  112.675000 -107.430000  111.825000 -107.430000 ;
      POLYGON  112.675000  -99.480000  116.225000  -99.480000  112.675000 -103.030000 ;
      POLYGON  112.680000  -79.130000  115.350000  -79.130000  112.680000  -81.800000 ;
      POLYGON  113.555000  -84.470000  113.555000  -88.015000  110.010000  -88.015000 ;
      POLYGON  113.610000  102.095000  117.160000   98.545000  113.610000   98.545000 ;
      POLYGON  113.615000  -63.185000  113.615000  -64.225000  112.575000  -64.225000 ;
      POLYGON  113.615000  -58.005000  115.245000  -58.005000  113.615000  -59.635000 ;
      POLYGON  113.615000   59.635000  116.280000   56.970000  113.615000   56.970000 ;
      POLYGON  113.615000   63.185000  117.165000   63.185000  117.165000   59.635000 ;
      POLYGON  113.615000   80.865000  116.285000   78.195000  113.615000   78.195000 ;
      POLYGON  114.485000   83.540000  117.160000   83.540000  117.160000   80.865000 ;
      POLYGON  114.490000  104.765000  117.160000  104.765000  117.160000  102.095000 ;
      POLYGON  114.490000  122.445000  118.035000  118.900000  114.490000  118.900000 ;
      POLYGON  114.490000  125.990000  118.035000  125.990000  118.035000  122.445000 ;
      POLYGON  114.525000 -125.955000  114.525000 -129.500000  110.980000 -129.500000 ;
      POLYGON  114.525000 -121.580000  115.355000 -121.580000  114.525000 -122.410000 ;
      POLYGON  115.245000  -55.330000  117.920000  -55.330000  115.245000  -58.005000 ;
      POLYGON  115.350000  -75.620000  118.860000  -75.620000  115.350000  -79.130000 ;
      POLYGON  115.355000 -118.035000  118.900000 -118.035000  115.355000 -121.580000 ;
      POLYGON  116.225000 -103.030000  116.225000 -106.580000  112.675000 -106.580000 ;
      POLYGON  116.225000  -96.810000  118.895000  -96.810000  116.225000  -99.480000 ;
      POLYGON  116.225000  -81.800000  116.225000  -84.470000  113.555000  -84.470000 ;
      POLYGON  116.280000   56.970000  118.950000   54.300000  116.280000   54.300000 ;
      POLYGON  116.285000   78.195000  119.830000   74.650000  116.285000   74.650000 ;
      POLYGON  117.160000   80.865000  119.830000   80.865000  119.830000   78.195000 ;
      POLYGON  117.160000   98.545000  120.710000   94.995000  117.160000   94.995000 ;
      POLYGON  117.160000  102.095000  120.710000  102.095000  120.710000   98.545000 ;
      POLYGON  117.165000  -59.635000  117.165000  -63.185000  113.615000  -63.185000 ;
      POLYGON  117.165000   59.635000  119.830000   59.635000  119.830000   56.970000 ;
      POLYGON  117.920000  -51.790000  121.460000  -51.790000  117.920000  -55.330000 ;
      POLYGON  118.035000  118.900000  121.580000  115.355000  118.035000  115.355000 ;
      POLYGON  118.035000  122.445000  121.580000  122.445000  121.580000  118.900000 ;
      POLYGON  118.035000  140.125000  135.715000  122.445000  118.035000  122.445000 ;
      POLYGON  118.070000 -122.410000  118.070000 -125.955000  114.525000 -125.955000 ;
      POLYGON  118.795000  -58.005000  118.795000  -59.635000  117.165000  -59.635000 ;
      POLYGON  118.860000  -72.075000  122.405000  -72.075000  118.860000  -75.620000 ;
      POLYGON  118.895000  -93.300000  122.405000  -93.300000  118.895000  -96.810000 ;
      POLYGON  118.895000  -79.130000  118.895000  -81.800000  116.225000  -81.800000 ;
      POLYGON  118.900000 -121.580000  118.900000 -122.410000  118.070000 -122.410000 ;
      POLYGON  118.900000 -114.490000  122.445000 -114.490000  118.900000 -118.035000 ;
      POLYGON  118.950000   54.300000  122.500000   50.750000  118.950000   50.750000 ;
      POLYGON  119.775000  -99.480000  119.775000 -103.030000  116.225000 -103.030000 ;
      POLYGON  119.830000   56.970000  122.500000   56.970000  122.500000   54.300000 ;
      POLYGON  119.830000   74.650000  123.375000   71.105000  119.830000   71.105000 ;
      POLYGON  119.830000   78.195000  123.375000   78.195000  123.375000   74.650000 ;
      POLYGON  120.710000   94.995000  122.405000   93.300000  120.710000   93.300000 ;
      POLYGON  120.710000   98.545000  124.260000   98.545000  124.260000   94.995000 ;
      POLYGON  121.460000  -50.750000  122.500000  -50.750000  121.460000  -51.790000 ;
      POLYGON  121.470000  -55.330000  121.470000  -58.005000  118.795000  -58.005000 ;
      POLYGON  121.580000  115.355000  125.115000  111.820000  121.580000  111.820000 ;
      POLYGON  121.580000  118.900000  125.125000  118.900000  125.125000  115.355000 ;
      POLYGON  122.405000  -89.750000  125.955000  -89.750000  122.405000  -93.300000 ;
      POLYGON  122.405000  -75.620000  122.405000  -79.130000  118.895000  -79.130000 ;
      POLYGON  122.405000  -70.335000  124.145000  -70.335000  122.405000  -72.075000 ;
      POLYGON  122.405000   93.300000  125.955000   89.750000  122.405000   89.750000 ;
      POLYGON  122.445000 -118.035000  122.445000 -121.580000  118.900000 -121.580000 ;
      POLYGON  122.445000 -111.820000  125.115000 -111.820000  122.445000 -114.490000 ;
      POLYGON  122.445000  -96.810000  122.445000  -99.480000  119.775000  -99.480000 ;
      POLYGON  122.500000   54.300000  125.010000   54.300000  125.010000   51.790000 ;
      POLYGON  123.375000   71.105000  125.075000   69.405000  123.375000   69.405000 ;
      POLYGON  123.375000   74.650000  126.920000   74.650000  126.920000   71.105000 ;
      POLYGON  124.145000  -66.790000  127.690000  -66.790000  124.145000  -70.335000 ;
      POLYGON  124.260000   94.995000  125.955000   94.995000  125.955000   93.300000 ;
      POLYGON  125.010000  -51.790000  125.010000  -55.330000  121.470000  -55.330000 ;
      POLYGON  125.075000   69.405000  128.620000   65.860000  125.075000   65.860000 ;
      POLYGON  125.115000 -108.275000  128.660000 -108.275000  125.115000 -111.820000 ;
      POLYGON  125.115000  111.820000  128.625000  108.310000  125.115000  108.310000 ;
      POLYGON  125.125000  115.355000  128.660000  115.355000  128.660000  111.820000 ;
      POLYGON  125.950000  -72.075000  125.950000  -75.620000  122.405000  -75.620000 ;
      POLYGON  125.955000  -93.300000  125.955000  -96.810000  122.445000  -96.810000 ;
      POLYGON  125.955000  -88.900000  126.805000  -88.900000  125.955000  -89.750000 ;
      POLYGON  125.955000   89.750000  128.620000   87.085000  125.955000   87.085000 ;
      POLYGON  125.955000   93.300000  129.505000   93.300000  129.505000   89.750000 ;
      POLYGON  125.990000 -114.490000  125.990000 -118.035000  122.445000 -118.035000 ;
      POLYGON  125.990000 -114.490000  143.670000 -114.490000  125.990000 -132.170000 ;
      POLYGON  126.805000  -85.350000  130.355000  -85.350000  126.805000  -88.900000 ;
      POLYGON  126.920000   71.105000  128.620000   71.105000  128.620000   69.405000 ;
      POLYGON  127.585000  -70.440000  127.585000  -72.075000  125.950000  -72.075000 ;
      POLYGON  127.690000  -70.335000  127.690000  -70.440000  127.585000  -70.440000 ;
      POLYGON  127.690000  -64.225000  130.255000  -64.225000  127.690000  -66.790000 ;
      POLYGON  128.620000   65.860000  131.295000   63.185000  128.620000   63.185000 ;
      POLYGON  128.620000   69.405000  132.165000   69.405000  132.165000   65.860000 ;
      POLYGON  128.620000   87.085000  131.290000   84.415000  128.620000   84.415000 ;
      POLYGON  128.625000  108.310000  132.170000  104.765000  128.625000  104.765000 ;
      POLYGON  128.660000 -111.820000  128.660000 -114.490000  125.990000 -114.490000 ;
      POLYGON  128.660000 -104.730000  132.205000 -104.730000  128.660000 -108.275000 ;
      POLYGON  128.660000  111.820000  132.170000  111.820000  132.170000  108.310000 ;
      POLYGON  129.505000  -89.750000  129.505000  -93.300000  125.955000  -93.300000 ;
      POLYGON  129.505000   89.750000  132.170000   89.750000  132.170000   87.085000 ;
      POLYGON  130.255000  -63.185000  131.295000  -63.185000  130.255000  -64.225000 ;
      POLYGON  130.355000  -88.900000  130.355000  -89.750000  129.505000  -89.750000 ;
      POLYGON  130.355000  -81.800000  133.905000  -81.800000  130.355000  -85.350000 ;
      POLYGON  131.235000  -66.790000  131.235000  -70.335000  127.690000  -70.335000 ;
      POLYGON  131.290000   84.415000  134.840000   80.865000  131.290000   80.865000 ;
      POLYGON  131.295000  -60.515000  133.965000  -60.515000  131.295000  -63.185000 ;
      POLYGON  131.295000   63.185000  133.965000   60.515000  131.295000   60.515000 ;
      POLYGON  132.165000   65.860000  134.840000   65.860000  134.840000   63.185000 ;
      POLYGON  132.170000   87.085000  134.840000   87.085000  134.840000   84.415000 ;
      POLYGON  132.170000  104.765000  135.715000  101.220000  132.170000  101.220000 ;
      POLYGON  132.170000  108.310000  135.715000  108.310000  135.715000  104.765000 ;
      POLYGON  132.205000 -108.275000  132.205000 -111.820000  128.660000 -111.820000 ;
      POLYGON  132.205000 -103.900000  133.035000 -103.900000  132.205000 -104.730000 ;
      POLYGON  133.035000 -100.355000  136.580000 -100.355000  133.035000 -103.900000 ;
      POLYGON  133.800000  -64.225000  133.800000  -66.790000  131.235000  -66.790000 ;
      POLYGON  133.905000  -85.350000  133.905000  -88.900000  130.355000  -88.900000 ;
      POLYGON  133.905000  -79.130000  136.575000  -79.130000  133.905000  -81.800000 ;
      POLYGON  133.965000  -56.970000  137.510000  -56.970000  133.965000  -60.515000 ;
      POLYGON  133.965000   60.515000  137.510000   56.970000  133.965000   56.970000 ;
      POLYGON  134.840000  -63.185000  134.840000  -64.225000  133.800000  -64.225000 ;
      POLYGON  134.840000   63.185000  137.510000   63.185000  137.510000   60.515000 ;
      POLYGON  134.840000   80.865000  138.390000   77.315000  134.840000   77.315000 ;
      POLYGON  134.840000   84.415000  138.390000   84.415000  138.390000   80.865000 ;
      POLYGON  135.715000  101.220000  139.260000   97.675000  135.715000   97.675000 ;
      POLYGON  135.715000  104.765000  139.260000  104.765000  139.260000  101.220000 ;
      POLYGON  135.715000  122.445000  153.395000  104.765000  135.715000  104.765000 ;
      POLYGON  135.750000 -104.730000  135.750000 -108.275000  132.205000 -108.275000 ;
      POLYGON  136.575000  -75.620000  140.085000  -75.620000  136.575000  -79.130000 ;
      POLYGON  136.580000 -103.900000  136.580000 -104.730000  135.750000 -104.730000 ;
      POLYGON  136.580000  -96.810000  140.125000  -96.810000  136.580000 -100.355000 ;
      POLYGON  137.455000  -81.800000  137.455000  -85.350000  133.905000  -85.350000 ;
      POLYGON  137.510000  -60.515000  137.510000  -63.185000  134.840000  -63.185000 ;
      POLYGON  137.510000   60.515000  140.020000   60.515000  140.020000   58.005000 ;
      POLYGON  138.390000   77.315000  140.085000   75.620000  138.390000   75.620000 ;
      POLYGON  138.390000   80.865000  141.940000   80.865000  141.940000   77.315000 ;
      POLYGON  139.260000   97.675000  142.795000   94.140000  139.260000   94.140000 ;
      POLYGON  139.260000  101.220000  142.805000  101.220000  142.805000   97.675000 ;
      POLYGON  140.020000  -58.005000  140.020000  -60.515000  137.510000  -60.515000 ;
      POLYGON  140.085000  -72.070000  143.635000  -72.070000  140.085000  -75.620000 ;
      POLYGON  140.085000   75.620000  143.635000   72.070000  140.085000   72.070000 ;
      POLYGON  140.125000 -100.355000  140.125000 -103.900000  136.580000 -103.900000 ;
      POLYGON  140.125000  -94.140000  142.795000  -94.140000  140.125000  -96.810000 ;
      POLYGON  140.125000  -79.130000  140.125000  -81.800000  137.455000  -81.800000 ;
      POLYGON  141.940000   77.315000  143.635000   77.315000  143.635000   75.620000 ;
      POLYGON  142.795000  -90.595000  146.340000  -90.595000  142.795000  -94.140000 ;
      POLYGON  142.795000   94.140000  146.305000   90.630000  142.795000   90.630000 ;
      POLYGON  142.805000   97.675000  146.340000   97.675000  146.340000   94.140000 ;
      POLYGON  143.635000  -75.620000  143.635000  -79.130000  140.125000  -79.130000 ;
      POLYGON  143.635000  -70.440000  145.265000  -70.440000  143.635000  -72.070000 ;
      POLYGON  143.635000   72.070000  146.300000   69.405000  143.635000   69.405000 ;
      POLYGON  143.635000   75.620000  147.185000   75.620000  147.185000   72.070000 ;
      POLYGON  143.670000  -96.810000  143.670000 -100.355000  140.125000 -100.355000 ;
      POLYGON  143.670000  -96.810000  161.350000  -96.810000  143.670000 -114.490000 ;
      POLYGON  145.265000  -67.670000  148.035000  -67.670000  145.265000  -70.440000 ;
      POLYGON  146.300000   69.405000  148.970000   66.735000  146.300000   66.735000 ;
      POLYGON  146.305000   90.630000  149.850000   87.085000  146.305000   87.085000 ;
      POLYGON  146.340000  -94.140000  146.340000  -96.810000  143.670000  -96.810000 ;
      POLYGON  146.340000  -87.050000  149.885000  -87.050000  146.340000  -90.595000 ;
      POLYGON  146.340000   94.140000  149.850000   94.140000  149.850000   90.630000 ;
      POLYGON  147.185000  -72.070000  147.185000  -75.620000  143.635000  -75.620000 ;
      POLYGON  147.185000   72.070000  149.850000   72.070000  149.850000   69.405000 ;
      POLYGON  148.035000  -64.225000  151.480000  -64.225000  148.035000  -67.670000 ;
      POLYGON  148.815000  -70.440000  148.815000  -72.070000  147.185000  -72.070000 ;
      POLYGON  148.970000   66.735000  152.520000   63.185000  148.970000   63.185000 ;
      POLYGON  149.850000   69.405000  152.520000   69.405000  152.520000   66.735000 ;
      POLYGON  149.850000   87.085000  153.395000   83.540000  149.850000   83.540000 ;
      POLYGON  149.850000   90.630000  153.395000   90.630000  153.395000   87.085000 ;
      POLYGON  149.885000  -90.595000  149.885000  -94.140000  146.340000  -94.140000 ;
      POLYGON  149.885000  -86.220000  150.715000  -86.220000  149.885000  -87.050000 ;
      POLYGON  150.715000  -82.675000  154.260000  -82.675000  150.715000  -86.220000 ;
      POLYGON  151.480000  -63.185000  152.520000  -63.185000  151.480000  -64.225000 ;
      POLYGON  151.585000  -67.670000  151.585000  -70.440000  148.815000  -70.440000 ;
      POLYGON  152.520000   66.735000  155.030000   66.735000  155.030000   64.225000 ;
      POLYGON  153.395000   83.540000  156.940000   79.995000  153.395000   79.995000 ;
      POLYGON  153.395000   87.085000  156.940000   87.085000  156.940000   83.540000 ;
      POLYGON  153.395000  104.765000  171.075000   87.085000  153.395000   87.085000 ;
      POLYGON  153.430000  -87.050000  153.430000  -90.595000  149.885000  -90.595000 ;
      POLYGON  154.260000  -86.220000  154.260000  -87.050000  153.430000  -87.050000 ;
      POLYGON  154.260000  -79.130000  157.805000  -79.130000  154.260000  -82.675000 ;
      POLYGON  155.030000  -64.225000  155.030000  -67.670000  151.585000  -67.670000 ;
      POLYGON  156.940000   79.995000  160.475000   76.460000  156.940000   76.460000 ;
      POLYGON  156.940000   83.540000  160.485000   83.540000  160.485000   79.995000 ;
      POLYGON  157.805000  -82.675000  157.805000  -86.220000  154.260000  -86.220000 ;
      POLYGON  157.805000  -76.460000  160.475000  -76.460000  157.805000  -79.130000 ;
      POLYGON  160.475000  -72.950000  163.985000  -72.950000  160.475000  -76.460000 ;
      POLYGON  160.475000   76.460000  163.985000   72.950000  160.475000   72.950000 ;
      POLYGON  160.485000   79.995000  164.020000   79.995000  164.020000   76.460000 ;
      POLYGON  161.350000  -79.130000  161.350000  -82.675000  157.805000  -82.675000 ;
      POLYGON  161.350000  -79.130000  179.030000  -79.130000  161.350000  -96.810000 ;
      POLYGON  163.985000  -69.405000  167.530000  -69.405000  163.985000  -72.950000 ;
      POLYGON  163.985000   72.950000  167.530000   69.405000  163.985000   69.405000 ;
      POLYGON  164.020000  -76.460000  164.020000  -79.130000  161.350000  -79.130000 ;
      POLYGON  164.020000   76.460000  167.530000   76.460000  167.530000   72.950000 ;
      POLYGON  167.530000  -72.950000  167.530000  -76.460000  164.020000  -76.460000 ;
      POLYGON  167.530000   72.950000  170.040000   72.950000  170.040000   70.440000 ;
      POLYGON  170.040000  -70.440000  170.040000  -72.950000  167.530000  -72.950000 ;
      POLYGON  171.075000   87.085000  182.540000   75.620000  171.075000   75.620000 ;
      POLYGON  179.030000  -75.620000  182.540000  -75.620000  179.030000  -79.130000 ;
      RECT -182.540000  -75.620000 -167.530000  -72.950000 ;
      RECT -182.540000  -72.950000 -170.040000   72.950000 ;
      RECT -182.540000   72.950000 -167.530000   75.620000 ;
      RECT -171.075000  -87.085000 -156.940000  -83.540000 ;
      RECT -171.075000  -83.540000 -160.475000  -80.005000 ;
      RECT -171.075000  -80.005000 -164.020000  -76.460000 ;
      RECT -171.075000  -76.460000 -167.530000  -75.620000 ;
      RECT -167.530000  -69.405000 -152.520000  -66.735000 ;
      RECT -167.530000  -66.735000 -155.030000   67.670000 ;
      RECT -167.530000   67.670000 -151.585000   69.405000 ;
      RECT -166.495000  -70.440000 -149.850000  -69.405000 ;
      RECT -166.495000   69.405000 -149.850000   70.440000 ;
      RECT -164.860000   79.130000 -161.350000   82.675000 ;
      RECT -164.860000   82.675000 -157.805000   86.220000 ;
      RECT -164.860000   86.220000 -154.260000   89.755000 ;
      RECT -164.860000   89.755000 -150.725000   93.300000 ;
      RECT -163.985000  -72.950000 -147.185000  -72.070000 ;
      RECT -163.985000  -72.070000 -149.850000  -70.440000 ;
      RECT -163.985000   70.440000 -149.850000   72.070000 ;
      RECT -163.985000   72.070000 -147.185000   72.950000 ;
      RECT -161.315000   72.950000 -147.185000   75.620000 ;
      RECT -160.475000  -76.460000 -143.635000  -75.620000 ;
      RECT -160.475000  -75.620000 -147.185000  -72.950000 ;
      RECT -157.805000   75.620000 -143.635000   79.130000 ;
      RECT -156.930000  -80.005000 -140.125000  -79.130000 ;
      RECT -156.930000  -79.130000 -143.635000  -76.460000 ;
      RECT -154.260000   79.130000 -140.125000   81.800000 ;
      RECT -154.260000   81.800000 -137.455000   82.675000 ;
      RECT -153.395000 -104.765000 -139.260000 -101.220000 ;
      RECT -153.395000 -101.220000 -142.795000  -97.685000 ;
      RECT -153.395000  -97.685000 -146.340000  -94.140000 ;
      RECT -153.395000  -94.140000 -149.850000  -90.630000 ;
      RECT -153.395000  -83.540000 -138.390000  -80.865000 ;
      RECT -153.395000  -80.865000 -140.125000  -80.005000 ;
      RECT -152.520000  -63.185000 -137.510000  -60.515000 ;
      RECT -152.520000  -60.515000 -140.020000   60.515000 ;
      RECT -152.520000   60.515000 -137.510000   63.185000 ;
      RECT -151.585000   63.185000 -134.840000   64.120000 ;
      RECT -151.480000  -64.225000 -134.840000  -63.185000 ;
      RECT -151.480000   64.120000 -133.905000   64.225000 ;
      RECT -150.715000   82.675000 -137.455000   85.350000 ;
      RECT -150.715000   85.350000 -133.905000   86.220000 ;
      RECT -149.850000  -87.085000 -134.840000  -84.415000 ;
      RECT -149.850000  -84.415000 -138.390000  -83.540000 ;
      RECT -148.970000  -66.735000 -132.165000  -65.860000 ;
      RECT -148.970000  -65.860000 -134.840000  -64.225000 ;
      RECT -148.035000   64.225000 -133.905000   66.790000 ;
      RECT -148.035000   66.790000 -131.235000   67.670000 ;
      RECT -147.180000   86.220000 -133.905000   87.085000 ;
      RECT -147.180000   87.085000 -132.170000   89.750000 ;
      RECT -147.180000   89.750000 -129.505000   89.755000 ;
      RECT -147.180000   96.810000 -143.670000  100.355000 ;
      RECT -147.180000  100.355000 -140.125000  103.900000 ;
      RECT -147.180000  103.900000 -136.580000  107.435000 ;
      RECT -147.180000  107.435000 -133.045000  110.980000 ;
      RECT -146.305000  -90.630000 -129.505000  -89.750000 ;
      RECT -146.305000  -89.750000 -132.170000  -87.085000 ;
      RECT -146.300000  -69.405000 -132.165000  -66.735000 ;
      RECT -146.300000   67.670000 -131.235000   69.405000 ;
      RECT -145.265000   69.405000 -128.620000   70.440000 ;
      RECT -143.635000  -72.070000 -126.920000  -71.105000 ;
      RECT -143.635000  -71.105000 -128.620000  -69.405000 ;
      RECT -143.635000   70.440000 -128.620000   72.070000 ;
      RECT -143.635000   89.755000 -129.505000   93.300000 ;
      RECT -142.795000  -94.140000 -125.955000  -93.300000 ;
      RECT -142.795000  -93.300000 -129.505000  -90.630000 ;
      RECT -140.125000   93.300000 -125.955000   96.810000 ;
      RECT -140.085000  -75.620000 -123.375000  -74.650000 ;
      RECT -140.085000  -74.650000 -126.920000  -72.070000 ;
      RECT -140.085000   72.070000 -128.620000   72.075000 ;
      RECT -140.085000   72.075000 -125.950000   75.620000 ;
      RECT -139.735000  110.980000 -129.500000  114.490000 ;
      RECT -139.735000  114.490000 -125.990000  118.035000 ;
      RECT -139.735000  118.035000 -122.445000  118.425000 ;
      RECT -139.250000  -97.685000 -122.445000  -96.810000 ;
      RECT -139.250000  -96.810000 -125.955000  -94.140000 ;
      RECT -137.510000  -56.970000 -122.500000  -54.300000 ;
      RECT -137.510000  -54.300000 -125.010000   55.330000 ;
      RECT -137.510000   55.330000 -121.470000   56.970000 ;
      RECT -136.580000   96.810000 -122.445000   99.480000 ;
      RECT -136.580000   99.480000 -119.775000  100.355000 ;
      RECT -136.575000  -79.130000 -119.830000  -78.195000 ;
      RECT -136.575000  -78.195000 -123.375000  -75.620000 ;
      RECT -136.575000   75.620000 -122.405000   79.130000 ;
      RECT -136.475000  -58.005000 -119.830000  -56.970000 ;
      RECT -136.475000   56.970000 -119.830000   58.005000 ;
      RECT -135.715000 -122.445000 -121.580000 -118.900000 ;
      RECT -135.715000 -118.900000 -125.115000 -115.365000 ;
      RECT -135.715000 -115.365000 -128.660000 -111.820000 ;
      RECT -135.715000 -111.820000 -132.170000 -108.310000 ;
      RECT -135.715000 -101.220000 -120.710000  -98.545000 ;
      RECT -135.715000  -98.545000 -122.445000  -97.685000 ;
      RECT -134.840000  -80.865000 -119.830000  -79.130000 ;
      RECT -133.965000  -60.515000 -117.165000  -59.635000 ;
      RECT -133.965000  -59.635000 -119.830000  -58.005000 ;
      RECT -133.965000   58.005000 -119.830000   59.635000 ;
      RECT -133.965000   59.635000 -117.165000   60.515000 ;
      RECT -133.905000   79.130000 -118.895000   81.800000 ;
      RECT -133.035000  100.355000 -119.775000  103.030000 ;
      RECT -133.035000  103.030000 -116.225000  103.900000 ;
      RECT -132.170000 -104.765000 -117.160000 -102.095000 ;
      RECT -132.170000 -102.095000 -120.710000 -101.220000 ;
      RECT -131.545000  118.425000 -122.445000  121.580000 ;
      RECT -131.545000  121.580000 -118.900000  125.115000 ;
      RECT -131.545000  125.115000 -115.365000  126.615000 ;
      RECT -131.295000  -63.185000 -117.165000  -60.515000 ;
      RECT -131.295000   60.515000 -117.165000   63.185000 ;
      RECT -131.290000  -84.415000 -114.485000  -83.540000 ;
      RECT -131.290000  -83.540000 -117.160000  -80.865000 ;
      RECT -130.360000   63.185000 -113.615000   64.120000 ;
      RECT -130.355000   81.800000 -116.225000   84.470000 ;
      RECT -130.355000   84.470000 -113.555000   85.350000 ;
      RECT -129.500000  103.900000 -116.225000  104.765000 ;
      RECT -129.500000  104.765000 -114.490000  107.430000 ;
      RECT -129.500000  107.430000 -111.825000  107.435000 ;
      RECT -128.625000 -108.310000 -111.825000 -107.430000 ;
      RECT -128.625000 -107.430000 -114.490000 -104.765000 ;
      RECT -128.620000  -87.085000 -114.485000  -84.415000 ;
      RECT -128.620000  -65.860000 -112.575000  -64.225000 ;
      RECT -128.620000  -64.225000 -113.615000  -63.185000 ;
      RECT -128.620000   85.350000 -113.555000   87.085000 ;
      RECT -127.690000   64.120000 -112.680000   66.790000 ;
      RECT -125.955000  -89.750000 -109.240000  -88.785000 ;
      RECT -125.955000  -88.785000 -110.940000  -87.085000 ;
      RECT -125.955000   87.085000 -110.940000   89.750000 ;
      RECT -125.955000  107.435000 -111.825000  110.980000 ;
      RECT -125.115000 -111.820000 -108.275000 -110.980000 ;
      RECT -125.115000 -110.980000 -111.825000 -108.310000 ;
      RECT -125.075000  -69.405000 -110.010000  -66.790000 ;
      RECT -125.075000  -66.790000 -112.575000  -65.860000 ;
      RECT -125.075000   66.790000 -110.010000   69.405000 ;
      RECT -124.145000   69.405000 -110.010000   69.460000 ;
      RECT -124.145000   69.460000 -107.340000   70.335000 ;
      RECT -123.375000  -71.105000 -107.395000  -69.405000 ;
      RECT -122.500000  -50.750000 -110.000000   -6.250000 ;
      RECT -122.500000   -6.250000  105.000000    6.250000 ;
      RECT -122.500000    6.250000 -110.000000   50.750000 ;
      RECT -122.445000  110.980000 -108.275000  112.885000 ;
      RECT -122.445000  112.885000 -106.370000  114.490000 ;
      RECT -122.405000  -93.300000 -105.695000  -92.330000 ;
      RECT -122.405000  -92.330000 -109.240000  -89.750000 ;
      RECT -122.405000   70.335000 -107.340000   72.075000 ;
      RECT -122.405000   89.750000 -110.940000   89.755000 ;
      RECT -122.405000   89.755000 -108.270000   93.300000 ;
      RECT -122.255000  126.615000 -115.365000  128.660000 ;
      RECT -122.255000  128.660000 -111.820000  132.170000 ;
      RECT -122.255000  132.170000 -108.310000  135.715000 ;
      RECT -122.255000  135.715000 -104.765000  135.905000 ;
      RECT -121.570000 -115.365000 -104.765000 -114.490000 ;
      RECT -121.570000 -114.490000 -108.275000 -111.820000 ;
      RECT -121.470000   50.750000 -110.000000   51.780000 ;
      RECT -121.460000  -51.790000 -110.000000  -50.750000 ;
      RECT -121.460000   51.780000 -110.000000   51.790000 ;
      RECT -119.830000  -74.650000 -104.820000  -71.980000 ;
      RECT -119.830000  -71.980000 -107.395000  -71.105000 ;
      RECT -119.830000   72.075000 -107.340000   73.010000 ;
      RECT -119.830000   73.010000 -103.790000   74.650000 ;
      RECT -118.950000  -54.300000 -110.000000  -51.790000 ;
      RECT -118.900000  114.490000 -106.370000  116.225000 ;
      RECT -118.900000  116.225000 -103.030000  118.035000 ;
      RECT -118.895000  -96.810000 -102.150000  -95.875000 ;
      RECT -118.895000  -95.875000 -105.695000  -93.300000 ;
      RECT -118.895000   93.300000 -104.725000   96.810000 ;
      RECT -118.860000   74.650000 -103.790000   75.620000 ;
      RECT -118.035000 -140.125000 -103.900000 -136.580000 ;
      RECT -118.035000 -136.580000 -107.435000 -133.045000 ;
      RECT -118.035000 -133.045000 -110.980000 -129.500000 ;
      RECT -118.035000 -129.500000 -114.490000 -125.990000 ;
      RECT -118.035000 -118.900000 -103.030000 -116.225000 ;
      RECT -118.035000 -116.225000 -104.765000 -115.365000 ;
      RECT -117.920000   51.790000 -110.000000   55.330000 ;
      RECT -117.160000  -98.545000 -102.150000  -96.810000 ;
      RECT -116.535000  135.905000 -104.765000  139.260000 ;
      RECT -116.535000  139.260000 -101.220000  141.625000 ;
      RECT -116.285000  -78.195000 -100.340000  -76.460000 ;
      RECT -116.285000  -76.460000 -102.150000  -74.650000 ;
      RECT -116.280000  -56.970000 -110.000000  -54.300000 ;
      RECT -116.280000   55.330000 -110.000000   56.970000 ;
      RECT -116.225000   96.810000 -101.215000   99.480000 ;
      RECT -116.040000  118.035000 -103.030000  119.615000 ;
      RECT -116.040000  119.615000  -99.640000  120.895000 ;
      RECT -115.355000  120.895000  -99.640000  121.580000 ;
      RECT -115.350000   75.620000 -101.180000   79.130000 ;
      RECT -115.255000  141.625000 -101.220000  142.795000 ;
      RECT -115.255000  142.795000  -97.685000  142.905000 ;
      RECT -114.490000 -122.445000  -99.480000 -119.775000 ;
      RECT -114.490000 -119.775000 -103.030000 -118.900000 ;
      RECT -113.615000  -80.865000  -97.670000  -79.130000 ;
      RECT -113.615000  -79.130000 -100.340000  -78.195000 ;
      RECT -113.615000  -59.635000 -110.000000  -56.970000 ;
      RECT -113.615000   56.970000 -110.000000   58.005000 ;
      RECT -113.615000   58.005000  -97.565000   59.635000 ;
      RECT -113.610000 -102.095000  -96.805000 -101.220000 ;
      RECT -113.610000 -101.220000  -99.480000  -98.545000 ;
      RECT -112.680000   79.130000  -97.670000   81.800000 ;
      RECT -112.675000   99.480000  -98.545000  102.150000 ;
      RECT -112.675000  102.150000  -95.875000  103.030000 ;
      RECT -111.820000  121.580000  -99.640000  122.445000 ;
      RECT -111.820000  122.445000  -96.810000  125.110000 ;
      RECT -111.820000  125.110000  -94.145000  125.115000 ;
      RECT -110.945000 -125.990000  -94.145000 -125.110000 ;
      RECT -110.945000 -125.110000  -96.810000 -122.445000 ;
      RECT -110.940000 -104.765000  -96.805000 -102.095000 ;
      RECT -110.940000  -83.540000  -95.000000  -81.800000 ;
      RECT -110.940000  -81.800000  -97.670000  -80.865000 ;
      RECT -110.940000  103.030000  -95.875000  104.765000 ;
      RECT -110.065000  -63.185000 -110.000000  -59.635000 ;
      RECT -110.065000   59.635000  -97.565000   63.185000 ;
      RECT -110.010000   81.800000  -95.000000   84.470000 ;
      RECT -109.130000   63.185000  -97.565000   64.120000 ;
      RECT -109.025000  -64.225000  -92.385000  -63.185000 ;
      RECT -108.275000 -107.430000  -91.560000 -106.465000 ;
      RECT -108.275000 -106.465000  -93.260000 -104.765000 ;
      RECT -108.275000  104.765000  -93.260000  107.430000 ;
      RECT -108.275000  125.115000  -94.145000  128.660000 ;
      RECT -107.435000 -129.500000  -90.595000 -128.660000 ;
      RECT -107.435000 -128.660000  -94.145000 -125.990000 ;
      RECT -107.395000  -87.085000  -92.330000  -84.470000 ;
      RECT -107.395000  -84.470000  -95.000000  -83.540000 ;
      RECT -107.395000   84.470000  -92.330000   87.085000 ;
      RECT -106.465000   87.085000  -92.330000   87.140000 ;
      RECT -106.465000   87.140000  -89.660000   88.015000 ;
      RECT -106.460000  -66.790000  -92.385000  -64.225000 ;
      RECT -106.460000   64.120000  -97.565000   66.790000 ;
      RECT -105.695000  -88.785000  -89.715000  -87.085000 ;
      RECT -104.765000  128.660000  -90.595000  132.155000 ;
      RECT -104.765000  132.155000  -87.100000  132.170000 ;
      RECT -104.725000 -110.980000  -88.015000 -110.010000 ;
      RECT -104.725000 -110.010000  -91.560000 -107.430000 ;
      RECT -104.725000   88.015000  -89.660000   89.755000 ;
      RECT -104.725000  107.430000  -93.260000  107.435000 ;
      RECT -104.725000  107.435000  -90.590000  110.010000 ;
      RECT -104.725000  110.010000  -88.015000  110.980000 ;
      RECT -103.890000 -133.045000  -87.085000 -132.170000 ;
      RECT -103.890000 -132.170000  -90.595000 -129.500000 ;
      RECT -103.845000  -69.405000  -92.385000  -66.790000 ;
      RECT -103.790000   66.790000  -97.565000   69.460000 ;
      RECT -102.820000  110.980000  -88.015000  112.885000 ;
      RECT -102.150000  -92.330000  -87.140000  -89.660000 ;
      RECT -102.150000  -89.660000  -89.715000  -88.785000 ;
      RECT -102.150000   89.755000  -89.660000   90.690000 ;
      RECT -102.150000   90.690000  -86.110000   92.330000 ;
      RECT -101.525000  142.905000  -97.685000  146.340000 ;
      RECT -101.525000  146.340000  -94.140000  149.850000 ;
      RECT -101.525000  149.850000  -90.630000  153.395000 ;
      RECT -101.525000  153.395000  -87.085000  156.635000 ;
      RECT -101.270000  -71.980000  -92.385000  -69.405000 ;
      RECT -101.220000  132.170000  -87.100000  134.840000 ;
      RECT -101.220000  134.840000  -84.415000  135.715000 ;
      RECT -101.215000 -114.490000  -84.470000 -113.555000 ;
      RECT -101.215000 -113.555000  -88.015000 -110.980000 ;
      RECT -101.180000   92.330000  -86.110000   93.300000 ;
      RECT -100.355000 -157.805000  -86.220000 -154.260000 ;
      RECT -100.355000 -154.260000  -89.755000 -150.725000 ;
      RECT -100.355000 -150.725000  -93.300000 -147.180000 ;
      RECT -100.355000 -147.180000  -96.810000 -143.670000 ;
      RECT -100.355000 -136.580000  -84.625000 -134.630000 ;
      RECT -100.355000 -134.630000  -87.085000 -133.045000 ;
      RECT -100.245000  156.635000  -87.085000  156.940000 ;
      RECT -100.245000  156.940000  -83.540000  157.915000 ;
      RECT -100.240000   69.460000  -97.565000   73.010000 ;
      RECT  -99.480000 -116.225000  -84.470000 -114.490000 ;
      RECT  -99.480000  112.885000  -85.140000  116.225000 ;
      RECT  -98.605000  -95.875000  -82.660000  -94.140000 ;
      RECT  -98.605000  -94.140000  -84.470000  -92.330000 ;
      RECT  -98.600000  -74.650000  -92.385000  -71.980000 ;
      RECT  -97.675000  135.715000  -84.415000  138.390000 ;
      RECT  -97.675000  138.390000  -80.865000  139.260000 ;
      RECT  -97.670000   93.300000  -83.500000   96.810000 ;
      RECT  -97.630000   73.010000  -97.565000   75.620000 ;
      RECT  -96.810000 -140.125000  -81.800000 -137.455000 ;
      RECT  -96.810000 -137.455000  -84.625000 -136.580000 ;
      RECT  -96.790000  -76.460000  -92.385000  -74.650000 ;
      RECT  -96.090000  116.225000  -81.800000  119.615000 ;
      RECT  -95.985000  157.915000  -83.540000  160.475000 ;
      RECT  -95.985000  160.475000  -80.005000  162.175000 ;
      RECT  -95.935000  -98.545000  -79.990000  -96.810000 ;
      RECT  -95.935000  -96.810000  -82.660000  -95.875000 ;
      RECT  -95.930000 -119.775000  -79.125000 -118.900000 ;
      RECT  -95.930000 -118.900000  -81.800000 -116.225000 ;
      RECT  -95.310000  139.260000  -80.865000  140.125000 ;
      RECT  -95.310000  140.125000  -79.130000  141.625000 ;
      RECT  -95.000000   96.810000  -79.990000   99.480000 ;
      RECT  -94.995000  119.615000  -78.410000  120.710000 ;
      RECT  -94.140000  141.625000  -79.130000  142.790000 ;
      RECT  -94.140000  142.790000  -76.465000  142.795000 ;
      RECT  -94.120000  -79.130000  -92.385000  -76.460000 ;
      RECT  -94.120000   75.620000  -79.950000   79.130000 ;
      RECT  -93.265000 -143.670000  -76.350000 -142.905000 ;
      RECT  -93.265000 -142.905000  -79.130000 -140.125000 ;
      RECT  -93.260000 -122.445000  -79.125000 -119.775000 ;
      RECT  -93.260000 -101.220000  -77.320000  -99.480000 ;
      RECT  -93.260000  -99.480000  -79.990000  -98.545000 ;
      RECT  -93.260000  120.710000  -78.410000  122.445000 ;
      RECT  -92.330000   99.480000  -77.320000  102.150000 ;
      RECT  -91.450000  -81.800000  -74.705000  -80.865000 ;
      RECT  -91.450000   79.130000  -79.950000   81.800000 ;
      RECT  -90.595000 -125.110000  -73.015000 -125.010000 ;
      RECT  -90.595000 -125.010000  -75.580000 -122.445000 ;
      RECT  -90.595000  122.445000  -75.580000  125.110000 ;
      RECT  -90.595000  142.795000  -76.465000  145.375000 ;
      RECT  -90.595000  145.375000  -73.880000  146.340000 ;
      RECT  -89.755000 -147.180000  -72.915000 -146.340000 ;
      RECT  -89.755000 -146.340000  -76.350000 -143.670000 ;
      RECT  -89.715000 -104.765000  -74.650000 -102.150000 ;
      RECT  -89.715000 -102.150000  -77.320000 -101.220000 ;
      RECT  -89.715000  102.150000  -74.650000  104.765000 ;
      RECT  -89.090000  125.110000  -75.580000  125.115000 ;
      RECT  -89.090000  125.115000  -72.910000  126.615000 ;
      RECT  -88.785000  104.765000  -74.650000  104.820000 ;
      RECT  -88.785000  104.820000  -71.980000  105.695000 ;
      RECT  -88.780000  -84.470000  -74.705000  -81.800000 ;
      RECT  -88.780000   81.800000  -79.950000   84.470000 ;
      RECT  -88.120000  162.175000  -80.005000  164.020000 ;
      RECT  -88.120000  164.020000  -76.460000  167.530000 ;
      RECT  -88.120000  167.530000  -72.950000  170.040000 ;
      RECT  -88.015000 -106.465000  -72.035000 -104.765000 ;
      RECT  -87.085000  146.340000  -73.880000  148.445000 ;
      RECT  -87.085000  148.445000  -70.810000  149.850000 ;
      RECT  -87.045000 -128.660000  -70.125000 -127.900000 ;
      RECT  -87.045000 -127.900000  -73.015000 -125.110000 ;
      RECT  -87.045000  105.695000  -71.980000  107.435000 ;
      RECT  -87.045000  126.615000  -72.910000  128.660000 ;
      RECT  -86.210000 -150.725000  -69.405000 -149.850000 ;
      RECT  -86.210000 -149.850000  -72.915000 -147.180000 ;
      RECT  -86.165000  -87.085000  -74.705000  -84.470000 ;
      RECT  -86.110000   84.470000  -79.950000   87.140000 ;
      RECT  -84.470000 -110.010000  -69.460000 -107.340000 ;
      RECT  -84.470000 -107.340000  -72.035000 -106.465000 ;
      RECT  -84.470000  107.435000  -71.980000  108.370000 ;
      RECT  -84.470000  108.370000  -68.430000  110.010000 ;
      RECT  -83.590000  -89.660000  -74.705000  -87.085000 ;
      RECT  -83.550000  128.660000  -69.365000  132.155000 ;
      RECT  -83.540000  149.850000  -70.810000  151.585000 ;
      RECT  -83.540000  151.585000  -67.670000  153.395000 ;
      RECT  -83.535000 -132.170000  -66.790000 -131.235000 ;
      RECT  -83.535000 -131.235000  -70.125000 -128.660000 ;
      RECT  -82.765000 -175.395000  -10.800000 -171.140000 ;
      RECT  -82.765000 -171.140000  -11.900000 -170.040000 ;
      RECT  -82.765000 -170.040000  -72.950000 -167.530000 ;
      RECT  -82.765000 -167.530000  -75.620000 -164.860000 ;
      RECT  -82.765000 -164.860000  -79.130000 -161.350000 ;
      RECT  -82.765000 -161.350000  -82.675000 -157.805000 ;
      RECT  -82.675000 -154.260000  -67.670000 -151.585000 ;
      RECT  -82.675000 -151.585000  -69.405000 -150.725000 ;
      RECT  -82.560000   87.140000  -79.950000   90.690000 ;
      RECT  -81.595000  110.010000  -68.430000  111.820000 ;
      RECT  -81.595000  111.820000  -64.980000  112.885000 ;
      RECT  -81.075000 -134.630000  -66.790000 -132.170000 ;
      RECT  -80.925000 -113.555000  -64.980000 -111.820000 ;
      RECT  -80.925000 -111.820000  -66.790000 -110.010000 ;
      RECT  -80.920000  -92.330000  -74.705000  -89.660000 ;
      RECT  -80.865000  132.155000  -65.870000  134.625000 ;
      RECT  -80.865000  134.625000  -63.400000  134.840000 ;
      RECT  -80.300000  153.395000  -67.670000  155.030000 ;
      RECT  -80.300000  155.030000  -11.340000  156.130000 ;
      RECT  -80.300000  156.130000  -10.240000  156.635000 ;
      RECT  -79.995000  156.635000  -10.240000  156.940000 ;
      RECT  -79.950000   92.330000  -63.240000   93.300000 ;
      RECT  -79.130000 -157.805000   -4.895000 -155.030000 ;
      RECT  -79.130000 -155.030000  -67.670000 -154.260000 ;
      RECT  -79.110000  -94.140000  -74.705000  -92.330000 ;
      RECT  -78.255000 -116.225000  -62.310000 -114.490000 ;
      RECT  -78.255000 -114.490000  -64.980000 -113.555000 ;
      RECT  -78.255000  112.885000  -64.980000  115.355000 ;
      RECT  -78.255000  115.355000  -61.445000  116.225000 ;
      RECT  -78.250000 -137.455000  -63.395000 -134.630000 ;
      RECT  -77.315000  134.840000  -63.400000  137.510000 ;
      RECT  -77.315000  137.510000  -60.515000  138.390000 ;
      RECT  -76.460000  156.940000  -10.240000  160.475000 ;
      RECT  -76.440000  -96.810000  -74.705000  -94.140000 ;
      RECT  -76.440000   93.300000  -63.240000   96.810000 ;
      RECT  -75.620000 -182.540000  -11.900000 -181.440000 ;
      RECT  -75.620000 -181.440000  -10.800000 -175.395000 ;
      RECT  -75.620000  170.040000   75.620000  182.540000 ;
      RECT  -75.585000 -161.350000   -4.895000 -157.805000 ;
      RECT  -75.580000 -140.125000  -11.900000 -140.020000 ;
      RECT  -75.580000 -140.020000  -60.515000 -137.510000 ;
      RECT  -75.580000 -137.510000  -63.395000 -137.455000 ;
      RECT  -75.580000 -118.900000  -59.640000 -117.160000 ;
      RECT  -75.580000 -117.160000  -62.310000 -116.225000 ;
      RECT  -75.580000  138.390000  -60.515000  140.020000 ;
      RECT  -75.580000  140.020000   -4.895000  140.125000 ;
      RECT  -74.865000  116.225000  -61.445000  118.425000 ;
      RECT  -74.865000  118.425000  -58.375000  119.615000 ;
      RECT  -73.770000  -99.480000  -57.025000  -98.545000 ;
      RECT  -73.770000   96.810000  -63.240000   99.480000 ;
      RECT  -72.915000  140.125000   -4.895000  142.790000 ;
      RECT  -72.915000  160.475000  -10.240000  164.020000 ;
      RECT  -72.800000 -142.905000  -10.800000 -141.120000 ;
      RECT  -72.800000 -141.120000  -11.900000 -140.125000 ;
      RECT  -72.075000 -164.860000   -4.895000 -161.350000 ;
      RECT  -72.035000 -122.445000  -56.970000 -119.830000 ;
      RECT  -72.035000 -119.830000  -59.640000 -118.900000 ;
      RECT  -72.035000  119.615000  -58.375000  121.470000 ;
      RECT  -72.035000  121.470000  -55.330000  122.445000 ;
      RECT  -71.105000  122.445000  -55.330000  123.375000 ;
      RECT  -71.100000 -102.150000  -57.025000  -99.480000 ;
      RECT  -71.100000   99.480000  -63.240000  102.150000 ;
      RECT  -70.330000  142.790000   -4.895000  145.375000 ;
      RECT  -69.470000 -125.010000  -54.355000 -122.445000 ;
      RECT  -69.405000 -167.530000   -4.895000 -164.860000 ;
      RECT  -69.405000  164.020000  -10.240000  166.430000 ;
      RECT  -69.405000  166.430000  -11.340000  167.530000 ;
      RECT  -69.365000 -146.340000  -10.800000 -142.905000 ;
      RECT  -69.365000  123.375000  -55.330000  125.010000 ;
      RECT  -69.365000  125.010000  -11.340000  125.115000 ;
      RECT  -68.485000 -104.765000  -57.025000 -102.150000 ;
      RECT  -68.430000  102.150000  -63.240000  104.820000 ;
      RECT  -67.865000  125.115000  -11.340000  126.110000 ;
      RECT  -67.865000  126.110000  -10.240000  126.615000 ;
      RECT  -67.260000  145.375000   -4.895000  146.340000 ;
      RECT  -67.260000  146.340000    1.425000  148.445000 ;
      RECT  -66.580000 -127.900000   -4.895000 -125.010000 ;
      RECT  -65.910000 -107.340000  -57.025000 -104.765000 ;
      RECT  -65.855000 -149.850000  -10.800000 -146.340000 ;
      RECT  -65.820000  126.615000  -10.240000  128.660000 ;
      RECT  -64.880000  104.820000  -63.240000  108.370000 ;
      RECT  -64.120000 -151.585000  -11.900000 -151.420000 ;
      RECT  -64.120000 -151.420000  -10.800000 -149.850000 ;
      RECT  -64.120000  148.445000    1.425000  151.585000 ;
      RECT  -63.245000 -131.235000   -4.895000 -127.900000 ;
      RECT  -63.240000 -110.010000   61.430000 -110.000000 ;
      RECT  -63.240000 -110.000000  -57.025000 -107.340000 ;
      RECT  -63.240000  110.000000   -4.895000  110.010000 ;
      RECT  -63.185000 -152.520000  -11.900000 -151.585000 ;
      RECT  -63.185000  151.585000    1.425000  152.520000 ;
      RECT  -62.325000  128.660000  -10.240000  132.155000 ;
      RECT  -61.430000 -111.820000   61.430000 -110.010000 ;
      RECT  -61.430000  110.010000   -4.895000  111.820000 ;
      RECT  -59.855000  132.155000  -10.240000  134.625000 ;
      RECT  -59.850000 -134.630000   -4.895000 -131.235000 ;
      RECT  -58.760000 -114.490000   58.760000 -111.820000 ;
      RECT  -57.895000  111.820000   -4.895000  114.490000 ;
      RECT  -57.895000  114.490000   -0.405000  115.355000 ;
      RECT  -56.970000 -137.510000   -4.895000 -134.630000 ;
      RECT  -56.970000  134.625000  -10.240000  136.410000 ;
      RECT  -56.970000  136.410000  -11.340000  137.510000 ;
      RECT  -56.090000 -117.160000   56.090000 -114.490000 ;
      RECT  -54.825000  115.355000   -0.405000  118.425000 ;
      RECT  -53.420000 -119.830000   53.420000 -117.160000 ;
      RECT  -51.780000  118.425000   -0.405000  121.470000 ;
      RECT  -50.805000 -122.445000   50.750000 -119.830000 ;
      RECT  -50.750000 -122.500000   50.750000 -122.445000 ;
      RECT  -50.750000  121.470000   -0.405000  122.500000 ;
      RECT   -7.565000 -170.040000   -4.895000 -167.530000 ;
      RECT   -7.565000 -140.020000   -4.895000 -137.510000 ;
      RECT   -7.565000  122.500000   -0.405000  125.010000 ;
      RECT   -7.565000  152.520000    1.425000  155.030000 ;
      RECT   -7.460000 -140.125000   73.765000 -140.020000 ;
      RECT   -0.405000  125.010000   66.790000  127.690000 ;
      RECT   -0.405000  127.690000   63.245000  131.235000 ;
      RECT   -0.405000  131.235000   60.515000  132.170000 ;
      RECT    1.425000  155.030000   79.130000  157.805000 ;
      RECT    1.425000  157.805000   75.585000  161.350000 ;
      RECT    1.425000  161.350000   72.915000  164.020000 ;
      RECT    2.265000  132.170000   60.515000  133.965000 ;
      RECT    2.265000  133.965000   56.970000  134.840000 ;
      RECT    4.935000 -182.540000   75.620000 -170.040000 ;
      RECT    4.935000 -152.520000   63.185000 -149.850000 ;
      RECT    4.935000 -149.850000   65.855000 -146.340000 ;
      RECT    4.935000 -146.340000   69.365000 -142.790000 ;
      RECT    4.935000 -142.790000   72.915000 -141.940000 ;
      RECT    4.935000 -141.940000   73.765000 -140.125000 ;
      RECT    4.935000  134.840000   56.970000  137.510000 ;
      RECT    4.935000  164.020000   69.405000  167.530000 ;
      RECT   11.455000 -166.430000   69.405000 -164.860000 ;
      RECT   11.455000 -164.860000   72.075000 -161.315000 ;
      RECT   11.455000 -161.315000   75.620000 -157.770000 ;
      RECT   11.455000 -157.770000   79.165000 -156.940000 ;
      RECT   11.455000 -156.940000   79.995000 -156.130000 ;
      RECT   11.455000 -136.410000   56.970000 -134.840000 ;
      RECT   11.455000 -134.840000   59.640000 -132.170000 ;
      RECT   11.455000 -132.170000   62.310000 -128.660000 ;
      RECT   11.455000 -128.660000   65.820000 -126.110000 ;
      RECT   12.015000  111.100000   58.760000  114.490000 ;
      RECT   12.015000  114.490000   56.090000  117.160000 ;
      RECT   12.015000  117.160000   53.420000  119.830000 ;
      RECT   12.015000  119.830000   51.780000  121.400000 ;
      RECT   12.015000  141.120000   72.915000  142.790000 ;
      RECT   12.015000  142.790000   69.365000  146.340000 ;
      RECT   12.015000  146.340000   65.855000  149.850000 ;
      RECT   12.015000  149.850000   64.120000  151.420000 ;
      RECT   12.555000 -167.530000   69.405000 -166.430000 ;
      RECT   12.555000 -156.130000   79.995000 -155.030000 ;
      RECT   12.555000 -137.510000   56.970000 -136.410000 ;
      RECT   12.555000 -126.110000   65.820000 -125.115000 ;
      RECT   12.555000 -125.115000   69.365000 -125.010000 ;
      RECT   13.115000  110.000000   63.240000  110.010000 ;
      RECT   13.115000  110.010000   62.270000  110.980000 ;
      RECT   13.115000  110.980000   58.760000  111.100000 ;
      RECT   13.115000  121.400000   51.780000  121.470000 ;
      RECT   13.115000  121.470000   50.750000  122.500000 ;
      RECT   13.115000  140.020000   75.580000  140.125000 ;
      RECT   13.115000  140.125000   72.915000  141.120000 ;
      RECT   13.115000  151.420000   64.120000  151.585000 ;
      RECT   13.115000  151.585000   63.185000  152.520000 ;
      RECT   50.750000 -110.000000   61.430000 -108.370000 ;
      RECT   50.750000 -108.370000   64.880000 -104.820000 ;
      RECT   54.300000 -125.010000   69.365000 -123.375000 ;
      RECT   54.300000 -123.375000   71.105000 -122.500000 ;
      RECT   54.300000  122.500000   70.335000  124.145000 ;
      RECT   54.300000  124.145000   66.790000  125.010000 ;
      RECT   55.330000  121.470000   72.035000  122.445000 ;
      RECT   55.330000  122.445000   70.335000  122.500000 ;
      RECT   56.970000 -122.500000   71.105000 -119.830000 ;
      RECT   56.970000  119.830000   72.035000  121.470000 ;
      RECT   57.025000 -104.820000   68.430000 -102.150000 ;
      RECT   57.025000 -102.150000   71.100000  -99.480000 ;
      RECT   57.025000  -99.480000   73.770000  -98.545000 ;
      RECT   59.640000 -119.830000   74.650000 -117.160000 ;
      RECT   59.640000  117.160000   75.580000  118.900000 ;
      RECT   59.640000  118.900000   72.035000  119.830000 ;
      RECT   60.515000 -140.020000   73.765000 -138.390000 ;
      RECT   60.515000 -138.390000   77.315000 -137.510000 ;
      RECT   60.515000  137.510000   75.580000  140.020000 ;
      RECT   62.310000 -117.160000   77.320000 -114.490000 ;
      RECT   62.310000  114.490000   78.255000  116.225000 ;
      RECT   62.310000  116.225000   75.580000  117.160000 ;
      RECT   63.185000 -137.510000   77.315000 -134.840000 ;
      RECT   63.240000   92.330000   79.950000   93.300000 ;
      RECT   63.240000   93.300000   76.440000   96.810000 ;
      RECT   63.240000   96.810000   73.010000  100.240000 ;
      RECT   63.240000  100.240000   69.460000  103.790000 ;
      RECT   63.240000  103.790000   65.910000  107.340000 ;
      RECT   64.060000  133.965000   78.250000  137.455000 ;
      RECT   64.060000  137.455000   75.580000  137.510000 ;
      RECT   64.980000 -114.490000   79.990000 -111.820000 ;
      RECT   65.820000  110.980000   80.925000  113.555000 ;
      RECT   65.820000  113.555000   78.255000  114.490000 ;
      RECT   65.855000 -134.840000   80.865000 -132.170000 ;
      RECT   66.735000 -155.030000   79.995000 -153.395000 ;
      RECT   66.735000 -153.395000   83.540000 -152.520000 ;
      RECT   66.735000  152.520000   82.675000  154.260000 ;
      RECT   66.735000  154.260000   79.130000  155.030000 ;
      RECT   66.790000  110.010000   80.925000  110.980000 ;
      RECT   66.790000  131.235000   81.800000  133.905000 ;
      RECT   66.790000  133.905000   78.250000  133.965000 ;
      RECT   67.670000  151.585000   82.675000  152.520000 ;
      RECT   68.430000 -111.820000   79.990000 -110.980000 ;
      RECT   68.430000 -110.980000   83.500000 -108.370000 ;
      RECT   68.430000  -98.545000   73.770000  -96.810000 ;
      RECT   68.430000  -96.810000   76.440000  -94.140000 ;
      RECT   68.430000  -94.140000   79.110000  -90.690000 ;
      RECT   68.430000  -90.690000   82.560000  -87.140000 ;
      RECT   69.365000 -132.170000   83.535000 -128.660000 ;
      RECT   69.405000 -152.520000   83.540000 -149.850000 ;
      RECT   69.405000  149.850000   86.220000  150.715000 ;
      RECT   69.405000  150.715000   82.675000  151.585000 ;
      RECT   69.460000  107.340000   84.470000  110.010000 ;
      RECT   70.335000  127.690000   87.045000  128.660000 ;
      RECT   70.335000  128.660000   85.350000  130.355000 ;
      RECT   70.335000  130.355000   81.800000  131.235000 ;
      RECT   71.980000 -108.370000   83.500000 -107.435000 ;
      RECT   71.980000 -107.435000   87.045000 -105.695000 ;
      RECT   71.980000 -105.695000   88.785000 -104.820000 ;
      RECT   72.910000 -128.660000   87.045000 -125.115000 ;
      RECT   72.915000 -149.850000   87.085000 -147.180000 ;
      RECT   72.915000 -147.180000   89.755000 -146.340000 ;
      RECT   72.915000  146.340000   89.755000  147.180000 ;
      RECT   72.915000  147.180000   86.220000  149.850000 ;
      RECT   72.950000 -170.040000   75.620000 -167.530000 ;
      RECT   72.950000  167.530000   88.120000  170.040000 ;
      RECT   73.010000  103.790000   89.715000  104.765000 ;
      RECT   73.010000  104.765000   88.015000  106.465000 ;
      RECT   73.010000  106.465000   84.470000  107.340000 ;
      RECT   73.015000 -125.115000   87.045000 -125.110000 ;
      RECT   73.015000 -125.110000   90.595000 -125.010000 ;
      RECT   73.880000  124.145000   90.595000  125.110000 ;
      RECT   73.880000  125.110000   87.045000  127.690000 ;
      RECT   74.650000 -125.010000   90.595000 -124.260000 ;
      RECT   74.650000 -124.260000   91.445000 -123.375000 ;
      RECT   74.650000 -104.820000   88.785000 -102.150000 ;
      RECT   74.705000  -87.140000   86.110000  -84.470000 ;
      RECT   74.705000  -84.470000   88.780000  -81.800000 ;
      RECT   74.705000  -81.800000   91.450000  -80.865000 ;
      RECT   75.580000  122.445000   90.595000  124.145000 ;
      RECT   75.620000 -167.530000   90.630000 -164.860000 ;
      RECT   76.460000  164.020000   88.120000  167.530000 ;
      RECT   76.465000 -146.340000   89.755000 -143.635000 ;
      RECT   76.465000 -143.635000   93.300000 -142.790000 ;
      RECT   76.465000  142.790000   93.265000  143.670000 ;
      RECT   76.465000  143.670000   89.755000  146.340000 ;
      RECT   76.560000  100.240000   93.260000  101.220000 ;
      RECT   76.560000  101.220000   89.715000  103.790000 ;
      RECT   77.315000 -142.790000   93.300000 -141.940000 ;
      RECT   77.320000 -102.150000   92.330000  -99.480000 ;
      RECT   78.195000 -123.375000   91.445000 -120.710000 ;
      RECT   78.195000 -120.710000   94.995000 -119.830000 ;
      RECT   79.125000  118.900000   95.930000  119.775000 ;
      RECT   79.125000  119.775000   93.260000  122.445000 ;
      RECT   79.130000  140.125000   93.265000  142.790000 ;
      RECT   79.130000  161.350000   88.120000  164.020000 ;
      RECT   79.165000 -164.860000   90.630000 -161.315000 ;
      RECT   79.235000 -141.940000   93.300000 -140.090000 ;
      RECT   79.235000 -140.090000   96.845000 -140.020000 ;
      RECT   79.950000   75.620000   94.120000   79.130000 ;
      RECT   79.950000   79.130000   90.690000   82.560000 ;
      RECT   79.950000   82.560000   87.140000   86.110000 ;
      RECT   79.950000   86.110000   83.590000   89.660000 ;
      RECT   79.950000   89.660000   80.920000   92.330000 ;
      RECT   79.990000  -99.480000   95.000000  -96.810000 ;
      RECT   79.990000   96.810000   95.935000   98.545000 ;
      RECT   79.990000   98.545000   93.260000  100.240000 ;
      RECT   80.865000 -140.020000   96.845000 -139.260000 ;
      RECT   80.865000 -139.260000   97.675000 -138.390000 ;
      RECT   80.865000 -119.830000   94.995000 -117.160000 ;
      RECT   80.920000   74.650000   97.630000   75.620000 ;
      RECT   81.800000  116.225000   95.930000  118.900000 ;
      RECT   81.800000  137.455000   96.810000  140.125000 ;
      RECT   82.660000  -96.810000   97.670000  -94.140000 ;
      RECT   82.675000  157.805000   88.120000  161.350000 ;
      RECT   82.710000 -161.315000   90.630000 -157.770000 ;
      RECT   83.500000   93.300000   98.605000   95.875000 ;
      RECT   83.500000   95.875000   95.935000   96.810000 ;
      RECT   83.535000 -117.160000   98.545000 -114.490000 ;
      RECT   83.540000 -157.770000   90.630000 -156.940000 ;
      RECT   84.415000 -138.390000   97.675000 -135.715000 ;
      RECT   84.415000 -135.715000  101.220000 -134.840000 ;
      RECT   84.470000   92.330000   98.605000   93.300000 ;
      RECT   84.470000  113.555000   99.480000  116.225000 ;
      RECT   85.130000  -80.865000   91.450000  -79.130000 ;
      RECT   85.130000  -79.130000   94.120000  -76.460000 ;
      RECT   85.130000  -76.460000   96.790000  -73.010000 ;
      RECT   85.130000  -73.010000  100.240000  -70.440000 ;
      RECT   85.350000  133.905000  100.355000  136.580000 ;
      RECT   85.350000  136.580000   96.810000  137.455000 ;
      RECT   86.110000  -94.140000   97.670000  -93.300000 ;
      RECT   86.110000  -93.300000  101.180000  -90.690000 ;
      RECT   86.220000  154.260000  100.355000  157.805000 ;
      RECT   87.045000 -114.490000  101.215000 -110.980000 ;
      RECT   87.085000 -156.940000   90.630000 -153.395000 ;
      RECT   87.085000 -134.840000  101.220000 -132.170000 ;
      RECT   87.140000   89.660000  102.150000   92.330000 ;
      RECT   88.015000  110.010000  104.725000  110.980000 ;
      RECT   88.015000  110.980000  103.030000  112.675000 ;
      RECT   88.015000  112.675000   99.480000  113.555000 ;
      RECT   88.900000  130.355000  103.900000  133.035000 ;
      RECT   88.900000  133.035000  100.355000  133.905000 ;
      RECT   89.660000  -90.690000  101.180000  -89.755000 ;
      RECT   89.660000  -89.755000  104.725000  -88.015000 ;
      RECT   89.660000  -88.015000  106.465000  -87.140000 ;
      RECT   89.765000  150.715000  100.355000  154.260000 ;
      RECT   90.590000 -110.980000  104.725000 -107.435000 ;
      RECT   90.595000 -132.170000  104.765000 -129.500000 ;
      RECT   90.595000 -129.500000  107.435000 -128.660000 ;
      RECT   90.595000  128.660000  107.435000  129.500000 ;
      RECT   90.595000  129.500000  103.900000  130.355000 ;
      RECT   90.690000   86.110000  107.395000   87.085000 ;
      RECT   90.690000   87.085000  105.695000   88.785000 ;
      RECT   90.690000   88.785000  102.150000   89.660000 ;
      RECT   91.560000  106.465000  108.275000  107.430000 ;
      RECT   91.560000  107.430000  104.725000  110.010000 ;
      RECT   92.330000 -107.435000  104.725000 -107.430000 ;
      RECT   92.330000 -107.430000  108.275000 -106.580000 ;
      RECT   92.330000 -106.580000  109.125000 -105.695000 ;
      RECT   92.330000  -87.140000  106.465000  -84.470000 ;
      RECT   92.385000  -70.440000  100.240000  -69.460000 ;
      RECT   92.385000  -69.460000  103.790000  -66.790000 ;
      RECT   92.385000  -66.790000  106.460000  -64.225000 ;
      RECT   92.385000  -64.225000  109.025000  -63.185000 ;
      RECT   93.260000  104.765000  108.275000  106.465000 ;
      RECT   93.300000 -149.850000  108.310000 -147.180000 ;
      RECT   93.300000  147.180000  100.355000  150.715000 ;
      RECT   94.145000 -128.660000  107.435000 -125.955000 ;
      RECT   94.145000 -125.955000  110.980000 -125.110000 ;
      RECT   94.145000  125.110000  110.945000  125.990000 ;
      RECT   94.145000  125.990000  107.435000  128.660000 ;
      RECT   94.240000   82.560000  110.940000   83.540000 ;
      RECT   94.240000   83.540000  107.395000   86.110000 ;
      RECT   94.995000 -125.110000  110.980000 -124.260000 ;
      RECT   95.000000  -84.470000  110.010000  -81.800000 ;
      RECT   95.875000 -105.695000  109.125000 -103.030000 ;
      RECT   95.875000 -103.030000  112.675000 -102.150000 ;
      RECT   96.805000  101.220000  113.610000  102.095000 ;
      RECT   96.805000  102.095000  110.940000  104.765000 ;
      RECT   96.810000  122.445000  110.945000  125.110000 ;
      RECT   96.810000  143.670000  100.355000  147.180000 ;
      RECT   96.845000 -147.180000  108.310000 -143.635000 ;
      RECT   97.565000  -63.185000  110.065000  -59.635000 ;
      RECT   97.565000  -59.635000  113.615000  -58.005000 ;
      RECT   97.565000   58.005000  113.615000   59.635000 ;
      RECT   97.565000   59.635000  110.065000   63.185000 ;
      RECT   97.565000   63.185000  108.370000   64.880000 ;
      RECT   97.565000   64.880000  104.820000   68.430000 ;
      RECT   97.565000   68.430000  101.270000   71.980000 ;
      RECT   97.565000   71.980000   98.600000   74.650000 ;
      RECT   97.670000  -81.800000  112.680000  -79.130000 ;
      RECT   97.670000   79.130000  113.615000   80.865000 ;
      RECT   97.670000   80.865000  110.940000   82.560000 ;
      RECT   98.545000 -124.260000  110.980000 -122.410000 ;
      RECT   98.545000 -122.410000  114.525000 -121.580000 ;
      RECT   98.545000 -121.580000  115.355000 -120.710000 ;
      RECT   98.545000 -102.150000  112.675000  -99.480000 ;
      RECT   98.600000   56.970000  113.615000   58.005000 ;
      RECT   99.480000   98.545000  113.610000  101.220000 ;
      RECT   99.480000  119.775000  114.490000  122.445000 ;
      RECT  100.340000  -79.130000  115.350000  -76.460000 ;
      RECT  100.390000 -143.635000  108.310000 -140.090000 ;
      RECT  101.180000   75.620000  116.285000   78.195000 ;
      RECT  101.180000   78.195000  113.615000   79.130000 ;
      RECT  101.215000  -99.480000  116.225000  -96.810000 ;
      RECT  101.220000 -140.090000  108.310000 -139.260000 ;
      RECT  102.095000 -120.710000  115.355000 -118.035000 ;
      RECT  102.095000 -118.035000  118.900000 -117.160000 ;
      RECT  102.150000   74.650000  116.285000   75.620000 ;
      RECT  102.150000   95.875000  117.160000   98.545000 ;
      RECT  103.030000  116.225000  118.035000  118.900000 ;
      RECT  103.030000  118.900000  114.490000  119.775000 ;
      RECT  103.780000  -58.005000  115.245000  -55.330000 ;
      RECT  103.780000  -55.330000  117.920000  -51.790000 ;
      RECT  103.790000  -76.460000  115.350000  -75.620000 ;
      RECT  103.790000  -75.620000  118.860000  -73.010000 ;
      RECT  103.900000  136.580000  118.035000  140.125000 ;
      RECT  104.725000  -96.810000  118.895000  -93.300000 ;
      RECT  104.765000 -139.260000  108.310000 -135.715000 ;
      RECT  104.765000 -117.160000  118.900000 -114.490000 ;
      RECT  104.820000   71.980000  119.830000   74.650000 ;
      RECT  105.695000   92.330000  122.405000   93.300000 ;
      RECT  105.695000   93.300000  120.710000   94.995000 ;
      RECT  105.695000   94.995000  117.160000   95.875000 ;
      RECT  106.360000  -73.010000  118.860000  -72.075000 ;
      RECT  106.360000  -72.075000  122.405000  -70.440000 ;
      RECT  106.580000  112.675000  121.580000  115.355000 ;
      RECT  106.580000  115.355000  118.035000  116.225000 ;
      RECT  107.340000  -70.440000  122.405000  -70.335000 ;
      RECT  107.340000  -70.335000  124.145000  -69.460000 ;
      RECT  107.445000  133.035000  118.035000  136.580000 ;
      RECT  108.270000  -93.300000  122.405000  -89.755000 ;
      RECT  108.275000 -114.490000  122.445000 -111.820000 ;
      RECT  108.275000 -111.820000  125.115000 -110.980000 ;
      RECT  108.275000  110.980000  125.115000  111.820000 ;
      RECT  108.275000  111.820000  121.580000  112.675000 ;
      RECT  108.370000   68.430000  125.075000   69.405000 ;
      RECT  108.370000   69.405000  123.375000   71.105000 ;
      RECT  108.370000   71.105000  119.830000   71.980000 ;
      RECT  109.240000   88.785000  125.955000   89.750000 ;
      RECT  109.240000   89.750000  122.405000   92.330000 ;
      RECT  110.000000  -51.790000  121.460000  -50.750000 ;
      RECT  110.000000  -50.750000  122.500000   50.750000 ;
      RECT  110.000000   50.750000  118.950000   54.300000 ;
      RECT  110.000000   54.300000  116.280000   56.970000 ;
      RECT  110.010000  -89.755000  122.405000  -89.750000 ;
      RECT  110.010000  -89.750000  125.955000  -88.900000 ;
      RECT  110.010000  -88.900000  126.805000  -88.015000 ;
      RECT  110.010000  -69.460000  124.145000  -66.790000 ;
      RECT  110.940000   87.085000  125.955000   88.785000 ;
      RECT  110.980000 -132.170000  125.990000 -129.500000 ;
      RECT  110.980000  129.500000  118.035000  133.035000 ;
      RECT  111.825000 -110.980000  125.115000 -108.275000 ;
      RECT  111.825000 -108.275000  128.660000 -107.430000 ;
      RECT  111.825000  107.430000  128.625000  108.310000 ;
      RECT  111.825000  108.310000  125.115000  110.980000 ;
      RECT  111.920000   64.880000  128.620000   65.860000 ;
      RECT  111.920000   65.860000  125.075000   68.430000 ;
      RECT  112.575000  -66.790000  127.690000  -64.225000 ;
      RECT  112.675000 -107.430000  128.660000 -106.580000 ;
      RECT  113.555000  -88.015000  126.805000  -85.350000 ;
      RECT  113.555000  -85.350000  130.355000  -84.470000 ;
      RECT  113.615000  -64.225000  130.255000  -63.185000 ;
      RECT  113.615000   63.185000  128.620000   64.880000 ;
      RECT  114.485000   83.540000  131.290000   84.415000 ;
      RECT  114.485000   84.415000  128.620000   87.085000 ;
      RECT  114.490000  104.765000  128.625000  107.430000 ;
      RECT  114.490000  125.990000  118.035000  129.500000 ;
      RECT  114.525000 -129.500000  125.990000 -125.955000 ;
      RECT  116.225000 -106.580000  128.660000 -104.730000 ;
      RECT  116.225000 -104.730000  132.205000 -103.900000 ;
      RECT  116.225000 -103.900000  133.035000 -103.030000 ;
      RECT  116.225000  -84.470000  130.355000  -81.800000 ;
      RECT  117.160000   80.865000  131.290000   83.540000 ;
      RECT  117.160000  102.095000  132.170000  104.765000 ;
      RECT  117.165000  -63.185000  131.295000  -60.515000 ;
      RECT  117.165000  -60.515000  133.965000  -59.635000 ;
      RECT  117.165000   59.635000  133.965000   60.515000 ;
      RECT  117.165000   60.515000  131.295000   63.185000 ;
      RECT  118.070000 -125.955000  125.990000 -122.410000 ;
      RECT  118.795000  -59.635000  133.965000  -58.005000 ;
      RECT  118.895000  -81.800000  133.905000  -79.130000 ;
      RECT  118.900000 -122.410000  125.990000 -121.580000 ;
      RECT  119.775000 -103.030000  133.035000 -100.355000 ;
      RECT  119.775000 -100.355000  136.580000  -99.480000 ;
      RECT  119.830000   56.970000  133.965000   59.635000 ;
      RECT  119.830000   78.195000  134.840000   80.865000 ;
      RECT  120.710000   98.545000  135.715000  101.220000 ;
      RECT  120.710000  101.220000  132.170000  102.095000 ;
      RECT  121.470000  -58.005000  133.965000  -56.970000 ;
      RECT  121.470000  -56.970000  137.510000  -55.330000 ;
      RECT  121.580000  118.900000  135.715000  122.445000 ;
      RECT  122.405000  -79.130000  136.575000  -75.620000 ;
      RECT  122.445000 -121.580000  125.990000 -118.035000 ;
      RECT  122.445000  -99.480000  136.580000  -96.810000 ;
      RECT  122.500000   54.300000  137.510000   56.970000 ;
      RECT  123.375000   74.650000  140.085000   75.620000 ;
      RECT  123.375000   75.620000  138.390000   77.315000 ;
      RECT  123.375000   77.315000  134.840000   78.195000 ;
      RECT  124.260000   94.995000  139.260000   97.675000 ;
      RECT  124.260000   97.675000  135.715000   98.545000 ;
      RECT  125.010000  -55.330000  137.510000   54.300000 ;
      RECT  125.125000  115.355000  135.715000  118.900000 ;
      RECT  125.950000  -75.620000  140.085000  -72.075000 ;
      RECT  125.955000  -96.810000  140.125000  -94.140000 ;
      RECT  125.955000  -94.140000  142.795000  -93.300000 ;
      RECT  125.955000   93.300000  142.795000   94.140000 ;
      RECT  125.955000   94.140000  139.260000   94.995000 ;
      RECT  126.920000   71.105000  143.635000   72.070000 ;
      RECT  126.920000   72.070000  140.085000   74.650000 ;
      RECT  127.585000  -72.075000  140.085000  -72.070000 ;
      RECT  127.585000  -72.070000  143.635000  -70.440000 ;
      RECT  127.690000  -70.440000  145.265000  -70.335000 ;
      RECT  128.620000   69.405000  143.635000   71.105000 ;
      RECT  128.660000 -114.490000  143.670000 -111.820000 ;
      RECT  128.660000  111.820000  135.715000  115.355000 ;
      RECT  129.505000  -93.300000  142.795000  -90.595000 ;
      RECT  129.505000  -90.595000  146.340000  -89.750000 ;
      RECT  129.505000   89.750000  146.305000   90.630000 ;
      RECT  129.505000   90.630000  142.795000   93.300000 ;
      RECT  130.355000  -89.750000  146.340000  -88.900000 ;
      RECT  131.235000  -70.335000  145.265000  -67.670000 ;
      RECT  131.235000  -67.670000  148.035000  -66.790000 ;
      RECT  132.165000   65.860000  148.970000   66.735000 ;
      RECT  132.165000   66.735000  146.300000   69.405000 ;
      RECT  132.170000   87.085000  146.305000   89.750000 ;
      RECT  132.170000  108.310000  135.715000  111.820000 ;
      RECT  132.205000 -111.820000  143.670000 -108.275000 ;
      RECT  133.800000  -66.790000  148.035000  -64.225000 ;
      RECT  133.905000  -88.900000  146.340000  -87.050000 ;
      RECT  133.905000  -87.050000  149.885000  -86.220000 ;
      RECT  133.905000  -86.220000  150.715000  -85.350000 ;
      RECT  134.840000  -64.225000  151.480000  -63.185000 ;
      RECT  134.840000   63.185000  148.970000   65.860000 ;
      RECT  134.840000   84.415000  149.850000   87.085000 ;
      RECT  135.750000 -108.275000  143.670000 -104.730000 ;
      RECT  136.580000 -104.730000  143.670000 -103.900000 ;
      RECT  137.455000  -85.350000  150.715000  -82.675000 ;
      RECT  137.455000  -82.675000  154.260000  -81.800000 ;
      RECT  137.510000  -63.185000  152.520000  -60.515000 ;
      RECT  137.510000   60.515000  152.520000   63.185000 ;
      RECT  138.390000   80.865000  153.395000   83.540000 ;
      RECT  138.390000   83.540000  149.850000   84.415000 ;
      RECT  139.260000  101.220000  153.395000  104.765000 ;
      RECT  140.020000  -60.515000  152.520000   60.515000 ;
      RECT  140.125000 -103.900000  143.670000 -100.355000 ;
      RECT  140.125000  -81.800000  154.260000  -79.130000 ;
      RECT  141.940000   77.315000  156.940000   79.995000 ;
      RECT  141.940000   79.995000  153.395000   80.865000 ;
      RECT  142.805000   97.675000  153.395000  101.220000 ;
      RECT  143.635000  -79.130000  157.805000  -76.460000 ;
      RECT  143.635000  -76.460000  160.475000  -75.620000 ;
      RECT  143.635000   75.620000  160.475000   76.460000 ;
      RECT  143.635000   76.460000  156.940000   77.315000 ;
      RECT  146.340000  -96.810000  161.350000  -94.140000 ;
      RECT  146.340000   94.140000  153.395000   97.675000 ;
      RECT  147.185000  -75.620000  160.475000  -72.950000 ;
      RECT  147.185000  -72.950000  163.985000  -72.070000 ;
      RECT  147.185000   72.070000  163.985000   72.950000 ;
      RECT  147.185000   72.950000  160.475000   75.620000 ;
      RECT  148.815000  -72.070000  163.985000  -70.440000 ;
      RECT  149.850000   69.405000  163.985000   72.070000 ;
      RECT  149.850000   90.630000  153.395000   94.140000 ;
      RECT  149.885000  -94.140000  161.350000  -90.595000 ;
      RECT  151.585000  -70.440000  163.985000  -69.405000 ;
      RECT  151.585000  -69.405000  167.530000  -67.670000 ;
      RECT  152.520000   66.735000  167.530000   69.405000 ;
      RECT  153.430000  -90.595000  161.350000  -87.050000 ;
      RECT  154.260000  -87.050000  161.350000  -86.220000 ;
      RECT  155.030000  -67.670000  167.530000   66.735000 ;
      RECT  156.940000   83.540000  171.075000   87.085000 ;
      RECT  157.805000  -86.220000  161.350000  -82.675000 ;
      RECT  160.485000   79.995000  171.075000   83.540000 ;
      RECT  164.020000  -79.130000  179.030000  -76.460000 ;
      RECT  164.020000   76.460000  171.075000   79.995000 ;
      RECT  167.530000  -76.460000  179.030000  -75.620000 ;
      RECT  167.530000  -75.620000  182.540000  -72.950000 ;
      RECT  167.530000   72.950000  182.540000   75.620000 ;
      RECT  167.530000   75.620000  171.075000   76.460000 ;
      RECT  170.040000  -72.950000  182.540000  -27.500000 ;
      RECT  170.040000  -27.500000  187.540000  -15.000000 ;
      RECT  170.040000   15.000000  187.540000   27.500000 ;
      RECT  170.040000   27.500000  182.540000   72.950000 ;
    LAYER via2 ;
      RECT -37.220000 -180.935000 -35.940000 -179.655000 ;
      RECT -37.220000 -178.465000 -35.940000 -177.185000 ;
      RECT -37.220000 -175.395000 -35.940000 -174.115000 ;
      RECT -37.220000 -172.925000 -35.940000 -171.645000 ;
      RECT -37.220000 -150.915000 -35.940000 -149.635000 ;
      RECT -37.220000 -148.445000 -35.940000 -147.165000 ;
      RECT -37.220000 -145.375000 -35.940000 -144.095000 ;
      RECT -37.220000 -142.905000 -35.940000 -141.625000 ;
      RECT -36.655000  126.615000 -35.375000  127.895000 ;
      RECT -36.655000  129.085000 -35.375000  130.365000 ;
      RECT -36.655000  132.155000 -35.375000  133.435000 ;
      RECT -36.655000  134.625000 -35.375000  135.905000 ;
      RECT -36.655000  156.635000 -35.375000  157.915000 ;
      RECT -36.655000  159.105000 -35.375000  160.385000 ;
      RECT -36.655000  162.175000 -35.375000  163.455000 ;
      RECT -36.655000  164.645000 -35.375000  165.925000 ;
      RECT -34.600000 -180.935000 -33.320000 -179.655000 ;
      RECT -34.600000 -178.465000 -33.320000 -177.185000 ;
      RECT -34.600000 -175.395000 -33.320000 -174.115000 ;
      RECT -34.600000 -172.925000 -33.320000 -171.645000 ;
      RECT -34.600000 -150.915000 -33.320000 -149.635000 ;
      RECT -34.600000 -148.445000 -33.320000 -147.165000 ;
      RECT -34.600000 -145.375000 -33.320000 -144.095000 ;
      RECT -34.600000 -142.905000 -33.320000 -141.625000 ;
      RECT -34.035000  126.615000 -32.755000  127.895000 ;
      RECT -34.035000  129.085000 -32.755000  130.365000 ;
      RECT -34.035000  132.155000 -32.755000  133.435000 ;
      RECT -34.035000  134.625000 -32.755000  135.905000 ;
      RECT -34.035000  156.635000 -32.755000  157.915000 ;
      RECT -34.035000  159.105000 -32.755000  160.385000 ;
      RECT -34.035000  162.175000 -32.755000  163.455000 ;
      RECT -34.035000  164.645000 -32.755000  165.925000 ;
      RECT -31.830000 -180.935000 -30.550000 -179.655000 ;
      RECT -31.830000 -178.465000 -30.550000 -177.185000 ;
      RECT -31.830000 -175.395000 -30.550000 -174.115000 ;
      RECT -31.830000 -172.925000 -30.550000 -171.645000 ;
      RECT -31.830000 -150.915000 -30.550000 -149.635000 ;
      RECT -31.830000 -148.445000 -30.550000 -147.165000 ;
      RECT -31.830000 -145.375000 -30.550000 -144.095000 ;
      RECT -31.830000 -142.905000 -30.550000 -141.625000 ;
      RECT -31.265000  126.615000 -29.985000  127.895000 ;
      RECT -31.265000  129.085000 -29.985000  130.365000 ;
      RECT -31.265000  132.155000 -29.985000  133.435000 ;
      RECT -31.265000  134.625000 -29.985000  135.905000 ;
      RECT -31.265000  156.635000 -29.985000  157.915000 ;
      RECT -31.265000  159.105000 -29.985000  160.385000 ;
      RECT -31.265000  162.175000 -29.985000  163.455000 ;
      RECT -31.265000  164.645000 -29.985000  165.925000 ;
      RECT -29.060000 -180.935000 -27.780000 -179.655000 ;
      RECT -29.060000 -178.465000 -27.780000 -177.185000 ;
      RECT -29.060000 -175.395000 -27.780000 -174.115000 ;
      RECT -29.060000 -172.925000 -27.780000 -171.645000 ;
      RECT -29.060000 -150.915000 -27.780000 -149.635000 ;
      RECT -29.060000 -148.445000 -27.780000 -147.165000 ;
      RECT -29.060000 -145.375000 -27.780000 -144.095000 ;
      RECT -29.060000 -142.905000 -27.780000 -141.625000 ;
      RECT -28.495000  126.615000 -27.215000  127.895000 ;
      RECT -28.495000  129.085000 -27.215000  130.365000 ;
      RECT -28.495000  132.155000 -27.215000  133.435000 ;
      RECT -28.495000  134.625000 -27.215000  135.905000 ;
      RECT -28.495000  156.635000 -27.215000  157.915000 ;
      RECT -28.495000  159.105000 -27.215000  160.385000 ;
      RECT -28.495000  162.175000 -27.215000  163.455000 ;
      RECT -28.495000  164.645000 -27.215000  165.925000 ;
      RECT -26.440000 -180.935000 -25.160000 -179.655000 ;
      RECT -26.440000 -178.465000 -25.160000 -177.185000 ;
      RECT -26.440000 -175.395000 -25.160000 -174.115000 ;
      RECT -26.440000 -172.925000 -25.160000 -171.645000 ;
      RECT -26.440000 -150.915000 -25.160000 -149.635000 ;
      RECT -26.440000 -148.445000 -25.160000 -147.165000 ;
      RECT -26.440000 -145.375000 -25.160000 -144.095000 ;
      RECT -26.440000 -142.905000 -25.160000 -141.625000 ;
      RECT -25.875000  126.615000 -24.595000  127.895000 ;
      RECT -25.875000  129.085000 -24.595000  130.365000 ;
      RECT -25.875000  132.155000 -24.595000  133.435000 ;
      RECT -25.875000  134.625000 -24.595000  135.905000 ;
      RECT -25.875000  156.635000 -24.595000  157.915000 ;
      RECT -25.875000  159.105000 -24.595000  160.385000 ;
      RECT -25.875000  162.175000 -24.595000  163.455000 ;
      RECT -25.875000  164.645000 -24.595000  165.925000 ;
      RECT -23.370000 -180.935000 -22.090000 -179.655000 ;
      RECT -23.370000 -178.465000 -22.090000 -177.185000 ;
      RECT -23.370000 -175.395000 -22.090000 -174.115000 ;
      RECT -23.370000 -172.925000 -22.090000 -171.645000 ;
      RECT -23.370000 -150.915000 -22.090000 -149.635000 ;
      RECT -23.370000 -148.445000 -22.090000 -147.165000 ;
      RECT -23.370000 -145.375000 -22.090000 -144.095000 ;
      RECT -23.370000 -142.905000 -22.090000 -141.625000 ;
      RECT -22.805000  126.615000 -21.525000  127.895000 ;
      RECT -22.805000  129.085000 -21.525000  130.365000 ;
      RECT -22.805000  132.155000 -21.525000  133.435000 ;
      RECT -22.805000  134.625000 -21.525000  135.905000 ;
      RECT -22.805000  156.635000 -21.525000  157.915000 ;
      RECT -22.805000  159.105000 -21.525000  160.385000 ;
      RECT -22.805000  162.175000 -21.525000  163.455000 ;
      RECT -22.805000  164.645000 -21.525000  165.925000 ;
      RECT -20.750000 -180.935000 -19.470000 -179.655000 ;
      RECT -20.750000 -178.465000 -19.470000 -177.185000 ;
      RECT -20.750000 -175.395000 -19.470000 -174.115000 ;
      RECT -20.750000 -172.925000 -19.470000 -171.645000 ;
      RECT -20.750000 -150.915000 -19.470000 -149.635000 ;
      RECT -20.750000 -148.445000 -19.470000 -147.165000 ;
      RECT -20.750000 -145.375000 -19.470000 -144.095000 ;
      RECT -20.750000 -142.905000 -19.470000 -141.625000 ;
      RECT -20.185000  126.615000 -18.905000  127.895000 ;
      RECT -20.185000  129.085000 -18.905000  130.365000 ;
      RECT -20.185000  132.155000 -18.905000  133.435000 ;
      RECT -20.185000  134.625000 -18.905000  135.905000 ;
      RECT -20.185000  156.635000 -18.905000  157.915000 ;
      RECT -20.185000  159.105000 -18.905000  160.385000 ;
      RECT -20.185000  162.175000 -18.905000  163.455000 ;
      RECT -20.185000  164.645000 -18.905000  165.925000 ;
      RECT -17.980000 -180.935000 -16.700000 -179.655000 ;
      RECT -17.980000 -178.465000 -16.700000 -177.185000 ;
      RECT -17.980000 -175.395000 -16.700000 -174.115000 ;
      RECT -17.980000 -172.925000 -16.700000 -171.645000 ;
      RECT -17.980000 -150.915000 -16.700000 -149.635000 ;
      RECT -17.980000 -148.445000 -16.700000 -147.165000 ;
      RECT -17.980000 -145.375000 -16.700000 -144.095000 ;
      RECT -17.980000 -142.905000 -16.700000 -141.625000 ;
      RECT -17.415000  126.615000 -16.135000  127.895000 ;
      RECT -17.415000  129.085000 -16.135000  130.365000 ;
      RECT -17.415000  132.155000 -16.135000  133.435000 ;
      RECT -17.415000  134.625000 -16.135000  135.905000 ;
      RECT -17.415000  156.635000 -16.135000  157.915000 ;
      RECT -17.415000  159.105000 -16.135000  160.385000 ;
      RECT -17.415000  162.175000 -16.135000  163.455000 ;
      RECT -17.415000  164.645000 -16.135000  165.925000 ;
      RECT -15.210000 -180.935000 -13.930000 -179.655000 ;
      RECT -15.210000 -178.465000 -13.930000 -177.185000 ;
      RECT -15.210000 -175.395000 -13.930000 -174.115000 ;
      RECT -15.210000 -172.925000 -13.930000 -171.645000 ;
      RECT -15.210000 -150.915000 -13.930000 -149.635000 ;
      RECT -15.210000 -148.445000 -13.930000 -147.165000 ;
      RECT -15.210000 -145.375000 -13.930000 -144.095000 ;
      RECT -15.210000 -142.905000 -13.930000 -141.625000 ;
      RECT -14.645000  126.615000 -13.365000  127.895000 ;
      RECT -14.645000  129.085000 -13.365000  130.365000 ;
      RECT -14.645000  132.155000 -13.365000  133.435000 ;
      RECT -14.645000  134.625000 -13.365000  135.905000 ;
      RECT -14.645000  156.635000 -13.365000  157.915000 ;
      RECT -14.645000  159.105000 -13.365000  160.385000 ;
      RECT -14.645000  162.175000 -13.365000  163.455000 ;
      RECT -14.645000  164.645000 -13.365000  165.925000 ;
      RECT -12.590000 -180.935000 -11.310000 -179.655000 ;
      RECT -12.590000 -178.465000 -11.310000 -177.185000 ;
      RECT -12.590000 -175.395000 -11.310000 -174.115000 ;
      RECT -12.590000 -172.925000 -11.310000 -171.645000 ;
      RECT -12.590000 -150.915000 -11.310000 -149.635000 ;
      RECT -12.590000 -148.445000 -11.310000 -147.165000 ;
      RECT -12.590000 -145.375000 -11.310000 -144.095000 ;
      RECT -12.590000 -142.905000 -11.310000 -141.625000 ;
      RECT -12.025000  126.615000 -10.745000  127.895000 ;
      RECT -12.025000  129.085000 -10.745000  130.365000 ;
      RECT -12.025000  132.155000 -10.745000  133.435000 ;
      RECT -12.025000  134.625000 -10.745000  135.905000 ;
      RECT -12.025000  156.635000 -10.745000  157.915000 ;
      RECT -12.025000  159.105000 -10.745000  160.385000 ;
      RECT -12.025000  162.175000 -10.745000  163.455000 ;
      RECT -12.025000  164.645000 -10.745000  165.925000 ;
      RECT  11.965000 -165.920000  13.245000 -164.640000 ;
      RECT  11.965000 -163.450000  13.245000 -162.170000 ;
      RECT  11.965000 -160.380000  13.245000 -159.100000 ;
      RECT  11.965000 -157.910000  13.245000 -156.630000 ;
      RECT  11.965000 -135.910000  13.245000 -134.630000 ;
      RECT  11.965000 -133.440000  13.245000 -132.160000 ;
      RECT  11.965000 -130.370000  13.245000 -129.090000 ;
      RECT  11.965000 -127.900000  13.245000 -126.620000 ;
      RECT  12.520000  111.605000  13.800000  112.885000 ;
      RECT  12.520000  114.075000  13.800000  115.355000 ;
      RECT  12.520000  117.145000  13.800000  118.425000 ;
      RECT  12.520000  119.615000  13.800000  120.895000 ;
      RECT  12.520000  141.625000  13.800000  142.905000 ;
      RECT  12.520000  144.095000  13.800000  145.375000 ;
      RECT  12.520000  147.165000  13.800000  148.445000 ;
      RECT  12.520000  149.635000  13.800000  150.915000 ;
      RECT  14.585000 -165.920000  15.865000 -164.640000 ;
      RECT  14.585000 -163.450000  15.865000 -162.170000 ;
      RECT  14.585000 -160.380000  15.865000 -159.100000 ;
      RECT  14.585000 -157.910000  15.865000 -156.630000 ;
      RECT  14.585000 -135.910000  15.865000 -134.630000 ;
      RECT  14.585000 -133.440000  15.865000 -132.160000 ;
      RECT  14.585000 -130.370000  15.865000 -129.090000 ;
      RECT  14.585000 -127.900000  15.865000 -126.620000 ;
      RECT  15.140000  111.605000  16.420000  112.885000 ;
      RECT  15.140000  114.075000  16.420000  115.355000 ;
      RECT  15.140000  117.145000  16.420000  118.425000 ;
      RECT  15.140000  119.615000  16.420000  120.895000 ;
      RECT  15.140000  141.625000  16.420000  142.905000 ;
      RECT  15.140000  144.095000  16.420000  145.375000 ;
      RECT  15.140000  147.165000  16.420000  148.445000 ;
      RECT  15.140000  149.635000  16.420000  150.915000 ;
      RECT  17.355000 -165.920000  18.635000 -164.640000 ;
      RECT  17.355000 -163.450000  18.635000 -162.170000 ;
      RECT  17.355000 -160.380000  18.635000 -159.100000 ;
      RECT  17.355000 -157.910000  18.635000 -156.630000 ;
      RECT  17.355000 -135.910000  18.635000 -134.630000 ;
      RECT  17.355000 -133.440000  18.635000 -132.160000 ;
      RECT  17.355000 -130.370000  18.635000 -129.090000 ;
      RECT  17.355000 -127.900000  18.635000 -126.620000 ;
      RECT  17.910000  111.605000  19.190000  112.885000 ;
      RECT  17.910000  114.075000  19.190000  115.355000 ;
      RECT  17.910000  117.145000  19.190000  118.425000 ;
      RECT  17.910000  119.615000  19.190000  120.895000 ;
      RECT  17.910000  141.625000  19.190000  142.905000 ;
      RECT  17.910000  144.095000  19.190000  145.375000 ;
      RECT  17.910000  147.165000  19.190000  148.445000 ;
      RECT  17.910000  149.635000  19.190000  150.915000 ;
      RECT  20.125000 -165.920000  21.405000 -164.640000 ;
      RECT  20.125000 -163.450000  21.405000 -162.170000 ;
      RECT  20.125000 -160.380000  21.405000 -159.100000 ;
      RECT  20.125000 -157.910000  21.405000 -156.630000 ;
      RECT  20.125000 -135.910000  21.405000 -134.630000 ;
      RECT  20.125000 -133.440000  21.405000 -132.160000 ;
      RECT  20.125000 -130.370000  21.405000 -129.090000 ;
      RECT  20.125000 -127.900000  21.405000 -126.620000 ;
      RECT  20.680000  111.605000  21.960000  112.885000 ;
      RECT  20.680000  114.075000  21.960000  115.355000 ;
      RECT  20.680000  117.145000  21.960000  118.425000 ;
      RECT  20.680000  119.615000  21.960000  120.895000 ;
      RECT  20.680000  141.625000  21.960000  142.905000 ;
      RECT  20.680000  144.095000  21.960000  145.375000 ;
      RECT  20.680000  147.165000  21.960000  148.445000 ;
      RECT  20.680000  149.635000  21.960000  150.915000 ;
      RECT  22.745000 -165.920000  24.025000 -164.640000 ;
      RECT  22.745000 -163.450000  24.025000 -162.170000 ;
      RECT  22.745000 -160.380000  24.025000 -159.100000 ;
      RECT  22.745000 -157.910000  24.025000 -156.630000 ;
      RECT  22.745000 -135.910000  24.025000 -134.630000 ;
      RECT  22.745000 -133.440000  24.025000 -132.160000 ;
      RECT  22.745000 -130.370000  24.025000 -129.090000 ;
      RECT  22.745000 -127.900000  24.025000 -126.620000 ;
      RECT  23.300000  111.605000  24.580000  112.885000 ;
      RECT  23.300000  114.075000  24.580000  115.355000 ;
      RECT  23.300000  117.145000  24.580000  118.425000 ;
      RECT  23.300000  119.615000  24.580000  120.895000 ;
      RECT  23.300000  141.625000  24.580000  142.905000 ;
      RECT  23.300000  144.095000  24.580000  145.375000 ;
      RECT  23.300000  147.165000  24.580000  148.445000 ;
      RECT  23.300000  149.635000  24.580000  150.915000 ;
      RECT  25.815000 -165.920000  27.095000 -164.640000 ;
      RECT  25.815000 -163.450000  27.095000 -162.170000 ;
      RECT  25.815000 -160.380000  27.095000 -159.100000 ;
      RECT  25.815000 -157.910000  27.095000 -156.630000 ;
      RECT  25.815000 -135.910000  27.095000 -134.630000 ;
      RECT  25.815000 -133.440000  27.095000 -132.160000 ;
      RECT  25.815000 -130.370000  27.095000 -129.090000 ;
      RECT  25.815000 -127.900000  27.095000 -126.620000 ;
      RECT  26.370000  111.605000  27.650000  112.885000 ;
      RECT  26.370000  114.075000  27.650000  115.355000 ;
      RECT  26.370000  117.145000  27.650000  118.425000 ;
      RECT  26.370000  119.615000  27.650000  120.895000 ;
      RECT  26.370000  141.625000  27.650000  142.905000 ;
      RECT  26.370000  144.095000  27.650000  145.375000 ;
      RECT  26.370000  147.165000  27.650000  148.445000 ;
      RECT  26.370000  149.635000  27.650000  150.915000 ;
      RECT  28.435000 -165.920000  29.715000 -164.640000 ;
      RECT  28.435000 -163.450000  29.715000 -162.170000 ;
      RECT  28.435000 -160.380000  29.715000 -159.100000 ;
      RECT  28.435000 -157.910000  29.715000 -156.630000 ;
      RECT  28.435000 -135.910000  29.715000 -134.630000 ;
      RECT  28.435000 -133.440000  29.715000 -132.160000 ;
      RECT  28.435000 -130.370000  29.715000 -129.090000 ;
      RECT  28.435000 -127.900000  29.715000 -126.620000 ;
      RECT  28.990000  111.605000  30.270000  112.885000 ;
      RECT  28.990000  114.075000  30.270000  115.355000 ;
      RECT  28.990000  117.145000  30.270000  118.425000 ;
      RECT  28.990000  119.615000  30.270000  120.895000 ;
      RECT  28.990000  141.625000  30.270000  142.905000 ;
      RECT  28.990000  144.095000  30.270000  145.375000 ;
      RECT  28.990000  147.165000  30.270000  148.445000 ;
      RECT  28.990000  149.635000  30.270000  150.915000 ;
      RECT  31.205000 -165.920000  32.485000 -164.640000 ;
      RECT  31.205000 -163.450000  32.485000 -162.170000 ;
      RECT  31.205000 -160.380000  32.485000 -159.100000 ;
      RECT  31.205000 -157.910000  32.485000 -156.630000 ;
      RECT  31.205000 -135.910000  32.485000 -134.630000 ;
      RECT  31.205000 -133.440000  32.485000 -132.160000 ;
      RECT  31.205000 -130.370000  32.485000 -129.090000 ;
      RECT  31.205000 -127.900000  32.485000 -126.620000 ;
      RECT  31.760000  111.605000  33.040000  112.885000 ;
      RECT  31.760000  114.075000  33.040000  115.355000 ;
      RECT  31.760000  117.145000  33.040000  118.425000 ;
      RECT  31.760000  119.615000  33.040000  120.895000 ;
      RECT  31.760000  141.625000  33.040000  142.905000 ;
      RECT  31.760000  144.095000  33.040000  145.375000 ;
      RECT  31.760000  147.165000  33.040000  148.445000 ;
      RECT  31.760000  149.635000  33.040000  150.915000 ;
      RECT  33.975000 -165.920000  35.255000 -164.640000 ;
      RECT  33.975000 -163.450000  35.255000 -162.170000 ;
      RECT  33.975000 -160.380000  35.255000 -159.100000 ;
      RECT  33.975000 -157.910000  35.255000 -156.630000 ;
      RECT  33.975000 -135.910000  35.255000 -134.630000 ;
      RECT  33.975000 -133.440000  35.255000 -132.160000 ;
      RECT  33.975000 -130.370000  35.255000 -129.090000 ;
      RECT  33.975000 -127.900000  35.255000 -126.620000 ;
      RECT  34.530000  111.605000  35.810000  112.885000 ;
      RECT  34.530000  114.075000  35.810000  115.355000 ;
      RECT  34.530000  117.145000  35.810000  118.425000 ;
      RECT  34.530000  119.615000  35.810000  120.895000 ;
      RECT  34.530000  141.625000  35.810000  142.905000 ;
      RECT  34.530000  144.095000  35.810000  145.375000 ;
      RECT  34.530000  147.165000  35.810000  148.445000 ;
      RECT  34.530000  149.635000  35.810000  150.915000 ;
      RECT  36.595000 -165.920000  37.875000 -164.640000 ;
      RECT  36.595000 -163.450000  37.875000 -162.170000 ;
      RECT  36.595000 -160.380000  37.875000 -159.100000 ;
      RECT  36.595000 -157.910000  37.875000 -156.630000 ;
      RECT  36.595000 -135.910000  37.875000 -134.630000 ;
      RECT  36.595000 -133.440000  37.875000 -132.160000 ;
      RECT  36.595000 -130.370000  37.875000 -129.090000 ;
      RECT  36.595000 -127.900000  37.875000 -126.620000 ;
      RECT  37.150000  111.605000  38.430000  112.885000 ;
      RECT  37.150000  114.075000  38.430000  115.355000 ;
      RECT  37.150000  117.145000  38.430000  118.425000 ;
      RECT  37.150000  119.615000  38.430000  120.895000 ;
      RECT  37.150000  141.625000  38.430000  142.905000 ;
      RECT  37.150000  144.095000  38.430000  145.375000 ;
      RECT  37.150000  147.165000  38.430000  148.445000 ;
      RECT  37.150000  149.635000  38.430000  150.915000 ;
      RECT  97.760000   -4.645000  99.040000   -3.365000 ;
      RECT  97.760000   -2.175000  99.040000   -0.895000 ;
      RECT  97.760000    0.895000  99.040000    2.175000 ;
      RECT  97.760000    3.365000  99.040000    4.645000 ;
      RECT 100.380000   -4.645000 101.660000   -3.365000 ;
      RECT 100.380000   -2.175000 101.660000   -0.895000 ;
      RECT 100.380000    0.895000 101.660000    2.175000 ;
      RECT 100.380000    3.365000 101.660000    4.645000 ;
      RECT 103.150000   -4.645000 104.430000   -3.365000 ;
      RECT 103.150000   -2.175000 104.430000   -0.895000 ;
      RECT 103.150000    0.895000 104.430000    2.175000 ;
      RECT 103.150000    3.365000 104.430000    4.645000 ;
  END
END sky130_fd_pr__rf_test_coil3
END LIBRARY
