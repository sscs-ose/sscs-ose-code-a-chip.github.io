# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.350000 BY  4.900000 ;
  PIN BULK
    ANTENNADIFFAREA  3.913000 ;
    ANTENNAGATEAREA  0.903000 ;
    PORT
      LAYER li1 ;
        RECT 0.205000 0.925000 0.800000 3.975000 ;
        RECT 0.600000 0.455000 0.930000 0.785000 ;
        RECT 0.600000 0.785000 0.800000 0.925000 ;
        RECT 0.600000 3.975000 0.800000 4.115000 ;
        RECT 0.600000 4.115000 0.930000 4.445000 ;
        RECT 2.420000 0.455000 2.750000 0.785000 ;
        RECT 2.420000 4.115000 2.750000 4.445000 ;
        RECT 2.550000 0.785000 2.750000 0.925000 ;
        RECT 2.550000 0.925000 3.145000 3.975000 ;
        RECT 2.550000 3.975000 2.750000 4.115000 ;
      LAYER mcon ;
        RECT 0.300000 1.105000 0.470000 1.275000 ;
        RECT 0.300000 1.465000 0.470000 1.635000 ;
        RECT 0.300000 1.825000 0.470000 1.995000 ;
        RECT 0.300000 2.185000 0.470000 2.355000 ;
        RECT 0.300000 2.545000 0.470000 2.715000 ;
        RECT 0.300000 2.905000 0.470000 3.075000 ;
        RECT 0.300000 3.265000 0.470000 3.435000 ;
        RECT 0.300000 3.625000 0.470000 3.795000 ;
        RECT 2.880000 1.105000 3.050000 1.275000 ;
        RECT 2.880000 1.465000 3.050000 1.635000 ;
        RECT 2.880000 1.825000 3.050000 1.995000 ;
        RECT 2.880000 2.185000 3.050000 2.355000 ;
        RECT 2.880000 2.545000 3.050000 2.715000 ;
        RECT 2.880000 2.905000 3.050000 3.075000 ;
        RECT 2.880000 3.265000 3.050000 3.435000 ;
        RECT 2.880000 3.625000 3.050000 3.795000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.205000 1.045000 0.500000 3.855000 ;
        RECT 2.850000 1.045000 3.145000 3.855000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  0.842800 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.575000 3.280000 3.855000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.505000 ;
    PORT
      LAYER li1 ;
        RECT 1.240000 0.000000 2.110000 0.695000 ;
        RECT 1.240000 4.205000 2.110000 4.900000 ;
      LAYER mcon ;
        RECT 1.380000 0.095000 1.550000 0.265000 ;
        RECT 1.380000 0.455000 1.550000 0.625000 ;
        RECT 1.380000 4.275000 1.550000 4.445000 ;
        RECT 1.380000 4.635000 1.550000 4.805000 ;
        RECT 1.800000 0.095000 1.970000 0.265000 ;
        RECT 1.800000 0.455000 1.970000 0.625000 ;
        RECT 1.800000 4.275000 1.970000 4.445000 ;
        RECT 1.800000 4.635000 1.970000 4.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.250000 0.000000 2.100000 0.685000 ;
        RECT 1.250000 4.215000 2.100000 4.900000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.685600 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.045000 3.280000 2.325000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 1.060000 0.925000 1.230000 3.975000 ;
      RECT 1.590000 0.925000 1.760000 3.975000 ;
      RECT 2.120000 0.925000 2.290000 3.975000 ;
    LAYER mcon ;
      RECT 1.060000 1.105000 1.230000 1.275000 ;
      RECT 1.060000 1.465000 1.230000 1.635000 ;
      RECT 1.060000 1.825000 1.230000 1.995000 ;
      RECT 1.060000 2.185000 1.230000 2.355000 ;
      RECT 1.060000 2.545000 1.230000 2.715000 ;
      RECT 1.060000 2.905000 1.230000 3.075000 ;
      RECT 1.060000 3.265000 1.230000 3.435000 ;
      RECT 1.060000 3.625000 1.230000 3.795000 ;
      RECT 1.590000 1.105000 1.760000 1.275000 ;
      RECT 1.590000 1.465000 1.760000 1.635000 ;
      RECT 1.590000 1.825000 1.760000 1.995000 ;
      RECT 1.590000 2.185000 1.760000 2.355000 ;
      RECT 1.590000 2.545000 1.760000 2.715000 ;
      RECT 1.590000 2.905000 1.760000 3.075000 ;
      RECT 1.590000 3.265000 1.760000 3.435000 ;
      RECT 1.590000 3.625000 1.760000 3.795000 ;
      RECT 2.120000 1.105000 2.290000 1.275000 ;
      RECT 2.120000 1.465000 2.290000 1.635000 ;
      RECT 2.120000 1.825000 2.290000 1.995000 ;
      RECT 2.120000 2.185000 2.290000 2.355000 ;
      RECT 2.120000 2.545000 2.290000 2.715000 ;
      RECT 2.120000 2.905000 2.290000 3.075000 ;
      RECT 2.120000 3.265000 2.290000 3.435000 ;
      RECT 2.120000 3.625000 2.290000 3.795000 ;
    LAYER met1 ;
      RECT 1.015000 1.045000 1.275000 3.855000 ;
      RECT 1.545000 1.045000 1.805000 3.855000 ;
      RECT 2.075000 1.045000 2.335000 3.855000 ;
    LAYER via ;
      RECT 1.015000 1.075000 1.275000 1.335000 ;
      RECT 1.015000 1.395000 1.275000 1.655000 ;
      RECT 1.015000 1.715000 1.275000 1.975000 ;
      RECT 1.015000 2.035000 1.275000 2.295000 ;
      RECT 1.545000 2.605000 1.805000 2.865000 ;
      RECT 1.545000 2.925000 1.805000 3.185000 ;
      RECT 1.545000 3.245000 1.805000 3.505000 ;
      RECT 1.545000 3.565000 1.805000 3.825000 ;
      RECT 2.075000 1.075000 2.335000 1.335000 ;
      RECT 2.075000 1.395000 2.335000 1.655000 ;
      RECT 2.075000 1.715000 2.335000 1.975000 ;
      RECT 2.075000 2.035000 2.335000 2.295000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25
END LIBRARY
