txt.md
