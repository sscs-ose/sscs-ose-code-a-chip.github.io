# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4_top
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4_top ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.430000 BY  8.850000 ;
  PIN C0
    PORT
      LAYER met3 ;
        RECT 0.000000 0.000000 8.430000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 4.260000 ;
        RECT 0.000000 4.260000 8.430000 4.590000 ;
        RECT 0.000000 4.590000 0.330000 8.520000 ;
        RECT 0.000000 8.520000 8.430000 8.850000 ;
        RECT 1.230000 0.330000 1.530000 1.830000 ;
        RECT 1.230000 2.760000 1.530000 4.260000 ;
        RECT 1.230000 4.590000 1.530000 6.090000 ;
        RECT 1.230000 7.020000 1.530000 8.520000 ;
        RECT 2.850000 0.330000 3.150000 1.830000 ;
        RECT 2.850000 2.760000 3.150000 4.260000 ;
        RECT 2.850000 4.590000 3.150000 6.090000 ;
        RECT 2.850000 7.020000 3.150000 8.520000 ;
        RECT 4.050000 0.330000 4.380000 4.260000 ;
        RECT 4.050000 4.590000 4.380000 8.520000 ;
        RECT 5.280000 0.330000 5.580000 1.830000 ;
        RECT 5.280000 2.760000 5.580000 4.260000 ;
        RECT 5.280000 4.590000 5.580000 6.090000 ;
        RECT 5.280000 7.020000 5.580000 8.520000 ;
        RECT 6.900000 0.330000 7.200000 1.830000 ;
        RECT 6.900000 2.760000 7.200000 4.260000 ;
        RECT 6.900000 4.590000 7.200000 6.090000 ;
        RECT 6.900000 7.020000 7.200000 8.520000 ;
        RECT 8.100000 0.330000 8.430000 4.260000 ;
        RECT 8.100000 4.590000 8.430000 8.520000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT 0.630000 0.630000 0.930000 2.130000 ;
        RECT 0.630000 2.130000 3.750000 2.460000 ;
        RECT 0.630000 2.460000 0.930000 3.960000 ;
        RECT 0.630000 4.890000 0.930000 6.390000 ;
        RECT 0.630000 6.390000 3.750000 6.720000 ;
        RECT 0.630000 6.720000 0.930000 8.220000 ;
        RECT 2.025000 0.630000 2.355000 2.130000 ;
        RECT 2.025000 2.460000 2.355000 3.960000 ;
        RECT 2.025000 4.890000 2.355000 6.390000 ;
        RECT 2.025000 6.720000 2.355000 8.220000 ;
        RECT 3.450000 0.630000 3.750000 2.130000 ;
        RECT 3.450000 2.460000 3.750000 3.960000 ;
        RECT 3.450000 4.890000 3.750000 6.390000 ;
        RECT 3.450000 6.720000 3.750000 8.220000 ;
        RECT 4.680000 0.630000 4.980000 2.130000 ;
        RECT 4.680000 2.130000 7.800000 2.460000 ;
        RECT 4.680000 2.460000 4.980000 3.960000 ;
        RECT 4.680000 4.890000 4.980000 6.390000 ;
        RECT 4.680000 6.390000 7.800000 6.720000 ;
        RECT 4.680000 6.720000 4.980000 8.220000 ;
        RECT 6.075000 0.630000 6.405000 2.130000 ;
        RECT 6.075000 2.460000 6.405000 3.960000 ;
        RECT 6.075000 4.890000 6.405000 6.390000 ;
        RECT 6.075000 6.720000 6.405000 8.220000 ;
        RECT 7.500000 0.630000 7.800000 2.130000 ;
        RECT 7.500000 2.460000 7.800000 3.960000 ;
        RECT 7.500000 4.890000 7.800000 6.390000 ;
        RECT 7.500000 6.720000 7.800000 8.220000 ;
    END
  END C1
  PIN M5
    PORT
      LAYER met5 ;
        RECT 0.000000 0.000000 8.430000 8.850000 ;
    END
  END M5
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 5.895000 6.345000 5.945000 6.395000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 8.430000 8.850000 ;
    LAYER mcon ;
      RECT 0.080000 0.410000 0.250000 0.580000 ;
      RECT 0.080000 0.770000 0.250000 0.940000 ;
      RECT 0.080000 1.130000 0.250000 1.300000 ;
      RECT 0.080000 1.490000 0.250000 1.660000 ;
      RECT 0.080000 1.850000 0.250000 2.020000 ;
      RECT 0.080000 2.210000 0.250000 2.380000 ;
      RECT 0.080000 2.570000 0.250000 2.740000 ;
      RECT 0.080000 2.930000 0.250000 3.100000 ;
      RECT 0.080000 3.290000 0.250000 3.460000 ;
      RECT 0.080000 3.650000 0.250000 3.820000 ;
      RECT 0.080000 4.010000 0.250000 4.180000 ;
      RECT 0.080000 4.670000 0.250000 4.840000 ;
      RECT 0.080000 5.030000 0.250000 5.200000 ;
      RECT 0.080000 5.390000 0.250000 5.560000 ;
      RECT 0.080000 5.750000 0.250000 5.920000 ;
      RECT 0.080000 6.110000 0.250000 6.280000 ;
      RECT 0.080000 6.470000 0.250000 6.640000 ;
      RECT 0.080000 6.830000 0.250000 7.000000 ;
      RECT 0.080000 7.190000 0.250000 7.360000 ;
      RECT 0.080000 7.550000 0.250000 7.720000 ;
      RECT 0.080000 7.910000 0.250000 8.080000 ;
      RECT 0.080000 8.270000 0.250000 8.440000 ;
      RECT 0.485000 0.080000 0.655000 0.250000 ;
      RECT 0.485000 4.340000 0.655000 4.510000 ;
      RECT 0.485000 8.600000 0.655000 8.770000 ;
      RECT 0.845000 0.080000 1.015000 0.250000 ;
      RECT 0.845000 4.340000 1.015000 4.510000 ;
      RECT 0.845000 8.600000 1.015000 8.770000 ;
      RECT 1.205000 0.080000 1.375000 0.250000 ;
      RECT 1.205000 4.340000 1.375000 4.510000 ;
      RECT 1.205000 8.600000 1.375000 8.770000 ;
      RECT 1.565000 0.080000 1.735000 0.250000 ;
      RECT 1.565000 4.340000 1.735000 4.510000 ;
      RECT 1.565000 8.600000 1.735000 8.770000 ;
      RECT 1.925000 0.080000 2.095000 0.250000 ;
      RECT 1.925000 4.340000 2.095000 4.510000 ;
      RECT 1.925000 8.600000 2.095000 8.770000 ;
      RECT 2.285000 0.080000 2.455000 0.250000 ;
      RECT 2.285000 4.340000 2.455000 4.510000 ;
      RECT 2.285000 8.600000 2.455000 8.770000 ;
      RECT 2.645000 0.080000 2.815000 0.250000 ;
      RECT 2.645000 4.340000 2.815000 4.510000 ;
      RECT 2.645000 8.600000 2.815000 8.770000 ;
      RECT 3.005000 0.080000 3.175000 0.250000 ;
      RECT 3.005000 4.340000 3.175000 4.510000 ;
      RECT 3.005000 8.600000 3.175000 8.770000 ;
      RECT 3.365000 0.080000 3.535000 0.250000 ;
      RECT 3.365000 4.340000 3.535000 4.510000 ;
      RECT 3.365000 8.600000 3.535000 8.770000 ;
      RECT 3.725000 0.080000 3.895000 0.250000 ;
      RECT 3.725000 4.340000 3.895000 4.510000 ;
      RECT 3.725000 8.600000 3.895000 8.770000 ;
      RECT 4.130000 0.410000 4.300000 0.580000 ;
      RECT 4.130000 0.770000 4.300000 0.940000 ;
      RECT 4.130000 1.130000 4.300000 1.300000 ;
      RECT 4.130000 1.490000 4.300000 1.660000 ;
      RECT 4.130000 1.850000 4.300000 2.020000 ;
      RECT 4.130000 2.210000 4.300000 2.380000 ;
      RECT 4.130000 2.570000 4.300000 2.740000 ;
      RECT 4.130000 2.930000 4.300000 3.100000 ;
      RECT 4.130000 3.290000 4.300000 3.460000 ;
      RECT 4.130000 3.650000 4.300000 3.820000 ;
      RECT 4.130000 4.010000 4.300000 4.180000 ;
      RECT 4.130000 4.670000 4.300000 4.840000 ;
      RECT 4.130000 5.030000 4.300000 5.200000 ;
      RECT 4.130000 5.390000 4.300000 5.560000 ;
      RECT 4.130000 5.750000 4.300000 5.920000 ;
      RECT 4.130000 6.110000 4.300000 6.280000 ;
      RECT 4.130000 6.470000 4.300000 6.640000 ;
      RECT 4.130000 6.830000 4.300000 7.000000 ;
      RECT 4.130000 7.190000 4.300000 7.360000 ;
      RECT 4.130000 7.550000 4.300000 7.720000 ;
      RECT 4.130000 7.910000 4.300000 8.080000 ;
      RECT 4.130000 8.270000 4.300000 8.440000 ;
      RECT 4.535000 0.080000 4.705000 0.250000 ;
      RECT 4.535000 4.340000 4.705000 4.510000 ;
      RECT 4.535000 8.600000 4.705000 8.770000 ;
      RECT 4.895000 0.080000 5.065000 0.250000 ;
      RECT 4.895000 4.340000 5.065000 4.510000 ;
      RECT 4.895000 8.600000 5.065000 8.770000 ;
      RECT 5.255000 0.080000 5.425000 0.250000 ;
      RECT 5.255000 4.340000 5.425000 4.510000 ;
      RECT 5.255000 8.600000 5.425000 8.770000 ;
      RECT 5.615000 0.080000 5.785000 0.250000 ;
      RECT 5.615000 4.340000 5.785000 4.510000 ;
      RECT 5.615000 8.600000 5.785000 8.770000 ;
      RECT 5.975000 0.080000 6.145000 0.250000 ;
      RECT 5.975000 4.340000 6.145000 4.510000 ;
      RECT 5.975000 8.600000 6.145000 8.770000 ;
      RECT 6.335000 0.080000 6.505000 0.250000 ;
      RECT 6.335000 4.340000 6.505000 4.510000 ;
      RECT 6.335000 8.600000 6.505000 8.770000 ;
      RECT 6.695000 0.080000 6.865000 0.250000 ;
      RECT 6.695000 4.340000 6.865000 4.510000 ;
      RECT 6.695000 8.600000 6.865000 8.770000 ;
      RECT 7.055000 0.080000 7.225000 0.250000 ;
      RECT 7.055000 4.340000 7.225000 4.510000 ;
      RECT 7.055000 8.600000 7.225000 8.770000 ;
      RECT 7.415000 0.080000 7.585000 0.250000 ;
      RECT 7.415000 4.340000 7.585000 4.510000 ;
      RECT 7.415000 8.600000 7.585000 8.770000 ;
      RECT 7.775000 0.080000 7.945000 0.250000 ;
      RECT 7.775000 4.340000 7.945000 4.510000 ;
      RECT 7.775000 8.600000 7.945000 8.770000 ;
      RECT 8.180000 0.410000 8.350000 0.580000 ;
      RECT 8.180000 0.770000 8.350000 0.940000 ;
      RECT 8.180000 1.130000 8.350000 1.300000 ;
      RECT 8.180000 1.490000 8.350000 1.660000 ;
      RECT 8.180000 1.850000 8.350000 2.020000 ;
      RECT 8.180000 2.210000 8.350000 2.380000 ;
      RECT 8.180000 2.570000 8.350000 2.740000 ;
      RECT 8.180000 2.930000 8.350000 3.100000 ;
      RECT 8.180000 3.290000 8.350000 3.460000 ;
      RECT 8.180000 3.650000 8.350000 3.820000 ;
      RECT 8.180000 4.010000 8.350000 4.180000 ;
      RECT 8.180000 4.670000 8.350000 4.840000 ;
      RECT 8.180000 5.030000 8.350000 5.200000 ;
      RECT 8.180000 5.390000 8.350000 5.560000 ;
      RECT 8.180000 5.750000 8.350000 5.920000 ;
      RECT 8.180000 6.110000 8.350000 6.280000 ;
      RECT 8.180000 6.470000 8.350000 6.640000 ;
      RECT 8.180000 6.830000 8.350000 7.000000 ;
      RECT 8.180000 7.190000 8.350000 7.360000 ;
      RECT 8.180000 7.550000 8.350000 7.720000 ;
      RECT 8.180000 7.910000 8.350000 8.080000 ;
      RECT 8.180000 8.270000 8.350000 8.440000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 8.430000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 4.260000 ;
      RECT 0.000000 4.260000 8.430000 4.590000 ;
      RECT 0.000000 4.590000 0.330000 8.520000 ;
      RECT 0.000000 8.520000 8.430000 8.850000 ;
      RECT 0.565000 0.470000 0.705000 2.135000 ;
      RECT 0.565000 2.135000 3.815000 2.455000 ;
      RECT 0.565000 2.455000 0.705000 4.120000 ;
      RECT 0.565000 4.730000 0.705000 6.395000 ;
      RECT 0.565000 6.395000 3.815000 6.715000 ;
      RECT 0.565000 6.715000 0.705000 8.380000 ;
      RECT 0.845000 0.330000 0.985000 1.995000 ;
      RECT 0.845000 2.595000 0.985000 4.260000 ;
      RECT 0.845000 4.590000 0.985000 6.255000 ;
      RECT 0.845000 6.855000 0.985000 8.520000 ;
      RECT 1.125000 0.470000 1.265000 2.135000 ;
      RECT 1.125000 2.455000 1.265000 4.120000 ;
      RECT 1.125000 4.730000 1.265000 6.395000 ;
      RECT 1.125000 6.715000 1.265000 8.380000 ;
      RECT 1.405000 0.330000 1.545000 1.995000 ;
      RECT 1.405000 2.595000 1.545000 4.260000 ;
      RECT 1.405000 4.590000 1.545000 6.255000 ;
      RECT 1.405000 6.855000 1.545000 8.520000 ;
      RECT 1.685000 0.470000 1.825000 2.135000 ;
      RECT 1.685000 2.455000 1.825000 4.120000 ;
      RECT 1.685000 4.730000 1.825000 6.395000 ;
      RECT 1.685000 6.715000 1.825000 8.380000 ;
      RECT 2.055000 0.470000 2.325000 2.135000 ;
      RECT 2.055000 2.455000 2.325000 4.120000 ;
      RECT 2.055000 4.730000 2.325000 6.395000 ;
      RECT 2.055000 6.715000 2.325000 8.380000 ;
      RECT 2.555000 0.470000 2.695000 2.135000 ;
      RECT 2.555000 2.455000 2.695000 4.120000 ;
      RECT 2.555000 4.730000 2.695000 6.395000 ;
      RECT 2.555000 6.715000 2.695000 8.380000 ;
      RECT 2.835000 0.330000 2.975000 1.995000 ;
      RECT 2.835000 2.595000 2.975000 4.260000 ;
      RECT 2.835000 4.590000 2.975000 6.255000 ;
      RECT 2.835000 6.855000 2.975000 8.520000 ;
      RECT 3.115000 0.470000 3.255000 2.135000 ;
      RECT 3.115000 2.455000 3.255000 4.120000 ;
      RECT 3.115000 4.730000 3.255000 6.395000 ;
      RECT 3.115000 6.715000 3.255000 8.380000 ;
      RECT 3.395000 0.330000 3.535000 1.995000 ;
      RECT 3.395000 2.595000 3.535000 4.260000 ;
      RECT 3.395000 4.590000 3.535000 6.255000 ;
      RECT 3.395000 6.855000 3.535000 8.520000 ;
      RECT 3.675000 0.470000 3.815000 2.135000 ;
      RECT 3.675000 2.455000 3.815000 4.120000 ;
      RECT 3.675000 4.730000 3.815000 6.395000 ;
      RECT 3.675000 6.715000 3.815000 8.380000 ;
      RECT 4.050000 0.330000 4.380000 4.260000 ;
      RECT 4.050000 4.590000 4.380000 8.520000 ;
      RECT 4.615000 0.470000 4.755000 2.135000 ;
      RECT 4.615000 2.135000 7.865000 2.455000 ;
      RECT 4.615000 2.455000 4.755000 4.120000 ;
      RECT 4.615000 4.730000 4.755000 6.395000 ;
      RECT 4.615000 6.395000 7.865000 6.715000 ;
      RECT 4.615000 6.715000 4.755000 8.380000 ;
      RECT 4.895000 0.330000 5.035000 1.995000 ;
      RECT 4.895000 2.595000 5.035000 4.260000 ;
      RECT 4.895000 4.590000 5.035000 6.255000 ;
      RECT 4.895000 6.855000 5.035000 8.520000 ;
      RECT 5.175000 0.470000 5.315000 2.135000 ;
      RECT 5.175000 2.455000 5.315000 4.120000 ;
      RECT 5.175000 4.730000 5.315000 6.395000 ;
      RECT 5.175000 6.715000 5.315000 8.380000 ;
      RECT 5.455000 0.330000 5.595000 1.995000 ;
      RECT 5.455000 2.595000 5.595000 4.260000 ;
      RECT 5.455000 4.590000 5.595000 6.255000 ;
      RECT 5.455000 6.855000 5.595000 8.520000 ;
      RECT 5.735000 0.470000 5.875000 2.135000 ;
      RECT 5.735000 2.455000 5.875000 4.120000 ;
      RECT 5.735000 4.730000 5.875000 6.395000 ;
      RECT 5.735000 6.715000 5.875000 8.380000 ;
      RECT 6.105000 0.470000 6.375000 2.135000 ;
      RECT 6.105000 2.455000 6.375000 4.120000 ;
      RECT 6.105000 4.730000 6.375000 6.395000 ;
      RECT 6.105000 6.715000 6.375000 8.380000 ;
      RECT 6.605000 0.470000 6.745000 2.135000 ;
      RECT 6.605000 2.455000 6.745000 4.120000 ;
      RECT 6.605000 4.730000 6.745000 6.395000 ;
      RECT 6.605000 6.715000 6.745000 8.380000 ;
      RECT 6.885000 0.330000 7.025000 1.995000 ;
      RECT 6.885000 2.595000 7.025000 4.260000 ;
      RECT 6.885000 4.590000 7.025000 6.255000 ;
      RECT 6.885000 6.855000 7.025000 8.520000 ;
      RECT 7.165000 0.470000 7.305000 2.135000 ;
      RECT 7.165000 2.455000 7.305000 4.120000 ;
      RECT 7.165000 4.730000 7.305000 6.395000 ;
      RECT 7.165000 6.715000 7.305000 8.380000 ;
      RECT 7.445000 0.330000 7.585000 1.995000 ;
      RECT 7.445000 2.595000 7.585000 4.260000 ;
      RECT 7.445000 4.590000 7.585000 6.255000 ;
      RECT 7.445000 6.855000 7.585000 8.520000 ;
      RECT 7.725000 0.470000 7.865000 2.135000 ;
      RECT 7.725000 2.455000 7.865000 4.120000 ;
      RECT 7.725000 4.730000 7.865000 6.395000 ;
      RECT 7.725000 6.715000 7.865000 8.380000 ;
      RECT 8.100000 0.330000 8.430000 4.260000 ;
      RECT 8.100000 4.590000 8.430000 8.520000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 1.915000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 0.750000 ;
      RECT 0.000000 0.750000 1.910000 0.890000 ;
      RECT 0.000000 0.890000 0.330000 1.310000 ;
      RECT 0.000000 1.310000 1.910000 1.450000 ;
      RECT 0.000000 1.450000 0.330000 1.870000 ;
      RECT 0.000000 1.870000 1.910000 2.010000 ;
      RECT 0.000000 2.010000 0.330000 2.020000 ;
      RECT 0.000000 2.160000 8.430000 2.430000 ;
      RECT 0.000000 2.570000 0.330000 2.580000 ;
      RECT 0.000000 2.580000 1.910000 2.720000 ;
      RECT 0.000000 2.720000 0.330000 3.140000 ;
      RECT 0.000000 3.140000 1.910000 3.280000 ;
      RECT 0.000000 3.280000 0.330000 3.700000 ;
      RECT 0.000000 3.700000 1.910000 3.840000 ;
      RECT 0.000000 3.840000 0.330000 4.260000 ;
      RECT 0.000000 4.260000 1.915000 4.590000 ;
      RECT 0.000000 4.590000 0.330000 5.010000 ;
      RECT 0.000000 5.010000 1.910000 5.150000 ;
      RECT 0.000000 5.150000 0.330000 5.570000 ;
      RECT 0.000000 5.570000 1.910000 5.710000 ;
      RECT 0.000000 5.710000 0.330000 6.130000 ;
      RECT 0.000000 6.130000 1.910000 6.270000 ;
      RECT 0.000000 6.270000 0.330000 6.280000 ;
      RECT 0.000000 6.420000 8.430000 6.690000 ;
      RECT 0.000000 6.830000 0.330000 6.840000 ;
      RECT 0.000000 6.840000 1.910000 6.980000 ;
      RECT 0.000000 6.980000 0.330000 7.400000 ;
      RECT 0.000000 7.400000 1.910000 7.540000 ;
      RECT 0.000000 7.540000 0.330000 7.960000 ;
      RECT 0.000000 7.960000 1.910000 8.100000 ;
      RECT 0.000000 8.100000 0.330000 8.520000 ;
      RECT 0.000000 8.520000 1.915000 8.850000 ;
      RECT 0.370000 2.155000 4.010000 2.160000 ;
      RECT 0.370000 2.430000 4.010000 2.435000 ;
      RECT 0.370000 6.415000 4.010000 6.420000 ;
      RECT 0.370000 6.690000 4.010000 6.695000 ;
      RECT 0.470000 0.470000 3.910000 0.610000 ;
      RECT 0.470000 1.030000 3.910000 1.170000 ;
      RECT 0.470000 1.590000 3.910000 1.730000 ;
      RECT 0.470000 2.860000 3.910000 3.000000 ;
      RECT 0.470000 3.420000 3.910000 3.560000 ;
      RECT 0.470000 3.980000 3.910000 4.120000 ;
      RECT 0.470000 4.730000 3.910000 4.870000 ;
      RECT 0.470000 5.290000 3.910000 5.430000 ;
      RECT 0.470000 5.850000 3.910000 5.990000 ;
      RECT 0.470000 7.120000 3.910000 7.260000 ;
      RECT 0.470000 7.680000 3.910000 7.820000 ;
      RECT 0.470000 8.240000 3.910000 8.380000 ;
      RECT 2.050000 0.610000 2.330000 1.030000 ;
      RECT 2.050000 1.170000 2.330000 1.590000 ;
      RECT 2.050000 1.730000 2.330000 2.155000 ;
      RECT 2.050000 2.435000 2.330000 2.860000 ;
      RECT 2.050000 3.000000 2.330000 3.420000 ;
      RECT 2.050000 3.560000 2.330000 3.980000 ;
      RECT 2.050000 4.870000 2.330000 5.290000 ;
      RECT 2.050000 5.430000 2.330000 5.850000 ;
      RECT 2.050000 5.990000 2.330000 6.415000 ;
      RECT 2.050000 6.695000 2.330000 7.120000 ;
      RECT 2.050000 7.260000 2.330000 7.680000 ;
      RECT 2.050000 7.820000 2.330000 8.240000 ;
      RECT 2.055000 0.000000 2.325000 0.470000 ;
      RECT 2.055000 4.120000 2.325000 4.730000 ;
      RECT 2.055000 8.380000 2.325000 8.850000 ;
      RECT 2.465000 0.000000 5.965000 0.330000 ;
      RECT 2.465000 4.260000 5.965000 4.590000 ;
      RECT 2.465000 8.520000 5.965000 8.850000 ;
      RECT 2.470000 0.750000 5.960000 0.890000 ;
      RECT 2.470000 1.310000 5.960000 1.450000 ;
      RECT 2.470000 1.870000 5.960000 2.010000 ;
      RECT 2.470000 2.580000 5.960000 2.720000 ;
      RECT 2.470000 3.140000 5.960000 3.280000 ;
      RECT 2.470000 3.700000 5.960000 3.840000 ;
      RECT 2.470000 5.010000 5.960000 5.150000 ;
      RECT 2.470000 5.570000 5.960000 5.710000 ;
      RECT 2.470000 6.130000 5.960000 6.270000 ;
      RECT 2.470000 6.840000 5.960000 6.980000 ;
      RECT 2.470000 7.400000 5.960000 7.540000 ;
      RECT 2.470000 7.960000 5.960000 8.100000 ;
      RECT 4.050000 0.330000 4.380000 0.750000 ;
      RECT 4.050000 0.890000 4.380000 1.310000 ;
      RECT 4.050000 1.450000 4.380000 1.870000 ;
      RECT 4.050000 2.010000 4.380000 2.020000 ;
      RECT 4.050000 2.570000 4.380000 2.580000 ;
      RECT 4.050000 2.720000 4.380000 3.140000 ;
      RECT 4.050000 3.280000 4.380000 3.700000 ;
      RECT 4.050000 3.840000 4.380000 4.260000 ;
      RECT 4.050000 4.590000 4.380000 5.010000 ;
      RECT 4.050000 5.150000 4.380000 5.570000 ;
      RECT 4.050000 5.710000 4.380000 6.130000 ;
      RECT 4.050000 6.270000 4.380000 6.280000 ;
      RECT 4.050000 6.830000 4.380000 6.840000 ;
      RECT 4.050000 6.980000 4.380000 7.400000 ;
      RECT 4.050000 7.540000 4.380000 7.960000 ;
      RECT 4.050000 8.100000 4.380000 8.520000 ;
      RECT 4.420000 2.155000 8.060000 2.160000 ;
      RECT 4.420000 2.430000 8.060000 2.435000 ;
      RECT 4.420000 6.415000 8.060000 6.420000 ;
      RECT 4.420000 6.690000 8.060000 6.695000 ;
      RECT 4.520000 0.470000 7.960000 0.610000 ;
      RECT 4.520000 1.030000 7.960000 1.170000 ;
      RECT 4.520000 1.590000 7.960000 1.730000 ;
      RECT 4.520000 2.860000 7.960000 3.000000 ;
      RECT 4.520000 3.420000 7.960000 3.560000 ;
      RECT 4.520000 3.980000 7.960000 4.120000 ;
      RECT 4.520000 4.730000 7.960000 4.870000 ;
      RECT 4.520000 5.290000 7.960000 5.430000 ;
      RECT 4.520000 5.850000 7.960000 5.990000 ;
      RECT 4.520000 7.120000 7.960000 7.260000 ;
      RECT 4.520000 7.680000 7.960000 7.820000 ;
      RECT 4.520000 8.240000 7.960000 8.380000 ;
      RECT 6.100000 0.610000 6.380000 1.030000 ;
      RECT 6.100000 1.170000 6.380000 1.590000 ;
      RECT 6.100000 1.730000 6.380000 2.155000 ;
      RECT 6.100000 2.435000 6.380000 2.860000 ;
      RECT 6.100000 3.000000 6.380000 3.420000 ;
      RECT 6.100000 3.560000 6.380000 3.980000 ;
      RECT 6.100000 4.870000 6.380000 5.290000 ;
      RECT 6.100000 5.430000 6.380000 5.850000 ;
      RECT 6.100000 5.990000 6.380000 6.415000 ;
      RECT 6.100000 6.695000 6.380000 7.120000 ;
      RECT 6.100000 7.260000 6.380000 7.680000 ;
      RECT 6.100000 7.820000 6.380000 8.240000 ;
      RECT 6.105000 0.000000 6.375000 0.470000 ;
      RECT 6.105000 4.120000 6.375000 4.730000 ;
      RECT 6.105000 8.380000 6.375000 8.850000 ;
      RECT 6.515000 0.000000 8.430000 0.330000 ;
      RECT 6.515000 4.260000 8.430000 4.590000 ;
      RECT 6.515000 8.520000 8.430000 8.850000 ;
      RECT 6.520000 0.750000 8.430000 0.890000 ;
      RECT 6.520000 1.310000 8.430000 1.450000 ;
      RECT 6.520000 1.870000 8.430000 2.010000 ;
      RECT 6.520000 2.580000 8.430000 2.720000 ;
      RECT 6.520000 3.140000 8.430000 3.280000 ;
      RECT 6.520000 3.700000 8.430000 3.840000 ;
      RECT 6.520000 5.010000 8.430000 5.150000 ;
      RECT 6.520000 5.570000 8.430000 5.710000 ;
      RECT 6.520000 6.130000 8.430000 6.270000 ;
      RECT 6.520000 6.840000 8.430000 6.980000 ;
      RECT 6.520000 7.400000 8.430000 7.540000 ;
      RECT 6.520000 7.960000 8.430000 8.100000 ;
      RECT 8.100000 0.330000 8.430000 0.750000 ;
      RECT 8.100000 0.890000 8.430000 1.310000 ;
      RECT 8.100000 1.450000 8.430000 1.870000 ;
      RECT 8.100000 2.010000 8.430000 2.020000 ;
      RECT 8.100000 2.570000 8.430000 2.580000 ;
      RECT 8.100000 2.720000 8.430000 3.140000 ;
      RECT 8.100000 3.280000 8.430000 3.700000 ;
      RECT 8.100000 3.840000 8.430000 4.260000 ;
      RECT 8.100000 4.590000 8.430000 5.010000 ;
      RECT 8.100000 5.150000 8.430000 5.570000 ;
      RECT 8.100000 5.710000 8.430000 6.130000 ;
      RECT 8.100000 6.270000 8.430000 6.280000 ;
      RECT 8.100000 6.830000 8.430000 6.840000 ;
      RECT 8.100000 6.980000 8.430000 7.400000 ;
      RECT 8.100000 7.540000 8.430000 7.960000 ;
      RECT 8.100000 8.100000 8.430000 8.520000 ;
    LAYER met4 ;
      RECT 0.370000 0.370000 1.870000 1.870000 ;
      RECT 0.370000 2.720000 1.870000 4.220000 ;
      RECT 0.370000 4.630000 1.870000 6.130000 ;
      RECT 0.370000 6.980000 1.870000 8.480000 ;
      RECT 2.510000 0.370000 4.010000 1.870000 ;
      RECT 2.510000 2.720000 4.010000 4.220000 ;
      RECT 2.510000 4.630000 4.010000 6.130000 ;
      RECT 2.510000 6.980000 4.010000 8.480000 ;
      RECT 4.420000 0.370000 5.920000 1.870000 ;
      RECT 4.420000 2.720000 5.920000 4.220000 ;
      RECT 4.420000 4.630000 5.920000 6.130000 ;
      RECT 4.420000 6.980000 5.920000 8.480000 ;
      RECT 6.560000 0.370000 8.060000 1.870000 ;
      RECT 6.560000 2.720000 8.060000 4.220000 ;
      RECT 6.560000 4.630000 8.060000 6.130000 ;
      RECT 6.560000 6.980000 8.060000 8.480000 ;
    LAYER pwell ;
      RECT 2.335000 1.750000 2.455000 2.005000 ;
      RECT 2.335000 6.010000 2.455000 6.265000 ;
      RECT 6.385000 1.750000 6.505000 2.005000 ;
      RECT 6.385000 6.010000 6.505000 6.265000 ;
    LAYER via ;
      RECT 0.035000 0.380000 0.295000 0.640000 ;
      RECT 0.035000 0.700000 0.295000 0.960000 ;
      RECT 0.035000 1.020000 0.295000 1.280000 ;
      RECT 0.035000 1.340000 0.295000 1.600000 ;
      RECT 0.035000 1.660000 0.295000 1.920000 ;
      RECT 0.035000 2.670000 0.295000 2.930000 ;
      RECT 0.035000 2.990000 0.295000 3.250000 ;
      RECT 0.035000 3.310000 0.295000 3.570000 ;
      RECT 0.035000 3.630000 0.295000 3.890000 ;
      RECT 0.035000 3.950000 0.295000 4.210000 ;
      RECT 0.035000 4.640000 0.295000 4.900000 ;
      RECT 0.035000 4.960000 0.295000 5.220000 ;
      RECT 0.035000 5.280000 0.295000 5.540000 ;
      RECT 0.035000 5.600000 0.295000 5.860000 ;
      RECT 0.035000 5.920000 0.295000 6.180000 ;
      RECT 0.035000 6.930000 0.295000 7.190000 ;
      RECT 0.035000 7.250000 0.295000 7.510000 ;
      RECT 0.035000 7.570000 0.295000 7.830000 ;
      RECT 0.035000 7.890000 0.295000 8.150000 ;
      RECT 0.035000 8.210000 0.295000 8.470000 ;
      RECT 0.260000 0.035000 0.520000 0.295000 ;
      RECT 0.260000 4.295000 0.520000 4.555000 ;
      RECT 0.260000 8.555000 0.520000 8.815000 ;
      RECT 0.580000 0.035000 0.840000 0.295000 ;
      RECT 0.580000 4.295000 0.840000 4.555000 ;
      RECT 0.580000 8.555000 0.840000 8.815000 ;
      RECT 0.595000 2.165000 0.855000 2.425000 ;
      RECT 0.595000 6.425000 0.855000 6.685000 ;
      RECT 0.900000 0.035000 1.160000 0.295000 ;
      RECT 0.900000 4.295000 1.160000 4.555000 ;
      RECT 0.900000 8.555000 1.160000 8.815000 ;
      RECT 0.915000 2.165000 1.175000 2.425000 ;
      RECT 0.915000 6.425000 1.175000 6.685000 ;
      RECT 1.220000 0.035000 1.480000 0.295000 ;
      RECT 1.220000 4.295000 1.480000 4.555000 ;
      RECT 1.220000 8.555000 1.480000 8.815000 ;
      RECT 1.235000 2.165000 1.495000 2.425000 ;
      RECT 1.235000 6.425000 1.495000 6.685000 ;
      RECT 1.540000 0.035000 1.800000 0.295000 ;
      RECT 1.540000 4.295000 1.800000 4.555000 ;
      RECT 1.540000 8.555000 1.800000 8.815000 ;
      RECT 1.555000 2.165000 1.815000 2.425000 ;
      RECT 1.555000 6.425000 1.815000 6.685000 ;
      RECT 2.060000 0.500000 2.320000 0.760000 ;
      RECT 2.060000 0.820000 2.320000 1.080000 ;
      RECT 2.060000 1.140000 2.320000 1.400000 ;
      RECT 2.060000 1.460000 2.320000 1.720000 ;
      RECT 2.060000 1.780000 2.320000 2.040000 ;
      RECT 2.060000 2.550000 2.320000 2.810000 ;
      RECT 2.060000 2.870000 2.320000 3.130000 ;
      RECT 2.060000 3.190000 2.320000 3.450000 ;
      RECT 2.060000 3.510000 2.320000 3.770000 ;
      RECT 2.060000 3.830000 2.320000 4.090000 ;
      RECT 2.060000 4.760000 2.320000 5.020000 ;
      RECT 2.060000 5.080000 2.320000 5.340000 ;
      RECT 2.060000 5.400000 2.320000 5.660000 ;
      RECT 2.060000 5.720000 2.320000 5.980000 ;
      RECT 2.060000 6.040000 2.320000 6.300000 ;
      RECT 2.060000 6.810000 2.320000 7.070000 ;
      RECT 2.060000 7.130000 2.320000 7.390000 ;
      RECT 2.060000 7.450000 2.320000 7.710000 ;
      RECT 2.060000 7.770000 2.320000 8.030000 ;
      RECT 2.060000 8.090000 2.320000 8.350000 ;
      RECT 2.565000 2.165000 2.825000 2.425000 ;
      RECT 2.565000 6.425000 2.825000 6.685000 ;
      RECT 2.580000 0.035000 2.840000 0.295000 ;
      RECT 2.580000 4.295000 2.840000 4.555000 ;
      RECT 2.580000 8.555000 2.840000 8.815000 ;
      RECT 2.885000 2.165000 3.145000 2.425000 ;
      RECT 2.885000 6.425000 3.145000 6.685000 ;
      RECT 2.900000 0.035000 3.160000 0.295000 ;
      RECT 2.900000 4.295000 3.160000 4.555000 ;
      RECT 2.900000 8.555000 3.160000 8.815000 ;
      RECT 3.205000 2.165000 3.465000 2.425000 ;
      RECT 3.205000 6.425000 3.465000 6.685000 ;
      RECT 3.220000 0.035000 3.480000 0.295000 ;
      RECT 3.220000 4.295000 3.480000 4.555000 ;
      RECT 3.220000 8.555000 3.480000 8.815000 ;
      RECT 3.525000 2.165000 3.785000 2.425000 ;
      RECT 3.525000 6.425000 3.785000 6.685000 ;
      RECT 3.540000 0.035000 3.800000 0.295000 ;
      RECT 3.540000 4.295000 3.800000 4.555000 ;
      RECT 3.540000 8.555000 3.800000 8.815000 ;
      RECT 3.860000 0.035000 4.120000 0.295000 ;
      RECT 3.860000 4.295000 4.120000 4.555000 ;
      RECT 3.860000 8.555000 4.120000 8.815000 ;
      RECT 4.085000 0.380000 4.345000 0.640000 ;
      RECT 4.085000 0.700000 4.345000 0.960000 ;
      RECT 4.085000 1.020000 4.345000 1.280000 ;
      RECT 4.085000 1.340000 4.345000 1.600000 ;
      RECT 4.085000 1.660000 4.345000 1.920000 ;
      RECT 4.085000 2.670000 4.345000 2.930000 ;
      RECT 4.085000 2.990000 4.345000 3.250000 ;
      RECT 4.085000 3.310000 4.345000 3.570000 ;
      RECT 4.085000 3.630000 4.345000 3.890000 ;
      RECT 4.085000 3.950000 4.345000 4.210000 ;
      RECT 4.085000 4.640000 4.345000 4.900000 ;
      RECT 4.085000 4.960000 4.345000 5.220000 ;
      RECT 4.085000 5.280000 4.345000 5.540000 ;
      RECT 4.085000 5.600000 4.345000 5.860000 ;
      RECT 4.085000 5.920000 4.345000 6.180000 ;
      RECT 4.085000 6.930000 4.345000 7.190000 ;
      RECT 4.085000 7.250000 4.345000 7.510000 ;
      RECT 4.085000 7.570000 4.345000 7.830000 ;
      RECT 4.085000 7.890000 4.345000 8.150000 ;
      RECT 4.085000 8.210000 4.345000 8.470000 ;
      RECT 4.310000 0.035000 4.570000 0.295000 ;
      RECT 4.310000 4.295000 4.570000 4.555000 ;
      RECT 4.310000 8.555000 4.570000 8.815000 ;
      RECT 4.630000 0.035000 4.890000 0.295000 ;
      RECT 4.630000 4.295000 4.890000 4.555000 ;
      RECT 4.630000 8.555000 4.890000 8.815000 ;
      RECT 4.645000 2.165000 4.905000 2.425000 ;
      RECT 4.645000 6.425000 4.905000 6.685000 ;
      RECT 4.950000 0.035000 5.210000 0.295000 ;
      RECT 4.950000 4.295000 5.210000 4.555000 ;
      RECT 4.950000 8.555000 5.210000 8.815000 ;
      RECT 4.965000 2.165000 5.225000 2.425000 ;
      RECT 4.965000 6.425000 5.225000 6.685000 ;
      RECT 5.270000 0.035000 5.530000 0.295000 ;
      RECT 5.270000 4.295000 5.530000 4.555000 ;
      RECT 5.270000 8.555000 5.530000 8.815000 ;
      RECT 5.285000 2.165000 5.545000 2.425000 ;
      RECT 5.285000 6.425000 5.545000 6.685000 ;
      RECT 5.590000 0.035000 5.850000 0.295000 ;
      RECT 5.590000 4.295000 5.850000 4.555000 ;
      RECT 5.590000 8.555000 5.850000 8.815000 ;
      RECT 5.605000 2.165000 5.865000 2.425000 ;
      RECT 5.605000 6.425000 5.865000 6.685000 ;
      RECT 6.110000 0.500000 6.370000 0.760000 ;
      RECT 6.110000 0.820000 6.370000 1.080000 ;
      RECT 6.110000 1.140000 6.370000 1.400000 ;
      RECT 6.110000 1.460000 6.370000 1.720000 ;
      RECT 6.110000 1.780000 6.370000 2.040000 ;
      RECT 6.110000 2.550000 6.370000 2.810000 ;
      RECT 6.110000 2.870000 6.370000 3.130000 ;
      RECT 6.110000 3.190000 6.370000 3.450000 ;
      RECT 6.110000 3.510000 6.370000 3.770000 ;
      RECT 6.110000 3.830000 6.370000 4.090000 ;
      RECT 6.110000 4.760000 6.370000 5.020000 ;
      RECT 6.110000 5.080000 6.370000 5.340000 ;
      RECT 6.110000 5.400000 6.370000 5.660000 ;
      RECT 6.110000 5.720000 6.370000 5.980000 ;
      RECT 6.110000 6.040000 6.370000 6.300000 ;
      RECT 6.110000 6.810000 6.370000 7.070000 ;
      RECT 6.110000 7.130000 6.370000 7.390000 ;
      RECT 6.110000 7.450000 6.370000 7.710000 ;
      RECT 6.110000 7.770000 6.370000 8.030000 ;
      RECT 6.110000 8.090000 6.370000 8.350000 ;
      RECT 6.615000 2.165000 6.875000 2.425000 ;
      RECT 6.615000 6.425000 6.875000 6.685000 ;
      RECT 6.630000 0.035000 6.890000 0.295000 ;
      RECT 6.630000 4.295000 6.890000 4.555000 ;
      RECT 6.630000 8.555000 6.890000 8.815000 ;
      RECT 6.935000 2.165000 7.195000 2.425000 ;
      RECT 6.935000 6.425000 7.195000 6.685000 ;
      RECT 6.950000 0.035000 7.210000 0.295000 ;
      RECT 6.950000 4.295000 7.210000 4.555000 ;
      RECT 6.950000 8.555000 7.210000 8.815000 ;
      RECT 7.255000 2.165000 7.515000 2.425000 ;
      RECT 7.255000 6.425000 7.515000 6.685000 ;
      RECT 7.270000 0.035000 7.530000 0.295000 ;
      RECT 7.270000 4.295000 7.530000 4.555000 ;
      RECT 7.270000 8.555000 7.530000 8.815000 ;
      RECT 7.575000 2.165000 7.835000 2.425000 ;
      RECT 7.575000 6.425000 7.835000 6.685000 ;
      RECT 7.590000 0.035000 7.850000 0.295000 ;
      RECT 7.590000 4.295000 7.850000 4.555000 ;
      RECT 7.590000 8.555000 7.850000 8.815000 ;
      RECT 7.910000 0.035000 8.170000 0.295000 ;
      RECT 7.910000 4.295000 8.170000 4.555000 ;
      RECT 7.910000 8.555000 8.170000 8.815000 ;
      RECT 8.135000 0.380000 8.395000 0.640000 ;
      RECT 8.135000 0.700000 8.395000 0.960000 ;
      RECT 8.135000 1.020000 8.395000 1.280000 ;
      RECT 8.135000 1.340000 8.395000 1.600000 ;
      RECT 8.135000 1.660000 8.395000 1.920000 ;
      RECT 8.135000 2.670000 8.395000 2.930000 ;
      RECT 8.135000 2.990000 8.395000 3.250000 ;
      RECT 8.135000 3.310000 8.395000 3.570000 ;
      RECT 8.135000 3.630000 8.395000 3.890000 ;
      RECT 8.135000 3.950000 8.395000 4.210000 ;
      RECT 8.135000 4.640000 8.395000 4.900000 ;
      RECT 8.135000 4.960000 8.395000 5.220000 ;
      RECT 8.135000 5.280000 8.395000 5.540000 ;
      RECT 8.135000 5.600000 8.395000 5.860000 ;
      RECT 8.135000 5.920000 8.395000 6.180000 ;
      RECT 8.135000 6.930000 8.395000 7.190000 ;
      RECT 8.135000 7.250000 8.395000 7.510000 ;
      RECT 8.135000 7.570000 8.395000 7.830000 ;
      RECT 8.135000 7.890000 8.395000 8.150000 ;
      RECT 8.135000 8.210000 8.395000 8.470000 ;
    LAYER via2 ;
      RECT 0.025000 0.495000 0.305000 0.775000 ;
      RECT 0.025000 0.895000 0.305000 1.175000 ;
      RECT 0.025000 1.295000 0.305000 1.575000 ;
      RECT 0.025000 1.695000 0.305000 1.975000 ;
      RECT 0.025000 2.615000 0.305000 2.895000 ;
      RECT 0.025000 3.015000 0.305000 3.295000 ;
      RECT 0.025000 3.415000 0.305000 3.695000 ;
      RECT 0.025000 3.815000 0.305000 4.095000 ;
      RECT 0.025000 4.755000 0.305000 5.035000 ;
      RECT 0.025000 5.155000 0.305000 5.435000 ;
      RECT 0.025000 5.555000 0.305000 5.835000 ;
      RECT 0.025000 5.955000 0.305000 6.235000 ;
      RECT 0.025000 6.875000 0.305000 7.155000 ;
      RECT 0.025000 7.275000 0.305000 7.555000 ;
      RECT 0.025000 7.675000 0.305000 7.955000 ;
      RECT 0.025000 8.075000 0.305000 8.355000 ;
      RECT 0.390000 0.025000 0.670000 0.305000 ;
      RECT 0.390000 4.285000 0.670000 4.565000 ;
      RECT 0.390000 8.545000 0.670000 8.825000 ;
      RECT 0.790000 0.025000 1.070000 0.305000 ;
      RECT 0.790000 4.285000 1.070000 4.565000 ;
      RECT 0.790000 8.545000 1.070000 8.825000 ;
      RECT 0.850000 2.155000 1.130000 2.435000 ;
      RECT 0.850000 6.415000 1.130000 6.695000 ;
      RECT 1.190000 0.025000 1.470000 0.305000 ;
      RECT 1.190000 4.285000 1.470000 4.565000 ;
      RECT 1.190000 8.545000 1.470000 8.825000 ;
      RECT 1.250000 2.155000 1.530000 2.435000 ;
      RECT 1.250000 6.415000 1.530000 6.695000 ;
      RECT 1.590000 0.025000 1.870000 0.305000 ;
      RECT 1.590000 4.285000 1.870000 4.565000 ;
      RECT 1.590000 8.545000 1.870000 8.825000 ;
      RECT 1.650000 2.155000 1.930000 2.435000 ;
      RECT 1.650000 6.415000 1.930000 6.695000 ;
      RECT 2.050000 0.955000 2.330000 1.235000 ;
      RECT 2.050000 1.355000 2.330000 1.635000 ;
      RECT 2.050000 1.755000 2.330000 2.035000 ;
      RECT 2.050000 2.155000 2.330000 2.435000 ;
      RECT 2.050000 2.555000 2.330000 2.835000 ;
      RECT 2.050000 2.955000 2.330000 3.235000 ;
      RECT 2.050000 3.355000 2.330000 3.635000 ;
      RECT 2.050000 5.215000 2.330000 5.495000 ;
      RECT 2.050000 5.615000 2.330000 5.895000 ;
      RECT 2.050000 6.015000 2.330000 6.295000 ;
      RECT 2.050000 6.415000 2.330000 6.695000 ;
      RECT 2.050000 6.815000 2.330000 7.095000 ;
      RECT 2.050000 7.215000 2.330000 7.495000 ;
      RECT 2.050000 7.615000 2.330000 7.895000 ;
      RECT 2.450000 2.155000 2.730000 2.435000 ;
      RECT 2.450000 6.415000 2.730000 6.695000 ;
      RECT 2.510000 0.025000 2.790000 0.305000 ;
      RECT 2.510000 4.285000 2.790000 4.565000 ;
      RECT 2.510000 8.545000 2.790000 8.825000 ;
      RECT 2.850000 2.155000 3.130000 2.435000 ;
      RECT 2.850000 6.415000 3.130000 6.695000 ;
      RECT 2.910000 0.025000 3.190000 0.305000 ;
      RECT 2.910000 4.285000 3.190000 4.565000 ;
      RECT 2.910000 8.545000 3.190000 8.825000 ;
      RECT 3.250000 2.155000 3.530000 2.435000 ;
      RECT 3.250000 6.415000 3.530000 6.695000 ;
      RECT 3.310000 0.025000 3.590000 0.305000 ;
      RECT 3.310000 4.285000 3.590000 4.565000 ;
      RECT 3.310000 8.545000 3.590000 8.825000 ;
      RECT 3.710000 0.025000 3.990000 0.305000 ;
      RECT 3.710000 4.285000 3.990000 4.565000 ;
      RECT 3.710000 8.545000 3.990000 8.825000 ;
      RECT 4.075000 0.495000 4.355000 0.775000 ;
      RECT 4.075000 0.895000 4.355000 1.175000 ;
      RECT 4.075000 1.295000 4.355000 1.575000 ;
      RECT 4.075000 1.695000 4.355000 1.975000 ;
      RECT 4.075000 2.615000 4.355000 2.895000 ;
      RECT 4.075000 3.015000 4.355000 3.295000 ;
      RECT 4.075000 3.415000 4.355000 3.695000 ;
      RECT 4.075000 3.815000 4.355000 4.095000 ;
      RECT 4.075000 4.755000 4.355000 5.035000 ;
      RECT 4.075000 5.155000 4.355000 5.435000 ;
      RECT 4.075000 5.555000 4.355000 5.835000 ;
      RECT 4.075000 5.955000 4.355000 6.235000 ;
      RECT 4.075000 6.875000 4.355000 7.155000 ;
      RECT 4.075000 7.275000 4.355000 7.555000 ;
      RECT 4.075000 7.675000 4.355000 7.955000 ;
      RECT 4.075000 8.075000 4.355000 8.355000 ;
      RECT 4.440000 0.025000 4.720000 0.305000 ;
      RECT 4.440000 4.285000 4.720000 4.565000 ;
      RECT 4.440000 8.545000 4.720000 8.825000 ;
      RECT 4.840000 0.025000 5.120000 0.305000 ;
      RECT 4.840000 4.285000 5.120000 4.565000 ;
      RECT 4.840000 8.545000 5.120000 8.825000 ;
      RECT 4.900000 2.155000 5.180000 2.435000 ;
      RECT 4.900000 6.415000 5.180000 6.695000 ;
      RECT 5.240000 0.025000 5.520000 0.305000 ;
      RECT 5.240000 4.285000 5.520000 4.565000 ;
      RECT 5.240000 8.545000 5.520000 8.825000 ;
      RECT 5.300000 2.155000 5.580000 2.435000 ;
      RECT 5.300000 6.415000 5.580000 6.695000 ;
      RECT 5.640000 0.025000 5.920000 0.305000 ;
      RECT 5.640000 4.285000 5.920000 4.565000 ;
      RECT 5.640000 8.545000 5.920000 8.825000 ;
      RECT 5.700000 2.155000 5.980000 2.435000 ;
      RECT 5.700000 6.415000 5.980000 6.695000 ;
      RECT 6.100000 0.955000 6.380000 1.235000 ;
      RECT 6.100000 1.355000 6.380000 1.635000 ;
      RECT 6.100000 1.755000 6.380000 2.035000 ;
      RECT 6.100000 2.155000 6.380000 2.435000 ;
      RECT 6.100000 2.555000 6.380000 2.835000 ;
      RECT 6.100000 2.955000 6.380000 3.235000 ;
      RECT 6.100000 3.355000 6.380000 3.635000 ;
      RECT 6.100000 5.215000 6.380000 5.495000 ;
      RECT 6.100000 5.615000 6.380000 5.895000 ;
      RECT 6.100000 6.015000 6.380000 6.295000 ;
      RECT 6.100000 6.415000 6.380000 6.695000 ;
      RECT 6.100000 6.815000 6.380000 7.095000 ;
      RECT 6.100000 7.215000 6.380000 7.495000 ;
      RECT 6.100000 7.615000 6.380000 7.895000 ;
      RECT 6.500000 2.155000 6.780000 2.435000 ;
      RECT 6.500000 6.415000 6.780000 6.695000 ;
      RECT 6.560000 0.025000 6.840000 0.305000 ;
      RECT 6.560000 4.285000 6.840000 4.565000 ;
      RECT 6.560000 8.545000 6.840000 8.825000 ;
      RECT 6.900000 2.155000 7.180000 2.435000 ;
      RECT 6.900000 6.415000 7.180000 6.695000 ;
      RECT 6.960000 0.025000 7.240000 0.305000 ;
      RECT 6.960000 4.285000 7.240000 4.565000 ;
      RECT 6.960000 8.545000 7.240000 8.825000 ;
      RECT 7.300000 2.155000 7.580000 2.435000 ;
      RECT 7.300000 6.415000 7.580000 6.695000 ;
      RECT 7.360000 0.025000 7.640000 0.305000 ;
      RECT 7.360000 4.285000 7.640000 4.565000 ;
      RECT 7.360000 8.545000 7.640000 8.825000 ;
      RECT 7.760000 0.025000 8.040000 0.305000 ;
      RECT 7.760000 4.285000 8.040000 4.565000 ;
      RECT 7.760000 8.545000 8.040000 8.825000 ;
      RECT 8.125000 0.495000 8.405000 0.775000 ;
      RECT 8.125000 0.895000 8.405000 1.175000 ;
      RECT 8.125000 1.295000 8.405000 1.575000 ;
      RECT 8.125000 1.695000 8.405000 1.975000 ;
      RECT 8.125000 2.615000 8.405000 2.895000 ;
      RECT 8.125000 3.015000 8.405000 3.295000 ;
      RECT 8.125000 3.415000 8.405000 3.695000 ;
      RECT 8.125000 3.815000 8.405000 4.095000 ;
      RECT 8.125000 4.755000 8.405000 5.035000 ;
      RECT 8.125000 5.155000 8.405000 5.435000 ;
      RECT 8.125000 5.555000 8.405000 5.835000 ;
      RECT 8.125000 5.955000 8.405000 6.235000 ;
      RECT 8.125000 6.875000 8.405000 7.155000 ;
      RECT 8.125000 7.275000 8.405000 7.555000 ;
      RECT 8.125000 7.675000 8.405000 7.955000 ;
      RECT 8.125000 8.075000 8.405000 8.355000 ;
  END
END sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4_top
END LIBRARY
