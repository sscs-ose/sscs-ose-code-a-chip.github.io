# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15 ;
  ORIGIN  0.000000 -0.020000 ;
  SIZE  4.420000 BY  6.160000 ;
  PIN DRAIN
    ANTENNADIFFAREA  6.262000 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1.980000 4.420000 4.220000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.030000 ;
    PORT
      LAYER met1 ;
        RECT 0.910000 0.040000 3.720000 0.330000 ;
        RECT 0.910000 5.870000 3.720000 6.160000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  6.034750 ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.560000 4.420000 1.840000 ;
        RECT 0.000000 4.360000 4.420000 5.645000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  1.464500 ;
    PORT
      LAYER met1 ;
        RECT 0.130000 0.615000 0.420000 5.585000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.190000 0.675000 0.360000 5.525000 ;
      RECT 0.745000 0.555000 0.915000 5.645000 ;
      RECT 0.970000 0.100000 3.680000 0.270000 ;
      RECT 0.970000 5.930000 3.680000 6.100000 ;
      RECT 1.165000 0.555000 1.695000 5.645000 ;
      RECT 1.935000 0.555000 2.465000 5.645000 ;
      RECT 2.705000 0.555000 3.235000 5.645000 ;
      RECT 3.485000 0.555000 3.655000 5.645000 ;
      RECT 4.055000 0.675000 4.225000 5.525000 ;
    LAYER mcon ;
      RECT 0.190000 1.035000 0.360000 1.205000 ;
      RECT 0.190000 1.395000 0.360000 1.565000 ;
      RECT 0.190000 1.755000 0.360000 1.925000 ;
      RECT 0.190000 2.115000 0.360000 2.285000 ;
      RECT 0.190000 2.475000 0.360000 2.645000 ;
      RECT 0.190000 2.835000 0.360000 3.005000 ;
      RECT 0.190000 3.195000 0.360000 3.365000 ;
      RECT 0.190000 3.555000 0.360000 3.725000 ;
      RECT 0.190000 3.915000 0.360000 4.085000 ;
      RECT 0.190000 4.275000 0.360000 4.445000 ;
      RECT 0.190000 4.635000 0.360000 4.805000 ;
      RECT 0.190000 4.995000 0.360000 5.165000 ;
      RECT 0.190000 5.355000 0.360000 5.525000 ;
      RECT 0.745000 0.675000 0.915000 0.845000 ;
      RECT 0.745000 1.035000 0.915000 1.205000 ;
      RECT 0.745000 1.395000 0.915000 1.565000 ;
      RECT 0.745000 1.755000 0.915000 1.925000 ;
      RECT 0.745000 2.115000 0.915000 2.285000 ;
      RECT 0.745000 2.475000 0.915000 2.645000 ;
      RECT 0.745000 2.835000 0.915000 3.005000 ;
      RECT 0.745000 3.195000 0.915000 3.365000 ;
      RECT 0.745000 3.555000 0.915000 3.725000 ;
      RECT 0.745000 3.915000 0.915000 4.085000 ;
      RECT 0.745000 4.275000 0.915000 4.445000 ;
      RECT 0.745000 4.635000 0.915000 4.805000 ;
      RECT 0.745000 4.995000 0.915000 5.165000 ;
      RECT 0.745000 5.355000 0.915000 5.525000 ;
      RECT 0.970000 0.100000 1.140000 0.270000 ;
      RECT 0.970000 5.930000 1.140000 6.100000 ;
      RECT 1.165000 0.675000 1.695000 5.525000 ;
      RECT 1.330000 0.100000 1.500000 0.270000 ;
      RECT 1.330000 5.930000 1.500000 6.100000 ;
      RECT 1.690000 0.100000 1.860000 0.270000 ;
      RECT 1.690000 5.930000 1.860000 6.100000 ;
      RECT 1.935000 0.675000 2.465000 5.525000 ;
      RECT 2.050000 0.100000 2.220000 0.270000 ;
      RECT 2.050000 5.930000 2.220000 6.100000 ;
      RECT 2.410000 0.100000 2.580000 0.270000 ;
      RECT 2.410000 5.930000 2.580000 6.100000 ;
      RECT 2.705000 0.675000 3.235000 5.525000 ;
      RECT 2.770000 0.100000 2.940000 0.270000 ;
      RECT 2.770000 5.930000 2.940000 6.100000 ;
      RECT 3.130000 0.100000 3.300000 0.270000 ;
      RECT 3.130000 5.930000 3.300000 6.100000 ;
      RECT 3.485000 0.675000 3.655000 0.845000 ;
      RECT 3.485000 1.035000 3.655000 1.205000 ;
      RECT 3.485000 1.395000 3.655000 1.565000 ;
      RECT 3.485000 1.755000 3.655000 1.925000 ;
      RECT 3.485000 2.115000 3.655000 2.285000 ;
      RECT 3.485000 2.475000 3.655000 2.645000 ;
      RECT 3.485000 2.835000 3.655000 3.005000 ;
      RECT 3.485000 3.195000 3.655000 3.365000 ;
      RECT 3.485000 3.555000 3.655000 3.725000 ;
      RECT 3.485000 3.915000 3.655000 4.085000 ;
      RECT 3.485000 4.275000 3.655000 4.445000 ;
      RECT 3.485000 4.635000 3.655000 4.805000 ;
      RECT 3.485000 4.995000 3.655000 5.165000 ;
      RECT 3.485000 5.355000 3.655000 5.525000 ;
      RECT 3.490000 0.100000 3.660000 0.270000 ;
      RECT 3.490000 5.930000 3.660000 6.100000 ;
      RECT 4.055000 1.035000 4.225000 1.205000 ;
      RECT 4.055000 1.395000 4.225000 1.565000 ;
      RECT 4.055000 1.755000 4.225000 1.925000 ;
      RECT 4.055000 2.115000 4.225000 2.285000 ;
      RECT 4.055000 2.475000 4.225000 2.645000 ;
      RECT 4.055000 2.835000 4.225000 3.005000 ;
      RECT 4.055000 3.195000 4.225000 3.365000 ;
      RECT 4.055000 3.555000 4.225000 3.725000 ;
      RECT 4.055000 3.915000 4.225000 4.085000 ;
      RECT 4.055000 4.275000 4.225000 4.445000 ;
      RECT 4.055000 4.635000 4.225000 4.805000 ;
      RECT 4.055000 4.995000 4.225000 5.165000 ;
      RECT 4.055000 5.355000 4.225000 5.525000 ;
    LAYER met1 ;
      RECT 0.700000 0.560000 0.960000 0.615000 ;
      RECT 0.700000 0.615000 0.975000 5.585000 ;
      RECT 0.700000 5.585000 0.960000 5.640000 ;
      RECT 1.115000 0.615000 1.745000 5.585000 ;
      RECT 1.885000 0.615000 2.515000 5.585000 ;
      RECT 1.910000 0.560000 2.490000 0.615000 ;
      RECT 1.910000 5.585000 2.490000 5.645000 ;
      RECT 2.655000 0.615000 3.285000 5.585000 ;
      RECT 3.425000 0.615000 3.715000 5.585000 ;
      RECT 3.440000 0.560000 3.700000 0.615000 ;
      RECT 3.440000 5.585000 3.700000 5.645000 ;
      RECT 3.995000 0.615000 4.285000 5.585000 ;
    LAYER via ;
      RECT 0.700000 0.590000 0.960000 0.850000 ;
      RECT 0.700000 0.910000 0.960000 1.170000 ;
      RECT 0.700000 1.230000 0.960000 1.490000 ;
      RECT 0.700000 1.550000 0.960000 1.810000 ;
      RECT 0.700000 4.390000 0.960000 4.650000 ;
      RECT 0.700000 4.710000 0.960000 4.970000 ;
      RECT 0.700000 5.030000 0.960000 5.290000 ;
      RECT 0.700000 5.350000 0.960000 5.610000 ;
      RECT 1.140000 2.010000 1.720000 4.190000 ;
      RECT 1.910000 0.590000 2.490000 1.810000 ;
      RECT 1.910000 4.395000 2.490000 5.615000 ;
      RECT 2.680000 2.010000 3.260000 4.190000 ;
      RECT 3.440000 0.590000 3.700000 0.850000 ;
      RECT 3.440000 0.910000 3.700000 1.170000 ;
      RECT 3.440000 1.230000 3.700000 1.490000 ;
      RECT 3.440000 1.550000 3.700000 1.810000 ;
      RECT 3.440000 4.395000 3.700000 4.655000 ;
      RECT 3.440000 4.715000 3.700000 4.975000 ;
      RECT 3.440000 5.035000 3.700000 5.295000 ;
      RECT 3.440000 5.355000 3.700000 5.615000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15
END LIBRARY
