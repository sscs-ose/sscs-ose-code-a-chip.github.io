* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 05
.param
+ sky130_fd_pr__nfet_g5v0d16v0__toxe_mult = 0.94
+ sky130_fd_pr__nfet_g5v0d16v0__toxp_mult = 1.0
+ sky130_fd_pr__nfet_g5v0d16v0__overlap_mult = 0.10246
+ sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult = 8.1753e-1
+ sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult = 7.7786e-1
+ sky130_fd_pr__nfet_g5v0d16v0__rdiff_mult = 6.4330e-1
+ sky130_fd_pr__nfet_g5v0d16v0__lint_diff = 1.7325e-8
+ sky130_fd_pr__nfet_g5v0d16v0__dlc_diff = 1.7325e-8
+ sky130_fd_pr__nfet_g5v0d16v0__wint_diff = -3.2175e-8
+ sky130_fd_pr__nfet_g5v0d16v0__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 000, W = 20.0, L = 0.7
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_0 = -1.3425e-1
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_0 = 2.2191e-2
+ sky130_fd_pr__nfet_g5v0d16v0__k2_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ua_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ub_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_0 = -0.2485
+ sky130_fd_pr__nfet_g5v0d16v0__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ute_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_0 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__keta_diff_0 = 0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 001, W = 5.0, L = 0.7
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_1 = -0.14054
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_1 = 0.015572
+ sky130_fd_pr__nfet_g5v0d16v0__k2_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ua_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ub_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__a0_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ags_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_1 = -0.2485
+ sky130_fd_pr__nfet_g5v0d16v0__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ute_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_1 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__keta_diff_1 = 0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 002, W = 50.0, L = 0.7
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_2 = -0.13714
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_2 = 0.016601
+ sky130_fd_pr__nfet_g5v0d16v0__k2_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ua_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ub_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_2 = -0.2485
+ sky130_fd_pr__nfet_g5v0d16v0__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ute_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_2 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__keta_diff_2 = 0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 003, W = 20.0, L = 2.2
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_3 = -0.097324
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_3 = 0.004226
+ sky130_fd_pr__nfet_g5v0d16v0__k2_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ua_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ub_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_3 = 0.667
+ sky130_fd_pr__nfet_g5v0d16v0__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ute_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_3 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__keta_diff_3 = 0.0
*
* sky130_fd_pr__nfet_g5v0d16v0, Bin 004, W = 20.0, L = 2.2
* --------------------------------
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_4 = -0.090898
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_4 = 0.0020803
+ sky130_fd_pr__nfet_g5v0d16v0__k2_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ua_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ub_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_4 = 1.16
+ sky130_fd_pr__nfet_g5v0d16v0__voff_diff_4 = -0.1
+ sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__ute_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_4 = 0.0
+ sky130_fd_pr__nfet_g5v0d16v0__keta_diff_4 = 0.0
.include "sky130_fd_pr__nfet_g5v0d16v0__subcircuit.pm3.spice"
.include "sky130_fd_pr__nfet_g5v0d16v0.pm3.spice"
