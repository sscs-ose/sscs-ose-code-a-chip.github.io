** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/tb_cm_ota_working_v2_extracted.sch
**.subckt tb_cm_ota_working_v2_extracted
V1 avdd_1v8_ext GND 1.8
C1 out_ext GND 250f m=1
V3 inn_ext GND DC 1 AC 1
V4 inp_ext GND 1
X1 iref_ext out_ext inn_ext inp_ext GND avdd_1v8_ext cm_ota_extracted
I1 GND iref_ext 25.2u

V10 vdd GND 1.8
C10 out GND 250f m=1
V30 inn GND DC 1
V40 inp GND DC 1 AC 1
X10 vdd out inp inn itail GND cm_ota w1_2=5.88 w3_4=10.08 w5_6=19.32 w7_8=35.28 w9_10=11.76 beta=1 nf1_2=1 nf3_4=1 nf5_6=1 nf7_8=1 nf9_10=1
I30 GND itail 26.2u


.lib /opt/pdk/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.temp 27

.save all
.control
	ac dec 100 1 1e15
	
	plot vdb(out) vdb(out_ext)vs frequency
	plot (180*cph(out)/pi) (180*cph(out_ext)/pi)vs frequency
	
	let phase_vector = 180*cph(out)/pi
	let gain_vector = vdb(out)
	
	meas ac unity_gain_freq_val when vdb(out)=0
	meas ac unity_gain_freq_val_ext when vdb(out_ext)=0

	meas ac dc_gain_val find vdb(out) at=10Hz
	meas ac dc_gain_val_ext find vdb(out_ext) at=10Hz


	write tb_cm_ota_working_v2_extracted.raw
	// set hcopyscolor=1 //v1
	echo 'GBWP = ' gbw
	echo 'DC Gain = ' dc_gain
	echo 'pole1 freq = ' pole1_freq
	echo 'pole2 freq = ' pole2_freq
	echo '3dB BW = ' bandwidth
.endc

.subckt cm_ota vdd out inp inn itail vss  w1_2=1 w3_4=1 w5_6=1 w7_8=1 w9_10=1 beta=2 nf1_2=2 nf3_4=2 nf5_6=2 nf7_8=2 nf9_10=2
XM1 ds1_3 inn source source sky130_fd_pr__nfet_01v8 L=0.15 W=w1_2 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM3 ds1_3 ds1_3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=w3_4 nf=nf3_4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 ds2_4 inp source source sky130_fd_pr__nfet_01v8 L=0.15 W=w1_2 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM4 ds2_4 ds2_4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=w3_4 nf=nf3_4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM7 ds5_7 ds1_3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=w7_8 nf=nf7_8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 ds5_7 ds5_7 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=w5_6 nf=nf5_6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 out ds5_7 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=w5_6 nf=nf5_6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM8 out ds2_4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=w7_8 nf=nf7_8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 source itail vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=w9_10 nf=nf9_10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 itail itail vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=w9_10 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.subckt cm_ota_extracted ID VOUT VINN VINP VSS VDD
X0 m1_2236_5516# VINP m2_746_2735# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X1 m1_2236_5516# VINP m2_746_2735# VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X2 m2_746_2735# VINP m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X3 m2_746_2735# VINP m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X4 m1_2236_5516# VINP m2_746_2735# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X5 m1_2236_5516# VINP m2_746_2735# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X6 m2_746_2735# VINP m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X7 m2_746_2735# VINP m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X8 m1_2236_5516# VINN m2_2810_2735# VSS sky130_fd_pr__nfet_01v8 ad=9.31 pd=89.4 as=0.941 ps=8.96 w=0.84 l=0.15
X9 m1_2236_5516# VINN m2_2810_2735# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X10 m2_2810_2735# VINN m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X11 m2_2810_2735# VINN m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X12 m1_2236_5516# VINN m2_2810_2735# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X13 m1_2236_5516# VINN m2_2810_2735# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X14 m2_2810_2735# VINN m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X15 m2_2810_2735# VINN m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X16 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X17 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X18 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X19 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X20 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X21 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X22 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X23 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X24 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X25 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X26 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X27 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X28 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X29 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X30 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X31 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X32 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X33 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X34 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X35 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X36 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X37 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X38 m1_2236_5516# m1_828_5348# m1_828_5348# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X39 m1_828_5348# m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X40 VSS ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X41 ID ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X42 VSS ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X43 VSS ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X44 ID ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X45 VSS ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X46 ID ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X47 ID ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X48 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X49 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X50 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X51 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X52 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X53 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X54 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X55 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X56 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X57 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X58 m2_746_2735# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X59 VDD m2_746_2735# m2_746_2735# VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X60 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.41 pd=13.4 as=14.8 ps=143 w=0.84 l=0.15
X61 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X62 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X63 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X64 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X65 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X66 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X67 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X68 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X69 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X70 m2_2810_2735# m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X71 VDD m2_2810_2735# m2_2810_2735# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X72 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X73 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X74 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X75 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X76 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X77 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X78 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X79 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X80 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X81 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X82 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X83 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X84 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X85 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X86 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X87 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X88 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X89 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X90 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X91 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X92 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X93 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X94 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X95 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X96 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X97 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X98 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X99 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X100 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X101 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X102 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X103 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X104 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X105 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X106 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X107 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X108 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X109 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X110 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X111 VOUT m2_2810_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X112 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X113 VDD m2_2810_2735# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X114 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=4.94 ps=47 w=0.84 l=0.15
X115 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X116 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X117 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X118 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X119 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X120 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X121 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X122 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X123 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X124 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X125 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X126 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X127 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X128 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X129 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X130 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X131 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X132 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X133 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X134 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X135 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X136 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X137 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X138 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X139 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X140 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X141 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X142 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X143 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X144 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X145 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X146 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X147 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X148 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X149 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X150 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X151 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X152 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X153 m1_828_5348# m2_746_2735# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X154 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X155 VDD m2_746_2735# m1_828_5348# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X156 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X157 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X158 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X159 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X160 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X161 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X162 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X163 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X164 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X165 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X166 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X167 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X168 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X169 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X170 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X171 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X172 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X173 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X174 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X175 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X176 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X177 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X178 m1_2236_5516# m1_828_5348# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X179 VOUT m1_828_5348# m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X180 VSS ID m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X181 m1_2236_5516# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X182 VSS ID m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X183 VSS ID m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X184 m1_2236_5516# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X185 VSS ID m1_2236_5516# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X186 m1_2236_5516# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X187 m1_2236_5516# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
C0 m2_2810_2735# m1_828_5348# 0.0192f
C1 VDD m1_828_5348# 17.1f
C2 m1_2236_5516# VOUT 8.41f
C3 ID m1_828_5348# 0.00106f
C4 m2_746_2735# m1_2236_5516# 3.56f
C5 VDD VINP 0.0529f
C6 ID VINP 0.038f
C7 m2_2810_2735# VOUT 3.84f
C8 m1_2236_5516# VINN 0.377f
C9 VDD VOUT 17f
C10 ID VOUT 1.82e-19
C11 m2_746_2735# m2_2810_2735# 0.102f
C12 m2_746_2735# VDD 23.5f
C13 m2_746_2735# ID 0.116f
C14 VOUT m1_828_5348# 1.15f
C15 m2_2810_2735# m1_2236_5516# 3.1f
C16 VDD m1_2236_5516# 2.13f
C17 ID m1_2236_5516# 1.27f
C18 m2_746_2735# m1_828_5348# 3.78f
C19 m2_2810_2735# VINN 0.388f
C20 VDD VINN 0.0546f
C21 ID VINN 0.038f
C22 m2_746_2735# VINP 0.388f
C23 m1_2236_5516# m1_828_5348# 11.2f
C24 VINP m1_2236_5516# 0.377f
C25 VDD m2_2810_2735# 23.6f
C26 ID m2_2810_2735# 0.0149f
C27 VDD ID 0.137f
C28 m2_746_2735# VOUT 2.31e-19
C29 ID VSS 11.4f
C30 VOUT VSS 1.24f
C31 m1_828_5348# VSS 13.7f
C32 VDD VSS 57.6f
C33 m2_2810_2735# VSS 2.35f
C34 m2_746_2735# VSS 2.48f
C35 VINN VSS 2.15f
C36 m1_2236_5516# VSS 8.59f
C37 VINP VSS 2.17f


.ends
.GLOBAL GND
.end
