** sch_path: /home/GmTune/src/spice/GmCMFF.sch
**.subckt GmCMFF
V1 VDD GND VDD
V2 VSS GND 0
V3 VI VSS dc 0 ac 1 sin 0 vi fi
XM4 V11 V14 VDD VDD sky130_fd_pr__pfet_01v8 L=LMB W=WMB nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
E1 VIP net1 VI VSS 0.5
E2 VIN net1 VSS VI 0.5
XM5 net2 V14 VDD VDD sky130_fd_pr__pfet_01v8 L=LMB W=WMB nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 V14 V14 VDD VDD sky130_fd_pr__pfet_01v8 L=LMB W=WMB nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I1 V14 VSS I_B
VI1 V11 net3 0
.save i(vi1)
XM16 net3 VIP V12 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 V12 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=LM3 W=WM3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net4 VG V12 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V5 net1 VSS VCM
V6 VG GND VG
XM19 V15 net7 VDD VDD sky130_fd_pr__pfet_01v8 L=LM4 W=WM4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 net8 VG V12 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 net2 VIN net5 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 net5 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=LM3 W=WM3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 net7 VG net5 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 net6 VG net5 VSS sky130_fd_pr__nfet_01v8 L=LM1 W=WM1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net6 V13 VDD VDD sky130_fd_pr__pfet_01v8 L=LM4 W=WM4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VI3 V15 net4 0
.save i(vi3)
XM1 V13 V13 VDD VDD sky130_fd_pr__pfet_01v8 L=LM4 W=WM4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net7 net7 VDD VDD sky130_fd_pr__pfet_01v8 L=LM4 W=WM4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VI2 V13 net8 0
.save i(vi2)
R1 VDD VO1 2k m=1
I2 VDD net9 I_CM
VIO1 V15 net11 0
.save i(vio1)
R2 VDD VO2 2k m=1
VIO2 net6 net12 0
.save i(vio2)
XM3 net10 net9 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net9 net9 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 VO2 net9 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VI4 VO1 net10 0
.save i(vi4)
C1 net11 VO1 10u m=1
E3 VO VSS VO1 VO2 1
C2 VO2 net12 10u m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

.param VDD=1.8 VG=0.9 VCM=0.9 I_B=50u RLOAD=2k I_CM=250u vi=0.01 fi=10000 WMB=20u LMB=0.5u WM1=12u LM1=0.5u WM2=12u LM2=0.5u WM3=10u LM3=0.5u WM4=20u LM4=0.5u
.include /home/GmTune/src/spice/para.spice

.control
run
save all

op
print i(VI1) i(VI2) i(VI3) i(VI4) i(VIO1)
wrdata ckpts/IB.txt i(VI1)
wrdata ckpts/I1.txt i(VI2)
wrdata ckpts/I2.txt i(VI3)

ac dec 1000 1e6 1e9
let Gm = (i(VIO1) - i(VIO2)) / V(VI)
wrdata ckpts/Gm.txt Gm
wrdata ckpts/Gain.txt (Gm*2k)

noise V(VO) V3 dec 100 1e7 1e8
setplot noise1
wrdata ckpts/IRN.txt inoise_spectrum

*tran 10p 0.5u
*plot V(VO1) V(VO)
*plot i(VIO1)

*fourier 10000000 vo
*let idx = 2
*let sum_mag_square = 0
*while idx < 10
*   let mag = fourier11[1][idx]
*    let sum_mag_square = sum_mag_square + mag * mag
*    let idx = idx + 1
*end
*let root_sum_mag_square = sqrt(sum_mag_square)
*let thd = root_sum_mag_square / fourier11[1][1] * 100
*print thd
*wrdata ckpts/THD.txt thd

.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
