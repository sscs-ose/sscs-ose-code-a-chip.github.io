module approxMult_signed8x8 (A, B, OUT);
  input  [7:0] A;
  input  [7:0] B;
  output [15:0] OUT;
  wire n1, n10, n11, n12, n13, n14, n15, n2, n3, n4, n5, n6, n7, v0_0, v100_0, v101_0, v102_0, v103_0, v104_0, v105_0, v106_0, v107_0, v108_0, v109_0, v10_0, v110_0, v111_0, v112_0, v113_0, v114_0, v115_0, v116_0, v117_0, v118_0, v119_0, v11_0, v120_0, v121_0, v122_0, v123_0, v124_0, v125_0, v126_0, v127_0, v128_0, v129_0, v12_0, v130_0, v131_0, v132_0, v133_0, v134_0, v135_0, v136_0, v137_0, v138_0, v139_0, v13_0, v140_0, v141_0, v142_0, v143_0, v144_0, v145_0, v146_0, v147_0, v148_0, v149_0, v14_0, v150_0, v151_0, v152_0, v153_0, v154_0, v155_0, v156_0, v157_0, v158_0, v159_0, v15_0, v160_0, v161_0, v162_0, v163_0, v164_0, v165_0, v166_0, v167_0, v168_0, v169_0, v16_0, v170_0, v171_0, v172_0, v173_0, v174_0, v175_0, v176_0, v177_0, v178_0, v179_0, v17_0, v180_0, v181_0, v182_0, v183_0, v184_0, v185_0, v186_0, v187_0, v188_0, v189_0, v18_0, v190_0, v191_0, v192_0, v193_0, v194_0, v195_0, v196_0, v197_0, v198_0, v199_0, v19_0, v1_0, v200_0, v201_0, v202_0, v203_0, v204_0, v205_0, v206_0, v207_0, v208_0, v209_0, v20_0, v210_0, v211_0, v212_0, v213_0, v214_0, v215_0, v216_0, v217_0, v218_0, v219_0, v21_0, v220_0, v221_0, v222_0, v223_0, v224_0, v225_0, v226_0, v227_0, v228_0, v229_0, v22_0, v230_0, v231_0, v232_0, v233_0, v234_0, v235_0, v236_0, v237_0, v23_0, v24_0, v25_0, v26_0, v27_0, v28_0, v29_0, v2_0, v30_0, v31_0, v32_0, v33_0, v34_0, v35_0, v36_0, v37_0, v38_0, v39_0, v3_0, v40_0, v41_0, v42_0, v43_0, v44_0, v45_0, v46_0, v47_0, v48_0, v49_0, v4_0, v50_0, v51_0, v52_0, v53_0, v54_0, v55_0, v56_0, v57_0, v58_0, v59_0, v5_0, v60_0, v61_0, v62_0, v63_0, v64_0, v65_0, v66_0, v67_0, v68_0, v69_0, v6_0, v70_0, v71_0, v72_0, v73_0, v74_0, v75_0, v76_0, v77_0, v78_0, v79_0, v7_0, v80_0, v81_0, v82_0, v83_0, v84_0, v85_0, v86_0, v87_0, v88_0, v89_0, v8_0, v90_0, v91_0, v92_0, v93_0, v94_0, v95_0, v96_0, v97_0, v98_0, v99_0, v9_0;

  // Map n0..n7 to A[0..7], n8..n15 to B[0..7]
  assign n0 = A[0];
  assign n1 = A[1];
  assign n2 = A[2];
  assign n3 = A[3];
  assign n4 = A[4];
  assign n5 = A[5];
  assign n6 = A[6];
  assign n7 = A[7];
  assign n8 = B[0];
  assign n9 = B[1];
  assign n10 = B[2];
  assign n11 = B[3];
  assign n12 = B[4];
  assign n13 = B[5];
  assign n14 = B[6];
  assign n15 = B[7];

  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0001_ (
    .I(n2),
    .ZN(v0_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0002_ (
    .A1(n7),
    .A2(n10),
    .ZN(v1_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0003_ (
    .I(n3),
    .ZN(v2_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0004_ (
    .I(n4),
    .ZN(v3_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0005_ (
    .I(n11),
    .ZN(v4_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0006_ (
    .I(n15),
    .ZN(v5_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0007_ (
    .A1(n5),
    .A2(n11),
    .ZN(v6_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0008_ (
    .A1(v3_0),
    .A2(v4_0),
    .Z(v7_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0009_ (
    .I(n5),
    .ZN(v8_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0010_ (
    .I(n1),
    .ZN(v9_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0011_ (
    .I(n10),
    .ZN(v10_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0012_ (
    .I(v9_0),
    .ZN(v11_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0013_ (
    .A1(n5),
    .A2(n12),
    .ZN(v12_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0014_ (
    .A1(v7_0),
    .A2(v12_0),
    .Z(v13_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0015_ (
    .A1(n4),
    .A2(n12),
    .ZN(v14_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0016_ (
    .A1(v6_0),
    .A2(v14_0),
    .ZN(v15_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0017_ (
    .A1(v13_0),
    .A2(v15_0),
    .ZN(v16_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0018_ (
    .A1(n3),
    .A2(n13),
    .ZN(v17_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0019_ (
    .A1(v16_0),
    .A2(v17_0),
    .Z(v18_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0020_ (
    .A1(v16_0),
    .A2(v17_0),
    .ZN(v19_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0021_ (
    .I(n7),
    .ZN(v20_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0022_ (
    .I(n6),
    .ZN(v21_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0023_ (
    .A1(v20_0),
    .A2(v21_0),
    .Z(v22_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0024_ (
    .I(v19_0),
    .ZN(v23_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0025_ (
    .A1(n2),
    .A2(n14),
    .ZN(v24_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0026_ (
    .A1(v9_0),
    .A2(n15),
    .ZN(v25_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0027_ (
    .A1(v24_0),
    .A2(v25_0),
    .Z(v26_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0028_ (
    .A1(v3_0),
    .A2(v26_0),
    .ZN(v27_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0029_ (
    .I(v26_0),
    .ZN(v28_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0030_ (
    .A1(v3_0),
    .A2(v28_0),
    .Z(v29_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0031_ (
    .A1(v11_0),
    .A2(v29_0),
    .Z(v30_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0032_ (
    .A1(v10_0),
    .A2(v30_0),
    .Z(v31_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0033_ (
    .A1(v31_0),
    .A2(v31_0),
    .Z(v32_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0034_ (
    .I(v7_0),
    .ZN(v33_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0035_ (
    .A1(v32_0),
    .A2(v33_0),
    .Z(v34_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0036_ (
    .I(v23_0),
    .ZN(v35_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0037_ (
    .A1(n11),
    .A2(n6),
    .ZN(v36_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0038_ (
    .A1(v12_0),
    .A2(v36_0),
    .Z(v37_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0039_ (
    .I(v37_0),
    .ZN(v38_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0040_ (
    .A1(n4),
    .A2(n13),
    .ZN(v39_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0041_ (
    .A1(v38_0),
    .A2(v39_0),
    .Z(v40_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0042_ (
    .A1(v38_0),
    .A2(v39_0),
    .ZN(v41_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0043_ (
    .A1(v40_0),
    .A2(v41_0),
    .ZN(v42_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0044_ (
    .A1(v1_0),
    .A2(v20_0),
    .Z(v43_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0045_ (
    .I(v22_0),
    .ZN(v44_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0046_ (
    .A1(v43_0),
    .A2(v44_0),
    .Z(v45_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0047_ (
    .A1(v42_0),
    .A2(v45_0),
    .Z(v46_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0048_ (
    .A1(v46_0),
    .A2(v46_0),
    .Z(v47_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0049_ (
    .A1(v25_0),
    .A2(v24_0),
    .Z(v48_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0050_ (
    .A1(n3),
    .A2(n14),
    .ZN(v49_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0051_ (
    .A1(v0_0),
    .A2(n15),
    .ZN(v50_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0052_ (
    .A1(v49_0),
    .A2(v50_0),
    .Z(v51_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0053_ (
    .A1(v18_0),
    .A2(v13_0),
    .ZN(v52_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0054_ (
    .A1(v51_0),
    .A2(v52_0),
    .Z(v53_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0055_ (
    .I(v53_0),
    .ZN(v54_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0056_ (
    .A1(v48_0),
    .A2(v54_0),
    .ZN(v55_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0057_ (
    .I(v55_0),
    .ZN(v56_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0058_ (
    .A1(v47_0),
    .A2(v56_0),
    .Z(v57_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0059_ (
    .A1(v47_0),
    .A2(v56_0),
    .ZN(v58_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0060_ (
    .A1(v57_0),
    .A2(v58_0),
    .ZN(v59_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0061_ (
    .A1(v35_0),
    .A2(v59_0),
    .Z(v60_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0062_ (
    .A1(v27_0),
    .A2(v60_0),
    .Z(v61_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0063_ (
    .A1(v30_0),
    .A2(v10_0),
    .Z(v62_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0064_ (
    .A1(v30_0),
    .A2(v11_0),
    .ZN(v63_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0065_ (
    .A1(v62_0),
    .A2(v63_0),
    .ZN(v64_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0066_ (
    .A1(v61_0),
    .A2(v64_0),
    .Z(v65_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0067_ (
    .A1(v61_0),
    .A2(v64_0),
    .ZN(v66_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0068_ (
    .A1(v65_0),
    .A2(v66_0),
    .Z(v67_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0069_ (
    .A1(v33_0),
    .A2(v32_0),
    .Z(v68_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0070_ (
    .A1(v67_0),
    .A2(v68_0),
    .Z(v69_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0071_ (
    .A1(v60_0),
    .A2(v27_0),
    .Z(v70_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0072_ (
    .A1(v60_0),
    .A2(v35_0),
    .ZN(v71_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0073_ (
    .A1(v70_0),
    .A2(v71_0),
    .ZN(v72_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0074_ (
    .A1(v54_0),
    .A2(v48_0),
    .Z(v73_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0075_ (
    .A1(v52_0),
    .A2(v51_0),
    .ZN(v74_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0076_ (
    .A1(v73_0),
    .A2(v74_0),
    .ZN(v75_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0077_ (
    .A1(n4),
    .A2(n14),
    .ZN(v76_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0078_ (
    .A1(v2_0),
    .A2(n15),
    .ZN(v77_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0079_ (
    .A1(v76_0),
    .A2(v77_0),
    .Z(v78_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0080_ (
    .A1(n12),
    .A2(n6),
    .ZN(v79_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0081_ (
    .A1(v6_0),
    .A2(v79_0),
    .Z(v80_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0082_ (
    .A1(v40_0),
    .A2(v80_0),
    .ZN(v81_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0083_ (
    .A1(v78_0),
    .A2(v81_0),
    .Z(v82_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0084_ (
    .I(v82_0),
    .ZN(v83_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0085_ (
    .A1(v50_0),
    .A2(v49_0),
    .Z(v84_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0086_ (
    .A1(v83_0),
    .A2(v84_0),
    .Z(v85_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0087_ (
    .A1(v83_0),
    .A2(v84_0),
    .ZN(v86_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0088_ (
    .A1(v85_0),
    .A2(v86_0),
    .ZN(v87_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0089_ (
    .A1(v45_0),
    .A2(v46_0),
    .ZN(v88_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0090_ (
    .I(v88_0),
    .ZN(v89_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0091_ (
    .I(v20_0),
    .ZN(v90_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0092_ (
    .I(v90_0),
    .ZN(v91_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0093_ (
    .A1(n11),
    .A2(n7),
    .ZN(v92_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0094_ (
    .A1(v79_0),
    .A2(v92_0),
    .Z(v93_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0095_ (
    .I(v93_0),
    .ZN(v94_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0096_ (
    .A1(n5),
    .A2(n13),
    .ZN(v95_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0097_ (
    .A1(v94_0),
    .A2(v95_0),
    .Z(v96_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0098_ (
    .A1(v94_0),
    .A2(v95_0),
    .ZN(v97_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0099_ (
    .A1(v96_0),
    .A2(v97_0),
    .Z(v98_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0100_ (
    .I(v98_0),
    .ZN(v99_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0101_ (
    .A1(v91_0),
    .A2(v99_0),
    .Z(v100_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0102_ (
    .A1(v89_0),
    .A2(v100_0),
    .Z(v101_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0103_ (
    .A1(v89_0),
    .A2(v99_0),
    .ZN(v102_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0104_ (
    .A1(v101_0),
    .A2(v102_0),
    .ZN(v103_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0105_ (
    .A1(v87_0),
    .A2(v103_0),
    .Z(v104_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0106_ (
    .I(v57_0),
    .ZN(v105_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0107_ (
    .A1(v104_0),
    .A2(v105_0),
    .Z(v106_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0108_ (
    .A1(v75_0),
    .A2(v106_0),
    .Z(v107_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0109_ (
    .A1(v72_0),
    .A2(v107_0),
    .Z(v108_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0110_ (
    .A1(v68_0),
    .A2(v67_0),
    .ZN(v109_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0111_ (
    .A1(v109_0),
    .A2(v66_0),
    .ZN(v110_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0112_ (
    .A1(v108_0),
    .A2(v110_0),
    .Z(v111_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0113_ (
    .A1(v81_0),
    .A2(v78_0),
    .ZN(v112_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0114_ (
    .A1(v85_0),
    .A2(v112_0),
    .ZN(v113_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0115_ (
    .A1(v103_0),
    .A2(v87_0),
    .Z(v114_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0116_ (
    .A1(v114_0),
    .A2(v102_0),
    .ZN(v115_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0117_ (
    .A1(n5),
    .A2(n14),
    .ZN(v116_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0118_ (
    .A1(v3_0),
    .A2(n15),
    .ZN(v117_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0119_ (
    .A1(v116_0),
    .A2(v117_0),
    .Z(v118_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0120_ (
    .A1(v79_0),
    .A2(v92_0),
    .Z(v119_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0121_ (
    .A1(v96_0),
    .A2(v119_0),
    .ZN(v120_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0122_ (
    .A1(v118_0),
    .A2(v120_0),
    .Z(v121_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0123_ (
    .I(v121_0),
    .ZN(v122_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0124_ (
    .A1(v77_0),
    .A2(v76_0),
    .Z(v123_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0125_ (
    .A1(v122_0),
    .A2(v123_0),
    .Z(v124_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0126_ (
    .A1(v122_0),
    .A2(v123_0),
    .ZN(v125_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0127_ (
    .A1(v124_0),
    .A2(v125_0),
    .Z(v126_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0128_ (
    .A1(v90_0),
    .A2(v98_0),
    .ZN(v127_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0129_ (
    .I(v127_0),
    .ZN(v128_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0130_ (
    .I(v92_0),
    .ZN(v129_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0131_ (
    .A1(v129_0),
    .A2(n12),
    .ZN(v130_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0132_ (
    .A1(n12),
    .A2(n7),
    .ZN(v131_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0133_ (
    .A1(v92_0),
    .A2(v131_0),
    .ZN(v132_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0134_ (
    .A1(v130_0),
    .A2(v132_0),
    .ZN(v133_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0135_ (
    .A1(n13),
    .A2(n6),
    .ZN(v134_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0136_ (
    .A1(v133_0),
    .A2(v134_0),
    .Z(v135_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0137_ (
    .A1(v133_0),
    .A2(v134_0),
    .ZN(v136_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0138_ (
    .A1(v135_0),
    .A2(v136_0),
    .Z(v137_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0139_ (
    .I(v137_0),
    .ZN(v138_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0140_ (
    .A1(v138_0),
    .A2(v91_0),
    .Z(v139_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0141_ (
    .A1(v128_0),
    .A2(v139_0),
    .Z(v140_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0142_ (
    .A1(v128_0),
    .A2(v139_0),
    .ZN(v141_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0143_ (
    .A1(v140_0),
    .A2(v141_0),
    .Z(v142_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0144_ (
    .A1(v126_0),
    .A2(v142_0),
    .Z(v143_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0145_ (
    .A1(v115_0),
    .A2(v143_0),
    .Z(v144_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0146_ (
    .A1(v113_0),
    .A2(v144_0),
    .Z(v145_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0147_ (
    .A1(v106_0),
    .A2(v75_0),
    .ZN(v146_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0148_ (
    .A1(v105_0),
    .A2(v104_0),
    .ZN(v147_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0149_ (
    .A1(v146_0),
    .A2(v147_0),
    .ZN(v148_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0150_ (
    .A1(v145_0),
    .A2(v148_0),
    .Z(v149_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0151_ (
    .A1(v145_0),
    .A2(v148_0),
    .ZN(v150_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0152_ (
    .A1(v149_0),
    .A2(v150_0),
    .Z(v151_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0153_ (
    .A1(v110_0),
    .A2(v108_0),
    .ZN(v152_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0154_ (
    .A1(v107_0),
    .A2(v72_0),
    .ZN(v153_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0155_ (
    .A1(v152_0),
    .A2(v153_0),
    .ZN(v154_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0156_ (
    .A1(v151_0),
    .A2(v154_0),
    .Z(v155_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0157_ (
    .A1(v144_0),
    .A2(v113_0),
    .ZN(v156_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0158_ (
    .A1(v143_0),
    .A2(v115_0),
    .ZN(v157_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0159_ (
    .A1(v156_0),
    .A2(v157_0),
    .ZN(v158_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0160_ (
    .A1(v122_0),
    .A2(v118_0),
    .ZN(v159_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0161_ (
    .A1(v124_0),
    .A2(v159_0),
    .ZN(v160_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0162_ (
    .A1(v142_0),
    .A2(v126_0),
    .ZN(v161_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0163_ (
    .A1(v161_0),
    .A2(v141_0),
    .ZN(v162_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0164_ (
    .A1(n6),
    .A2(n14),
    .ZN(v163_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0165_ (
    .A1(v8_0),
    .A2(n15),
    .ZN(v164_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0166_ (
    .A1(v163_0),
    .A2(v164_0),
    .Z(v165_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0167_ (
    .A1(v135_0),
    .A2(v130_0),
    .ZN(v166_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0168_ (
    .A1(v165_0),
    .A2(v166_0),
    .Z(v167_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0169_ (
    .I(v167_0),
    .ZN(v168_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0170_ (
    .A1(v117_0),
    .A2(v116_0),
    .Z(v169_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0171_ (
    .A1(v168_0),
    .A2(v169_0),
    .Z(v170_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0172_ (
    .A1(v168_0),
    .A2(v169_0),
    .ZN(v171_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0173_ (
    .A1(v170_0),
    .A2(v171_0),
    .Z(v172_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0174_ (
    .A1(v90_0),
    .A2(v137_0),
    .ZN(v173_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0175_ (
    .I(v173_0),
    .ZN(v174_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0176_ (
    .A1(n13),
    .A2(n7),
    .ZN(v175_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0177_ (
    .A1(v175_0),
    .A2(v133_0),
    .Z(v176_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0178_ (
    .I(v176_0),
    .ZN(v177_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0179_ (
    .A1(v177_0),
    .A2(v91_0),
    .Z(v178_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0180_ (
    .A1(v174_0),
    .A2(v178_0),
    .Z(v179_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0181_ (
    .A1(v174_0),
    .A2(v178_0),
    .ZN(v180_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0182_ (
    .A1(v179_0),
    .A2(v180_0),
    .Z(v181_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0183_ (
    .A1(v172_0),
    .A2(v181_0),
    .Z(v182_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0184_ (
    .A1(v162_0),
    .A2(v182_0),
    .Z(v183_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0185_ (
    .A1(v160_0),
    .A2(v183_0),
    .Z(v184_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0186_ (
    .A1(v158_0),
    .A2(v184_0),
    .Z(v185_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0187_ (
    .A1(v152_0),
    .A2(v155_0),
    .ZN(v186_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0188_ (
    .A1(v186_0),
    .A2(v149_0),
    .Z(v187_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0189_ (
    .A1(v185_0),
    .A2(v187_0),
    .Z(v188_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0190_ (
    .A1(v166_0),
    .A2(v165_0),
    .ZN(v189_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0191_ (
    .A1(v170_0),
    .A2(v189_0),
    .ZN(v190_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0192_ (
    .A1(v181_0),
    .A2(v172_0),
    .ZN(v191_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0193_ (
    .A1(v191_0),
    .A2(v180_0),
    .ZN(v192_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0194_ (
    .A1(v133_0),
    .A2(v175_0),
    .Z(v193_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0195_ (
    .A1(v193_0),
    .A2(v130_0),
    .ZN(v194_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0196_ (
    .I(v194_0),
    .ZN(v195_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0197_ (
    .A1(n14),
    .A2(n7),
    .ZN(v196_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0198_ (
    .I(v196_0),
    .ZN(v197_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0199_ (
    .A1(v5_0),
    .A2(n6),
    .Z(v198_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0200_ (
    .A1(v197_0),
    .A2(v198_0),
    .Z(v199_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0201_ (
    .A1(v195_0),
    .A2(v199_0),
    .Z(v200_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0202_ (
    .A1(v195_0),
    .A2(v199_0),
    .ZN(v201_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0203_ (
    .A1(v200_0),
    .A2(v201_0),
    .Z(v202_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0204_ (
    .I(v202_0),
    .ZN(v203_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0205_ (
    .A1(v164_0),
    .A2(v163_0),
    .Z(v204_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0206_ (
    .A1(v203_0),
    .A2(v204_0),
    .Z(v205_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0207_ (
    .A1(v203_0),
    .A2(v204_0),
    .ZN(v206_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0208_ (
    .A1(v205_0),
    .A2(v206_0),
    .Z(v207_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0209_ (
    .A1(v90_0),
    .A2(v207_0),
    .Z(v208_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0210_ (
    .A1(v192_0),
    .A2(v208_0),
    .Z(v209_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0211_ (
    .A1(v190_0),
    .A2(v209_0),
    .Z(v210_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0212_ (
    .A1(v183_0),
    .A2(v160_0),
    .ZN(v211_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0213_ (
    .A1(v182_0),
    .A2(v162_0),
    .ZN(v212_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0214_ (
    .A1(v211_0),
    .A2(v212_0),
    .ZN(v213_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0215_ (
    .A1(v210_0),
    .A2(v213_0),
    .Z(v214_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0216_ (
    .A1(v210_0),
    .A2(v213_0),
    .ZN(v215_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0217_ (
    .A1(v214_0),
    .A2(v215_0),
    .Z(v216_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0218_ (
    .A1(v187_0),
    .A2(v185_0),
    .ZN(v217_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0219_ (
    .A1(v184_0),
    .A2(v158_0),
    .ZN(v218_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0220_ (
    .A1(v217_0),
    .A2(v218_0),
    .ZN(v219_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0221_ (
    .A1(v216_0),
    .A2(v219_0),
    .Z(v220_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0222_ (
    .A1(v205_0),
    .A2(v200_0),
    .ZN(v221_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0223_ (
    .A1(v198_0),
    .A2(v197_0),
    .ZN(v222_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0224_ (
    .A1(v5_0),
    .A2(n7),
    .Z(v223_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0225_ (
    .A1(v222_0),
    .A2(v223_0),
    .ZN(v224_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0226_ (
    .A1(v224_0),
    .A2(v194_0),
    .Z(v225_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0227_ (
    .A1(v225_0),
    .A2(v90_0),
    .Z(v226_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0228_ (
    .A1(v207_0),
    .A2(v90_0),
    .ZN(v227_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0229_ (
    .I(v227_0),
    .ZN(v228_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0230_ (
    .A1(v226_0),
    .A2(v228_0),
    .Z(v229_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0231_ (
    .A1(v221_0),
    .A2(v229_0),
    .Z(v230_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0232_ (
    .A1(v209_0),
    .A2(v190_0),
    .ZN(v231_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0233_ (
    .A1(v208_0),
    .A2(v192_0),
    .ZN(v232_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0234_ (
    .A1(v231_0),
    .A2(v232_0),
    .ZN(v233_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0235_ (
    .A1(v230_0),
    .A2(v233_0),
    .Z(v234_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0236_ (
    .A1(v219_0),
    .A2(v214_0),
    .ZN(v235_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0237_ (
    .A1(v235_0),
    .A2(v215_0),
    .ZN(v236_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0238_ (
    .A1(v234_0),
    .A2(v236_0),
    .Z(v237_0)
  );

  assign OUT[0] = v206_0;
  assign OUT[1] = v101_0;
  assign OUT[2] = v121_0;
  assign OUT[3] = v131_0;
  assign OUT[4] = v184_0;
  assign OUT[5] = v155_0;
  assign OUT[6] = n2;
  assign OUT[7] = v23_0;
  assign OUT[8] = v34_0;
  assign OUT[9] = v69_0;
  assign OUT[10] = v111_0;
  assign OUT[11] = v155_0;
  assign OUT[12] = v188_0;
  assign OUT[13] = v220_0;
  assign OUT[14] = v237_0;
  assign OUT[15] = v237_0;
endmodule
