# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3 ;
  ORIGIN  1.055000  1.055000 ;
  SIZE  3.880000 BY  3.880000 ;
  PIN C0
    PORT
      LAYER met2 ;
        RECT 0.000000 0.000000 0.610000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 0.610000 ;
        RECT 0.000000 1.160000 0.330000 1.440000 ;
        RECT 0.000000 1.440000 0.610000 1.770000 ;
        RECT 1.160000 0.000000 1.770000 0.330000 ;
        RECT 1.160000 1.440000 1.770000 1.770000 ;
        RECT 1.440000 0.330000 1.770000 0.610000 ;
        RECT 1.440000 1.160000 1.770000 1.440000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met2 ;
        RECT 0.000000 0.750000 1.770000 1.020000 ;
        RECT 0.470000 0.470000 1.300000 0.610000 ;
        RECT 0.470000 1.160000 1.300000 1.300000 ;
        RECT 0.750000 0.000000 1.020000 0.470000 ;
        RECT 0.750000 0.610000 1.020000 0.750000 ;
        RECT 0.750000 1.020000 1.020000 1.160000 ;
        RECT 0.750000 1.300000 1.020000 1.770000 ;
    END
  END C1
  PIN MET3
    PORT
      LAYER met3 ;
        RECT -1.055000 -1.055000 2.825000 2.825000 ;
    END
  END MET3
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 1.255000 1.190000 1.375000 1.445000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1.770000 1.770000 ;
    LAYER mcon ;
      RECT 0.080000 0.080000 0.250000 0.250000 ;
      RECT 0.080000 0.440000 0.250000 0.610000 ;
      RECT 0.080000 0.800000 0.250000 0.970000 ;
      RECT 0.080000 1.160000 0.250000 1.330000 ;
      RECT 0.080000 1.520000 0.250000 1.690000 ;
      RECT 0.440000 0.080000 0.610000 0.250000 ;
      RECT 0.440000 1.520000 0.610000 1.690000 ;
      RECT 0.800000 0.080000 0.970000 0.250000 ;
      RECT 0.800000 1.520000 0.970000 1.690000 ;
      RECT 1.160000 0.080000 1.330000 0.250000 ;
      RECT 1.160000 1.520000 1.330000 1.690000 ;
      RECT 1.520000 0.080000 1.690000 0.250000 ;
      RECT 1.520000 0.440000 1.690000 0.610000 ;
      RECT 1.520000 0.800000 1.690000 0.970000 ;
      RECT 1.520000 1.160000 1.690000 1.330000 ;
      RECT 1.520000 1.520000 1.690000 1.690000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1.770000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 1.440000 ;
      RECT 0.000000 1.440000 1.770000 1.770000 ;
      RECT 0.470000 0.470000 0.610000 0.750000 ;
      RECT 0.470000 0.750000 1.300000 1.020000 ;
      RECT 0.470000 1.020000 0.610000 1.300000 ;
      RECT 0.750000 0.470000 1.020000 0.750000 ;
      RECT 0.750000 1.020000 1.020000 1.300000 ;
      RECT 1.160000 0.470000 1.300000 0.750000 ;
      RECT 1.160000 1.020000 1.300000 1.300000 ;
      RECT 1.440000 0.330000 1.770000 1.440000 ;
    LAYER via ;
      RECT 0.035000 0.320000 0.295000 0.580000 ;
      RECT 0.035000 1.190000 0.295000 1.450000 ;
      RECT 0.320000 0.035000 0.580000 0.295000 ;
      RECT 0.320000 1.475000 0.580000 1.735000 ;
      RECT 0.470000 0.755000 0.730000 1.015000 ;
      RECT 0.755000 0.500000 1.015000 0.760000 ;
      RECT 0.755000 1.010000 1.015000 1.270000 ;
      RECT 1.040000 0.755000 1.300000 1.015000 ;
      RECT 1.190000 0.035000 1.450000 0.295000 ;
      RECT 1.190000 1.475000 1.450000 1.735000 ;
      RECT 1.475000 0.320000 1.735000 0.580000 ;
      RECT 1.475000 1.190000 1.735000 1.450000 ;
  END
END sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3
END LIBRARY
