* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 38
.param
+ sky130_fd_pr__nfet_01v8_lvt__toxe_mult = 1.0365
+ sky130_fd_pr__nfet_01v8_lvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_01v8_lvt__overlap_mult = 0.9632
+ sky130_fd_pr__nfet_01v8_lvt__ajunction_mult = 1.1229
+ sky130_fd_pr__nfet_01v8_lvt__pjunction_mult = 1.0009
+ sky130_fd_pr__nfet_01v8_lvt__lint_diff = -1.21275e-8
+ sky130_fd_pr__nfet_01v8_lvt__wint_diff = 2.252e-8
+ sky130_fd_pr__nfet_01v8_lvt__dlc_diff = -1.1228e-8
+ sky130_fd_pr__nfet_01v8_lvt__dwc_diff = 2.252e-8
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 000, W = 1.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_0 = -0.098172
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_0 = 0.0084685
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_0 = -0.0027071
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_0 = -0.17335
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_0 = 2.3712e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_0 = -8.8501e-21
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0 = 1.0585
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0 = -0.0025154
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 001, W = 1.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_1 = -0.090752
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_1 = 0.0070719
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_1 = -0.19831
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_1 = -0.0036953
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_1 = 7.0103e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_1 = 7.0368e-21
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1 = 0.47034
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1 = -0.0032454
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 002, W = 1.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2 = -0.0067259
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_2 = 0.0054653
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_2 = 0.0097562
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_2 = 0.042661
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_2 = -0.0038874
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_2 = 1.2427e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_2 = 1.7645e-20
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2 = 1.0266
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 003, W = 1.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3 = 1.713
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3 = 0.050867
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_3 = -0.013593
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_3 = 0.0012164
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_3 = -5.9367e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3 = 15330.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_3 = 1.6856e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 004, W = 1.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4 = 1.7318
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4 = 0.0083694
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_4 = -0.0099683
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_4 = -0.0014096
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_4 = -1.8383e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4 = 8402.2
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_4 = -7.5484e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 005, W = 1.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_5 = -2.0786e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5 = 1.2552
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5 = 0.010815
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_5 = 0.0053313
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_5 = -0.0061101
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_5 = -3.88e-11
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5 = -7222.9
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_5 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 006, W = 1.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_6 = -1.0226e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6 = 1.0513
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6 = -0.00281
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_6 = 0.0035231
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_6 = -0.0025486
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_6 = -1.0269e-11
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6 = 16049.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_6 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 007, W = 3.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_7 = 1.5569e-20
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7 = 0.92324
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7 = 1.1738e-5
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_7 = -0.10554
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_7 = 0.0059516
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_7 = -0.13065
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_7 = -0.00046542
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_7 = 2.4008e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 008, W = 3.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_8 = -0.13812
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_8 = -2.3907e-5
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_8 = 1.6561e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_8 = 1.1444e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8 = 0.43557
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8 = -0.0063361
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_8 = -0.090119
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_8 = 0.0044571
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 009, W = 3.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_9 = -0.023592
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_9 = -0.00084689
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_9 = -4.9665e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_9 = 4.2142e-20
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9 = 0.58545
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9 = -0.004977
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_9 = 0.010882
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_9 = 0.0070278
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 010, W = 3.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_10 = 3.6117e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_10 = 1.7405e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_10 = -0.0013865
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10 = 15652.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10 = 0.00059676
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10 = 1.5258
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_10 = -0.016009
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 011, W = 3.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_11 = -0.010413
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_11 = -5.3155e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_11 = 1.2312e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_11 = 0.00048662
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11 = 13003.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11 = 0.0075839
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11 = 1.5575
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 012, W = 3.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_12 = 0.0039021
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_12 = -1.7494e-10
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_12 = 1.1247e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_12 = -0.0051672
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12 = 12431.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12 = 0.0051902
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12 = 1.1333
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_12 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 013, W = 3.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_13 = 0.0104
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_13 = -2.3811e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_13 = 1.0065e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_13 = 0.00033753
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13 = 14111.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13 = -0.00056285
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13 = 1.279
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_13 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 014, W = 5.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14 = 0.74776
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_14 = 0.0035119
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_14 = 1.6765e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_14 = 1.0295e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_14 = -0.099705
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_14 = -0.14352
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_14 = 0.00063825
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14 = -0.0054958
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 015, W = 5.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15 = -0.0017086
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15 = 0.73762
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_15 = -0.0057065
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_15 = -1.1419e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_15 = 9.3017e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_15 = -0.024227
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_15 = -0.082489
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_15 = 0.00019125
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 016, W = 5.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_16 = -0.080836
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_16 = 8.6876e-6
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16 = -0.0065941
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16 = 0.183
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_16 = 0.010658
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_16 = 5.1068e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_16 = 9.1242e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_16 = 0.013681
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 017, W = 5.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_17 = 0.0012046
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17 = 18998.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17 = 0.012659
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17 = 1.5543
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_17 = -0.018618
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_17 = -1.1738e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_17 = 2.5304e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 018, W = 5.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_18 = -5.424e-5
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18 = 6404.6
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18 = 0.018672
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18 = 1.3805
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_18 = -0.0095611
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_18 = -1.1464e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_18 = 1.2294e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 019, W = 5.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_19 = -7.353e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_19 = -0.0062942
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19 = 4955.1
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19 = -0.0078181
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19 = 1.283
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_19 = 0.0015267
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_19 = -5.7263e-11
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 020, W = 5.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_20 = -4.4186e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_20 = 2.0425e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_20 = 0.0020151
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20 = 11267.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20 = -0.00695
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20 = 0.93542
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_20 = 0.0041501
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 021, W = 7.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_21 = -1.3594e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_21 = 1.2003e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_21 = -0.064846
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_21 = -0.086538
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_21 = 0.00086992
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21 = 0.00054786
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21 = 0.77157
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_21 = -0.0026262
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 022, W = 7.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_22 = 0.0093323
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_22 = 1.6144e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_22 = 9.0254e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_22 = -0.052987
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_22 = -0.13444
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_22 = 0.00026651
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22 = -0.0041849
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22 = 0.54697
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 023, W = 7.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_23 = 0.0083777
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_23 = -2.0667e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_23 = 1.6404e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_23 = 0.0085815
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_23 = -0.019173
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_23 = 0.00054736
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23 = -0.0040589
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23 = 0.44065
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_23 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 024, W = 7.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_24 = -0.010133
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_24 = 1.4921e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_24 = -1.0826e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_24 = -0.0025741
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24 = 10821.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24 = -0.005643
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24 = 1.5902
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_24 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 025, W = 7.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25 = 1.3778
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_25 = -0.0041947
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_25 = 1.2222e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_25 = 2.2389e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_25 = 0.00098004
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25 = 14700.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25 = -0.0043489
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 026, W = 7.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26 = -0.0096463
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26 = 1.3279
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_26 = 0.0030222
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_26 = 3.6823e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_26 = 8.5274e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_26 = -0.0037483
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26 = 20625.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 027, W = 7.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_27 = 0.0014067
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27 = -1191.1
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27 = -0.0016752
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27 = 1.1766
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_27 = 0.004209
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_27 = -4.7665e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_27 = 1.7991e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 028, W = 0.42, L = 1.0
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_28 = -0.010195
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28 = -0.0092111
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28 = 0.90829
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_28 = 1.1349e-7
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_28 = 4.3235e-8
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_28 = 0.0032889
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_28 = 4.8417e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_28 = -2.9607e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 029, W = 0.42, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_29 = -0.0014056
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29 = 32108.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29 = 0.053117
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29 = 1.7096
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_29 = -0.014845
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_29 = 2.011e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_29 = -1.5106e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 030, W = 0.42, L = 0.18
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_30 = 1.4221e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_30 = -0.00018398
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30 = 12891.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30 = 0.0079808
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30 = 1.5134
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_30 = -0.007809
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_30 = -2.8719e-12
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 031, W = 0.55, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_31 = 5.5377e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_31 = -6.1658e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_31 = -0.0013544
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31 = 26129.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31 = 0.068002
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31 = 1.9341
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_31 = -0.011808
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 032, W = 0.64, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_32 = -7.0929e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_32 = -3.2957e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_32 = -0.0022473
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32 = 9062.8
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32 = 0.054854
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32 = 2.1603
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_32 = -0.013718
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 033, W = 0.84, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_33 = -0.014456
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_33 = 8.4874e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_33 = -2.0231e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_33 = -0.001638
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33 = 7361.5
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33 = 0.061442
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33 = 2.0665
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 034, W = 1.65, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_34 = -0.011173
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_34 = 2.3351e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_34 = -8.8282e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_34 = -0.0020995
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34 = 14209.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34 = 0.028282
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34 = 1.3017
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_34 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 035, W = 3.01, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_35 = -0.016762
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_35 = 1.6664e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_35 = 1.0295e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_35 = -0.001361
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35 = 12105.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35 = 0.0027356
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35 = 1.5776
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_35 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 036, W = 5.05, L = 0.15
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36 = 1.7146
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_36 = -0.018098
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_36 = -5.6502e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_36 = 2.684e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_36 = 0.0013112
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36 = 19178.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36 = 0.014455
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 037, W = 5.05, L = 0.25
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37 = -0.0030604
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37 = 1.3479
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_37 = 0.0017424
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_37 = 5.0e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_37 = -1.2547e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_37 = -0.005
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37 = 7446.6
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
