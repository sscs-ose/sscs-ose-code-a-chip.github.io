* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope= .80e-2
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1= 2.05e-2 $ All W with L=0.5um
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2= 1.00e-2 $ W=3 L=1 um All W with L=0.8um & L=0.6um
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3= 0.67e-2 $ All W with L=4.0um
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope=0.000  $ All devices
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope=0.13  $ All devices
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope=0.12  $ All devices
.param sky130_fd_pr__nfet_g5v0d10v5__lint_slope=0.0  $ All devices
.param sky130_fd_pr__nfet_g5v0d10v5__wint_slope=0.0  $ All devices
