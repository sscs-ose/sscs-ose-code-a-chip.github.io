* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope= 1.20e-2
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1= 2.00e-2
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2= 2.30e-2
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3= 1.40e-2
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope=0.00e-2  $ All devices
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope=0.009  $ All devices
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope=0.02  $ All devices
.param sky130_fd_pr__pfet_g5v0d10v5__lint_slope=0.0  $ All devices
.param sky130_fd_pr__pfet_g5v0d10v5__wint_slope=0.0  $ All devices
