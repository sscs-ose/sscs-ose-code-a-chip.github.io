MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 25.07 BY 35.03 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.18 2.78 10.46 13.18 ;
      LAYER M3 ;
        RECT 13.62 2.78 13.9 8.98 ;
      LAYER M3 ;
        RECT 10.18 6.115 10.46 6.485 ;
      LAYER M2 ;
        RECT 10.32 6.16 13.76 6.44 ;
      LAYER M3 ;
        RECT 13.62 6.115 13.9 6.485 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 19.64 14.54 19.92 26.62 ;
      LAYER M2 ;
        RECT 13.16 27.16 22.96 27.44 ;
      LAYER M3 ;
        RECT 19.64 26.46 19.92 27.3 ;
      LAYER M2 ;
        RECT 19.62 27.16 19.94 27.44 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 2.8 19.52 3.08 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 4.56 2.8 7.48 3.08 ;
    END
  END VINP
  OBS 
  LAYER M2 ;
        RECT 16.6 7 19.52 7.28 ;
  LAYER M3 ;
        RECT 20.07 10.34 20.35 22.42 ;
  LAYER M3 ;
        RECT 14.05 13.7 14.33 24.1 ;
  LAYER M2 ;
        RECT 19.35 7 20.21 7.28 ;
  LAYER M3 ;
        RECT 20.07 7.14 20.35 10.5 ;
  LAYER M3 ;
        RECT 20.07 13.675 20.35 14.045 ;
  LAYER M4 ;
        RECT 14.19 13.46 20.21 14.26 ;
  LAYER M3 ;
        RECT 14.05 13.675 14.33 14.045 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M3 ;
        RECT 14.05 13.675 14.33 14.045 ;
  LAYER M4 ;
        RECT 14.025 13.46 14.355 14.26 ;
  LAYER M3 ;
        RECT 20.07 13.675 20.35 14.045 ;
  LAYER M4 ;
        RECT 20.045 13.46 20.375 14.26 ;
  LAYER M2 ;
        RECT 20.05 7 20.37 7.28 ;
  LAYER M3 ;
        RECT 20.07 6.98 20.35 7.3 ;
  LAYER M3 ;
        RECT 14.05 13.675 14.33 14.045 ;
  LAYER M4 ;
        RECT 14.025 13.46 14.355 14.26 ;
  LAYER M3 ;
        RECT 20.07 13.675 20.35 14.045 ;
  LAYER M4 ;
        RECT 20.045 13.46 20.375 14.26 ;
  LAYER M2 ;
        RECT 4.56 7 7.48 7.28 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 22.42 ;
  LAYER M3 ;
        RECT 9.75 13.7 10.03 24.1 ;
  LAYER M2 ;
        RECT 3.87 7 4.73 7.28 ;
  LAYER M3 ;
        RECT 3.73 7.14 4.01 10.5 ;
  LAYER M3 ;
        RECT 3.73 13.675 4.01 14.045 ;
  LAYER M4 ;
        RECT 3.87 13.46 9.89 14.26 ;
  LAYER M3 ;
        RECT 9.75 13.675 10.03 14.045 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M3 ;
        RECT 3.73 13.675 4.01 14.045 ;
  LAYER M4 ;
        RECT 3.705 13.46 4.035 14.26 ;
  LAYER M3 ;
        RECT 9.75 13.675 10.03 14.045 ;
  LAYER M4 ;
        RECT 9.725 13.46 10.055 14.26 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M3 ;
        RECT 3.73 13.675 4.01 14.045 ;
  LAYER M4 ;
        RECT 3.705 13.46 4.035 14.26 ;
  LAYER M3 ;
        RECT 9.75 13.675 10.03 14.045 ;
  LAYER M4 ;
        RECT 9.725 13.46 10.055 14.26 ;
  LAYER M2 ;
        RECT 4.13 6.58 7.91 6.86 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 13.18 ;
  LAYER M2 ;
        RECT 16.17 6.58 19.95 6.86 ;
  LAYER M2 ;
        RECT 0.69 27.58 11.35 27.86 ;
  LAYER M2 ;
        RECT 12.73 27.58 23.39 27.86 ;
  LAYER M2 ;
        RECT 7.74 6.58 8.6 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.72 8.74 7.56 ;
  LAYER M2 ;
        RECT 8.6 7.42 13.33 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M2 ;
        RECT 13.33 7.42 15.48 7.7 ;
  LAYER M1 ;
        RECT 15.355 6.72 15.605 7.56 ;
  LAYER M2 ;
        RECT 15.48 6.58 16.34 6.86 ;
  LAYER M3 ;
        RECT 13.19 13.02 13.47 16.8 ;
  LAYER M2 ;
        RECT 8.6 16.66 13.33 16.94 ;
  LAYER M3 ;
        RECT 8.46 16.8 8.74 27.72 ;
  LAYER M2 ;
        RECT 8.44 27.58 8.76 27.86 ;
  LAYER M2 ;
        RECT 11.18 27.58 12.9 27.86 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 8.44 16.66 8.76 16.94 ;
  LAYER M3 ;
        RECT 8.46 16.64 8.74 16.96 ;
  LAYER M2 ;
        RECT 8.44 27.58 8.76 27.86 ;
  LAYER M3 ;
        RECT 8.46 27.56 8.74 27.88 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 13.17 16.66 13.49 16.94 ;
  LAYER M3 ;
        RECT 13.19 16.64 13.47 16.96 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 8.44 16.66 8.76 16.94 ;
  LAYER M3 ;
        RECT 8.46 16.64 8.74 16.96 ;
  LAYER M2 ;
        RECT 8.44 27.58 8.76 27.86 ;
  LAYER M3 ;
        RECT 8.46 27.56 8.74 27.88 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 13.17 16.66 13.49 16.94 ;
  LAYER M3 ;
        RECT 13.19 16.64 13.47 16.96 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 8.44 16.66 8.76 16.94 ;
  LAYER M3 ;
        RECT 8.46 16.64 8.74 16.96 ;
  LAYER M2 ;
        RECT 8.44 27.58 8.76 27.86 ;
  LAYER M3 ;
        RECT 8.46 27.56 8.74 27.88 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 13.17 16.66 13.49 16.94 ;
  LAYER M3 ;
        RECT 13.19 16.64 13.47 16.96 ;
  LAYER M1 ;
        RECT 15.355 6.635 15.605 6.805 ;
  LAYER M2 ;
        RECT 15.31 6.58 15.65 6.86 ;
  LAYER M1 ;
        RECT 15.355 7.475 15.605 7.645 ;
  LAYER M2 ;
        RECT 15.31 7.42 15.65 7.7 ;
  LAYER M2 ;
        RECT 8.44 6.58 8.76 6.86 ;
  LAYER M3 ;
        RECT 8.46 6.56 8.74 6.88 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 8.44 16.66 8.76 16.94 ;
  LAYER M3 ;
        RECT 8.46 16.64 8.74 16.96 ;
  LAYER M2 ;
        RECT 8.44 27.58 8.76 27.86 ;
  LAYER M3 ;
        RECT 8.46 27.56 8.74 27.88 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 13.17 16.66 13.49 16.94 ;
  LAYER M3 ;
        RECT 13.19 16.64 13.47 16.96 ;
  LAYER M3 ;
        RECT 4.16 14.54 4.44 26.62 ;
  LAYER M3 ;
        RECT 5.45 27.14 5.73 31.66 ;
  LAYER M2 ;
        RECT 13.16 31.36 22.96 31.64 ;
  LAYER M3 ;
        RECT 4.16 26.46 4.44 26.88 ;
  LAYER M2 ;
        RECT 4.3 26.74 5.59 27.02 ;
  LAYER M3 ;
        RECT 5.45 26.88 5.73 27.3 ;
  LAYER M3 ;
        RECT 5.45 31.315 5.73 31.685 ;
  LAYER M4 ;
        RECT 5.59 31.1 11.61 31.9 ;
  LAYER M3 ;
        RECT 11.47 31.379 11.75 31.621 ;
  LAYER M2 ;
        RECT 11.61 31.36 13.33 31.64 ;
  LAYER M2 ;
        RECT 4.14 26.74 4.46 27.02 ;
  LAYER M3 ;
        RECT 4.16 26.72 4.44 27.04 ;
  LAYER M2 ;
        RECT 5.43 26.74 5.75 27.02 ;
  LAYER M3 ;
        RECT 5.45 26.72 5.73 27.04 ;
  LAYER M2 ;
        RECT 4.14 26.74 4.46 27.02 ;
  LAYER M3 ;
        RECT 4.16 26.72 4.44 27.04 ;
  LAYER M2 ;
        RECT 5.43 26.74 5.75 27.02 ;
  LAYER M3 ;
        RECT 5.45 26.72 5.73 27.04 ;
  LAYER M2 ;
        RECT 4.14 26.74 4.46 27.02 ;
  LAYER M3 ;
        RECT 4.16 26.72 4.44 27.04 ;
  LAYER M2 ;
        RECT 5.43 26.74 5.75 27.02 ;
  LAYER M3 ;
        RECT 5.45 26.72 5.73 27.04 ;
  LAYER M2 ;
        RECT 11.45 31.36 11.77 31.64 ;
  LAYER M3 ;
        RECT 11.47 31.34 11.75 31.66 ;
  LAYER M3 ;
        RECT 5.45 31.315 5.73 31.685 ;
  LAYER M4 ;
        RECT 5.425 31.1 5.755 31.9 ;
  LAYER M3 ;
        RECT 11.47 31.315 11.75 31.685 ;
  LAYER M4 ;
        RECT 11.445 31.1 11.775 31.9 ;
  LAYER M2 ;
        RECT 4.14 26.74 4.46 27.02 ;
  LAYER M3 ;
        RECT 4.16 26.72 4.44 27.04 ;
  LAYER M2 ;
        RECT 5.43 26.74 5.75 27.02 ;
  LAYER M3 ;
        RECT 5.45 26.72 5.73 27.04 ;
  LAYER M3 ;
        RECT 5.45 31.315 5.73 31.685 ;
  LAYER M4 ;
        RECT 5.425 31.1 5.755 31.9 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.72 8.68 10.92 8.96 ;
  LAYER M2 ;
        RECT 9.72 12.88 10.92 13.16 ;
  LAYER M2 ;
        RECT 9.29 12.46 11.35 12.74 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.29 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M3 ;
        RECT 10.18 2.78 10.46 13.18 ;
  LAYER M3 ;
        RECT 9.75 0.68 10.03 12.76 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M1 ;
        RECT 14.925 17.555 15.175 18.565 ;
  LAYER M1 ;
        RECT 14.925 19.655 15.175 23.185 ;
  LAYER M1 ;
        RECT 14.925 23.435 15.175 24.445 ;
  LAYER M1 ;
        RECT 14.925 25.535 15.175 26.545 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 15.355 19.655 15.605 23.185 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 17.305 ;
  LAYER M1 ;
        RECT 14.495 19.655 14.745 23.185 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 17.305 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 19.655 14.315 23.185 ;
  LAYER M1 ;
        RECT 14.065 23.435 14.315 24.445 ;
  LAYER M1 ;
        RECT 14.065 25.535 14.315 26.545 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 13.635 19.655 13.885 23.185 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 17.305 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 19.655 13.455 23.185 ;
  LAYER M1 ;
        RECT 13.205 23.435 13.455 24.445 ;
  LAYER M1 ;
        RECT 13.205 25.535 13.455 26.545 ;
  LAYER M1 ;
        RECT 12.775 13.775 13.025 17.305 ;
  LAYER M1 ;
        RECT 12.775 19.655 13.025 23.185 ;
  LAYER M2 ;
        RECT 13.16 17.92 15.22 18.2 ;
  LAYER M2 ;
        RECT 13.16 13.72 15.22 14 ;
  LAYER M2 ;
        RECT 12.73 14.14 15.65 14.42 ;
  LAYER M2 ;
        RECT 13.16 23.8 15.22 24.08 ;
  LAYER M2 ;
        RECT 13.16 19.6 15.22 19.88 ;
  LAYER M2 ;
        RECT 12.73 20.02 15.65 20.3 ;
  LAYER M2 ;
        RECT 13.16 25.9 15.22 26.18 ;
  LAYER M3 ;
        RECT 14.05 13.7 14.33 24.1 ;
  LAYER M3 ;
        RECT 13.62 14.12 13.9 26.2 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 17.305 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 19.655 9.155 23.185 ;
  LAYER M1 ;
        RECT 8.905 23.435 9.155 24.445 ;
  LAYER M1 ;
        RECT 8.905 25.535 9.155 26.545 ;
  LAYER M1 ;
        RECT 8.475 13.775 8.725 17.305 ;
  LAYER M1 ;
        RECT 8.475 19.655 8.725 23.185 ;
  LAYER M1 ;
        RECT 9.335 13.775 9.585 17.305 ;
  LAYER M1 ;
        RECT 9.335 19.655 9.585 23.185 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 17.305 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 19.655 10.015 23.185 ;
  LAYER M1 ;
        RECT 9.765 23.435 10.015 24.445 ;
  LAYER M1 ;
        RECT 9.765 25.535 10.015 26.545 ;
  LAYER M1 ;
        RECT 10.195 13.775 10.445 17.305 ;
  LAYER M1 ;
        RECT 10.195 19.655 10.445 23.185 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 17.305 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 19.655 10.875 23.185 ;
  LAYER M1 ;
        RECT 10.625 23.435 10.875 24.445 ;
  LAYER M1 ;
        RECT 10.625 25.535 10.875 26.545 ;
  LAYER M1 ;
        RECT 11.055 13.775 11.305 17.305 ;
  LAYER M1 ;
        RECT 11.055 19.655 11.305 23.185 ;
  LAYER M2 ;
        RECT 8.86 17.92 10.92 18.2 ;
  LAYER M2 ;
        RECT 8.86 13.72 10.92 14 ;
  LAYER M2 ;
        RECT 8.43 14.14 11.35 14.42 ;
  LAYER M2 ;
        RECT 8.86 23.8 10.92 24.08 ;
  LAYER M2 ;
        RECT 8.86 19.6 10.92 19.88 ;
  LAYER M2 ;
        RECT 8.43 20.02 11.35 20.3 ;
  LAYER M2 ;
        RECT 8.86 25.9 10.92 26.18 ;
  LAYER M3 ;
        RECT 9.75 13.7 10.03 24.1 ;
  LAYER M3 ;
        RECT 10.18 14.12 10.46 26.2 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M2 ;
        RECT 13.16 12.88 14.36 13.16 ;
  LAYER M2 ;
        RECT 13.16 8.68 14.36 8.96 ;
  LAYER M2 ;
        RECT 12.73 12.46 14.79 12.74 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 14.36 3.08 ;
  LAYER M2 ;
        RECT 12.73 6.58 14.79 6.86 ;
  LAYER M2 ;
        RECT 13.16 0.7 14.36 0.98 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 13.18 ;
  LAYER M3 ;
        RECT 13.62 2.78 13.9 8.98 ;
  LAYER M3 ;
        RECT 14.05 0.68 14.33 12.76 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 6.325 21.755 6.575 22.765 ;
  LAYER M1 ;
        RECT 6.325 17.135 6.575 20.665 ;
  LAYER M1 ;
        RECT 6.325 15.875 6.575 16.885 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 6.755 17.135 7.005 20.665 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M1 ;
        RECT 5.895 17.135 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 5.465 23.015 5.715 26.545 ;
  LAYER M1 ;
        RECT 5.465 21.755 5.715 22.765 ;
  LAYER M1 ;
        RECT 5.465 17.135 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.465 15.875 5.715 16.885 ;
  LAYER M1 ;
        RECT 5.465 11.255 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.465 9.995 5.715 11.005 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 8.905 ;
  LAYER M1 ;
        RECT 5.035 23.015 5.285 26.545 ;
  LAYER M1 ;
        RECT 5.035 17.135 5.285 20.665 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 26.545 ;
  LAYER M1 ;
        RECT 4.605 21.755 4.855 22.765 ;
  LAYER M1 ;
        RECT 4.605 17.135 4.855 20.665 ;
  LAYER M1 ;
        RECT 4.605 15.875 4.855 16.885 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M1 ;
        RECT 4.175 17.135 4.425 20.665 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 21.755 3.995 22.765 ;
  LAYER M1 ;
        RECT 3.745 17.135 3.995 20.665 ;
  LAYER M1 ;
        RECT 3.745 15.875 3.995 16.885 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M1 ;
        RECT 3.315 17.135 3.565 20.665 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 2.885 23.015 3.135 26.545 ;
  LAYER M1 ;
        RECT 2.885 21.755 3.135 22.765 ;
  LAYER M1 ;
        RECT 2.885 17.135 3.135 20.665 ;
  LAYER M1 ;
        RECT 2.885 15.875 3.135 16.885 ;
  LAYER M1 ;
        RECT 2.885 11.255 3.135 14.785 ;
  LAYER M1 ;
        RECT 2.885 9.995 3.135 11.005 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.905 ;
  LAYER M1 ;
        RECT 2.455 23.015 2.705 26.545 ;
  LAYER M1 ;
        RECT 2.455 17.135 2.705 20.665 ;
  LAYER M1 ;
        RECT 2.455 11.255 2.705 14.785 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 26.545 ;
  LAYER M1 ;
        RECT 2.025 21.755 2.275 22.765 ;
  LAYER M1 ;
        RECT 2.025 17.135 2.275 20.665 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.885 ;
  LAYER M1 ;
        RECT 2.025 11.255 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.905 ;
  LAYER M1 ;
        RECT 1.595 23.015 1.845 26.545 ;
  LAYER M1 ;
        RECT 1.595 17.135 1.845 20.665 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M1 ;
        RECT 1.165 23.015 1.415 26.545 ;
  LAYER M1 ;
        RECT 1.165 21.755 1.415 22.765 ;
  LAYER M1 ;
        RECT 1.165 17.135 1.415 20.665 ;
  LAYER M1 ;
        RECT 1.165 15.875 1.415 16.885 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.165 9.995 1.415 11.005 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 8.905 ;
  LAYER M1 ;
        RECT 0.735 23.015 0.985 26.545 ;
  LAYER M1 ;
        RECT 0.735 17.135 0.985 20.665 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 1.12 26.32 6.62 26.6 ;
  LAYER M2 ;
        RECT 1.12 22.12 6.62 22.4 ;
  LAYER M2 ;
        RECT 0.69 25.9 7.05 26.18 ;
  LAYER M2 ;
        RECT 1.12 20.44 6.62 20.72 ;
  LAYER M2 ;
        RECT 1.12 16.24 6.62 16.52 ;
  LAYER M2 ;
        RECT 0.69 20.02 7.05 20.3 ;
  LAYER M2 ;
        RECT 1.12 14.56 6.62 14.84 ;
  LAYER M2 ;
        RECT 1.12 10.36 6.62 10.64 ;
  LAYER M2 ;
        RECT 0.69 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 1.12 8.26 6.62 8.54 ;
  LAYER M3 ;
        RECT 4.16 14.54 4.44 26.62 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 22.42 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 26.2 ;
  LAYER M1 ;
        RECT 17.505 23.015 17.755 26.545 ;
  LAYER M1 ;
        RECT 17.505 21.755 17.755 22.765 ;
  LAYER M1 ;
        RECT 17.505 17.135 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.505 15.875 17.755 16.885 ;
  LAYER M1 ;
        RECT 17.505 11.255 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.505 9.995 17.755 11.005 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 8.905 ;
  LAYER M1 ;
        RECT 17.075 23.015 17.325 26.545 ;
  LAYER M1 ;
        RECT 17.075 17.135 17.325 20.665 ;
  LAYER M1 ;
        RECT 17.075 11.255 17.325 14.785 ;
  LAYER M1 ;
        RECT 17.935 23.015 18.185 26.545 ;
  LAYER M1 ;
        RECT 17.935 17.135 18.185 20.665 ;
  LAYER M1 ;
        RECT 17.935 11.255 18.185 14.785 ;
  LAYER M1 ;
        RECT 18.365 23.015 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.365 21.755 18.615 22.765 ;
  LAYER M1 ;
        RECT 18.365 17.135 18.615 20.665 ;
  LAYER M1 ;
        RECT 18.365 15.875 18.615 16.885 ;
  LAYER M1 ;
        RECT 18.365 11.255 18.615 14.785 ;
  LAYER M1 ;
        RECT 18.365 9.995 18.615 11.005 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 8.905 ;
  LAYER M1 ;
        RECT 18.795 23.015 19.045 26.545 ;
  LAYER M1 ;
        RECT 18.795 17.135 19.045 20.665 ;
  LAYER M1 ;
        RECT 18.795 11.255 19.045 14.785 ;
  LAYER M1 ;
        RECT 19.225 23.015 19.475 26.545 ;
  LAYER M1 ;
        RECT 19.225 21.755 19.475 22.765 ;
  LAYER M1 ;
        RECT 19.225 17.135 19.475 20.665 ;
  LAYER M1 ;
        RECT 19.225 15.875 19.475 16.885 ;
  LAYER M1 ;
        RECT 19.225 11.255 19.475 14.785 ;
  LAYER M1 ;
        RECT 19.225 9.995 19.475 11.005 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 8.905 ;
  LAYER M1 ;
        RECT 19.655 23.015 19.905 26.545 ;
  LAYER M1 ;
        RECT 19.655 17.135 19.905 20.665 ;
  LAYER M1 ;
        RECT 19.655 11.255 19.905 14.785 ;
  LAYER M1 ;
        RECT 20.085 23.015 20.335 26.545 ;
  LAYER M1 ;
        RECT 20.085 21.755 20.335 22.765 ;
  LAYER M1 ;
        RECT 20.085 17.135 20.335 20.665 ;
  LAYER M1 ;
        RECT 20.085 15.875 20.335 16.885 ;
  LAYER M1 ;
        RECT 20.085 11.255 20.335 14.785 ;
  LAYER M1 ;
        RECT 20.085 9.995 20.335 11.005 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 8.905 ;
  LAYER M1 ;
        RECT 20.515 23.015 20.765 26.545 ;
  LAYER M1 ;
        RECT 20.515 17.135 20.765 20.665 ;
  LAYER M1 ;
        RECT 20.515 11.255 20.765 14.785 ;
  LAYER M1 ;
        RECT 20.945 23.015 21.195 26.545 ;
  LAYER M1 ;
        RECT 20.945 21.755 21.195 22.765 ;
  LAYER M1 ;
        RECT 20.945 17.135 21.195 20.665 ;
  LAYER M1 ;
        RECT 20.945 15.875 21.195 16.885 ;
  LAYER M1 ;
        RECT 20.945 11.255 21.195 14.785 ;
  LAYER M1 ;
        RECT 20.945 9.995 21.195 11.005 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 8.905 ;
  LAYER M1 ;
        RECT 21.375 23.015 21.625 26.545 ;
  LAYER M1 ;
        RECT 21.375 17.135 21.625 20.665 ;
  LAYER M1 ;
        RECT 21.375 11.255 21.625 14.785 ;
  LAYER M1 ;
        RECT 21.805 23.015 22.055 26.545 ;
  LAYER M1 ;
        RECT 21.805 21.755 22.055 22.765 ;
  LAYER M1 ;
        RECT 21.805 17.135 22.055 20.665 ;
  LAYER M1 ;
        RECT 21.805 15.875 22.055 16.885 ;
  LAYER M1 ;
        RECT 21.805 11.255 22.055 14.785 ;
  LAYER M1 ;
        RECT 21.805 9.995 22.055 11.005 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 8.905 ;
  LAYER M1 ;
        RECT 22.235 23.015 22.485 26.545 ;
  LAYER M1 ;
        RECT 22.235 17.135 22.485 20.665 ;
  LAYER M1 ;
        RECT 22.235 11.255 22.485 14.785 ;
  LAYER M1 ;
        RECT 22.665 23.015 22.915 26.545 ;
  LAYER M1 ;
        RECT 22.665 21.755 22.915 22.765 ;
  LAYER M1 ;
        RECT 22.665 17.135 22.915 20.665 ;
  LAYER M1 ;
        RECT 22.665 15.875 22.915 16.885 ;
  LAYER M1 ;
        RECT 22.665 11.255 22.915 14.785 ;
  LAYER M1 ;
        RECT 22.665 9.995 22.915 11.005 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 8.905 ;
  LAYER M1 ;
        RECT 23.095 23.015 23.345 26.545 ;
  LAYER M1 ;
        RECT 23.095 17.135 23.345 20.665 ;
  LAYER M1 ;
        RECT 23.095 11.255 23.345 14.785 ;
  LAYER M2 ;
        RECT 17.46 26.32 22.96 26.6 ;
  LAYER M2 ;
        RECT 17.46 22.12 22.96 22.4 ;
  LAYER M2 ;
        RECT 17.03 25.9 23.39 26.18 ;
  LAYER M2 ;
        RECT 17.46 20.44 22.96 20.72 ;
  LAYER M2 ;
        RECT 17.46 16.24 22.96 16.52 ;
  LAYER M2 ;
        RECT 17.03 20.02 23.39 20.3 ;
  LAYER M2 ;
        RECT 17.46 14.56 22.96 14.84 ;
  LAYER M2 ;
        RECT 17.46 10.36 22.96 10.64 ;
  LAYER M2 ;
        RECT 17.03 14.14 23.39 14.42 ;
  LAYER M2 ;
        RECT 17.46 8.26 22.96 8.54 ;
  LAYER M3 ;
        RECT 19.64 14.54 19.92 26.62 ;
  LAYER M3 ;
        RECT 20.07 10.34 20.35 22.42 ;
  LAYER M3 ;
        RECT 20.5 8.24 20.78 26.2 ;
  LAYER M1 ;
        RECT 1.165 27.215 1.415 30.745 ;
  LAYER M1 ;
        RECT 1.165 30.995 1.415 32.005 ;
  LAYER M1 ;
        RECT 1.165 33.095 1.415 34.105 ;
  LAYER M1 ;
        RECT 0.735 27.215 0.985 30.745 ;
  LAYER M1 ;
        RECT 1.595 27.215 1.845 30.745 ;
  LAYER M1 ;
        RECT 2.025 27.215 2.275 30.745 ;
  LAYER M1 ;
        RECT 2.025 30.995 2.275 32.005 ;
  LAYER M1 ;
        RECT 2.025 33.095 2.275 34.105 ;
  LAYER M1 ;
        RECT 2.455 27.215 2.705 30.745 ;
  LAYER M1 ;
        RECT 2.885 27.215 3.135 30.745 ;
  LAYER M1 ;
        RECT 2.885 30.995 3.135 32.005 ;
  LAYER M1 ;
        RECT 2.885 33.095 3.135 34.105 ;
  LAYER M1 ;
        RECT 3.315 27.215 3.565 30.745 ;
  LAYER M1 ;
        RECT 3.745 27.215 3.995 30.745 ;
  LAYER M1 ;
        RECT 3.745 30.995 3.995 32.005 ;
  LAYER M1 ;
        RECT 3.745 33.095 3.995 34.105 ;
  LAYER M1 ;
        RECT 4.175 27.215 4.425 30.745 ;
  LAYER M1 ;
        RECT 4.605 27.215 4.855 30.745 ;
  LAYER M1 ;
        RECT 4.605 30.995 4.855 32.005 ;
  LAYER M1 ;
        RECT 4.605 33.095 4.855 34.105 ;
  LAYER M1 ;
        RECT 5.035 27.215 5.285 30.745 ;
  LAYER M1 ;
        RECT 5.465 27.215 5.715 30.745 ;
  LAYER M1 ;
        RECT 5.465 30.995 5.715 32.005 ;
  LAYER M1 ;
        RECT 5.465 33.095 5.715 34.105 ;
  LAYER M1 ;
        RECT 5.895 27.215 6.145 30.745 ;
  LAYER M1 ;
        RECT 6.325 27.215 6.575 30.745 ;
  LAYER M1 ;
        RECT 6.325 30.995 6.575 32.005 ;
  LAYER M1 ;
        RECT 6.325 33.095 6.575 34.105 ;
  LAYER M1 ;
        RECT 6.755 27.215 7.005 30.745 ;
  LAYER M1 ;
        RECT 7.185 27.215 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 30.995 7.435 32.005 ;
  LAYER M1 ;
        RECT 7.185 33.095 7.435 34.105 ;
  LAYER M1 ;
        RECT 7.615 27.215 7.865 30.745 ;
  LAYER M1 ;
        RECT 8.045 27.215 8.295 30.745 ;
  LAYER M1 ;
        RECT 8.045 30.995 8.295 32.005 ;
  LAYER M1 ;
        RECT 8.045 33.095 8.295 34.105 ;
  LAYER M1 ;
        RECT 8.475 27.215 8.725 30.745 ;
  LAYER M1 ;
        RECT 8.905 27.215 9.155 30.745 ;
  LAYER M1 ;
        RECT 8.905 30.995 9.155 32.005 ;
  LAYER M1 ;
        RECT 8.905 33.095 9.155 34.105 ;
  LAYER M1 ;
        RECT 9.335 27.215 9.585 30.745 ;
  LAYER M1 ;
        RECT 9.765 27.215 10.015 30.745 ;
  LAYER M1 ;
        RECT 9.765 30.995 10.015 32.005 ;
  LAYER M1 ;
        RECT 9.765 33.095 10.015 34.105 ;
  LAYER M1 ;
        RECT 10.195 27.215 10.445 30.745 ;
  LAYER M1 ;
        RECT 10.625 27.215 10.875 30.745 ;
  LAYER M1 ;
        RECT 10.625 30.995 10.875 32.005 ;
  LAYER M1 ;
        RECT 10.625 33.095 10.875 34.105 ;
  LAYER M1 ;
        RECT 11.055 27.215 11.305 30.745 ;
  LAYER M2 ;
        RECT 1.12 31.36 10.92 31.64 ;
  LAYER M2 ;
        RECT 1.12 27.16 10.92 27.44 ;
  LAYER M2 ;
        RECT 1.12 33.46 10.92 33.74 ;
  LAYER M3 ;
        RECT 5.45 27.14 5.73 31.66 ;
  LAYER M2 ;
        RECT 0.69 27.58 11.35 27.86 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M2 ;
        RECT 16.6 0.7 19.52 0.98 ;
  LAYER M2 ;
        RECT 16.6 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 16.6 2.8 19.52 3.08 ;
  LAYER M2 ;
        RECT 16.17 6.58 19.95 6.86 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 4.56 0.7 7.48 0.98 ;
  LAYER M2 ;
        RECT 4.56 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 4.13 6.58 7.91 6.86 ;
  LAYER M1 ;
        RECT 22.665 27.215 22.915 30.745 ;
  LAYER M1 ;
        RECT 22.665 30.995 22.915 32.005 ;
  LAYER M1 ;
        RECT 22.665 33.095 22.915 34.105 ;
  LAYER M1 ;
        RECT 23.095 27.215 23.345 30.745 ;
  LAYER M1 ;
        RECT 22.235 27.215 22.485 30.745 ;
  LAYER M1 ;
        RECT 21.805 27.215 22.055 30.745 ;
  LAYER M1 ;
        RECT 21.805 30.995 22.055 32.005 ;
  LAYER M1 ;
        RECT 21.805 33.095 22.055 34.105 ;
  LAYER M1 ;
        RECT 21.375 27.215 21.625 30.745 ;
  LAYER M1 ;
        RECT 20.945 27.215 21.195 30.745 ;
  LAYER M1 ;
        RECT 20.945 30.995 21.195 32.005 ;
  LAYER M1 ;
        RECT 20.945 33.095 21.195 34.105 ;
  LAYER M1 ;
        RECT 20.515 27.215 20.765 30.745 ;
  LAYER M1 ;
        RECT 20.085 27.215 20.335 30.745 ;
  LAYER M1 ;
        RECT 20.085 30.995 20.335 32.005 ;
  LAYER M1 ;
        RECT 20.085 33.095 20.335 34.105 ;
  LAYER M1 ;
        RECT 19.655 27.215 19.905 30.745 ;
  LAYER M1 ;
        RECT 19.225 27.215 19.475 30.745 ;
  LAYER M1 ;
        RECT 19.225 30.995 19.475 32.005 ;
  LAYER M1 ;
        RECT 19.225 33.095 19.475 34.105 ;
  LAYER M1 ;
        RECT 18.795 27.215 19.045 30.745 ;
  LAYER M1 ;
        RECT 18.365 27.215 18.615 30.745 ;
  LAYER M1 ;
        RECT 18.365 30.995 18.615 32.005 ;
  LAYER M1 ;
        RECT 18.365 33.095 18.615 34.105 ;
  LAYER M1 ;
        RECT 17.935 27.215 18.185 30.745 ;
  LAYER M1 ;
        RECT 17.505 27.215 17.755 30.745 ;
  LAYER M1 ;
        RECT 17.505 30.995 17.755 32.005 ;
  LAYER M1 ;
        RECT 17.505 33.095 17.755 34.105 ;
  LAYER M1 ;
        RECT 17.075 27.215 17.325 30.745 ;
  LAYER M1 ;
        RECT 16.645 27.215 16.895 30.745 ;
  LAYER M1 ;
        RECT 16.645 30.995 16.895 32.005 ;
  LAYER M1 ;
        RECT 16.645 33.095 16.895 34.105 ;
  LAYER M1 ;
        RECT 16.215 27.215 16.465 30.745 ;
  LAYER M1 ;
        RECT 15.785 27.215 16.035 30.745 ;
  LAYER M1 ;
        RECT 15.785 30.995 16.035 32.005 ;
  LAYER M1 ;
        RECT 15.785 33.095 16.035 34.105 ;
  LAYER M1 ;
        RECT 15.355 27.215 15.605 30.745 ;
  LAYER M1 ;
        RECT 14.925 27.215 15.175 30.745 ;
  LAYER M1 ;
        RECT 14.925 30.995 15.175 32.005 ;
  LAYER M1 ;
        RECT 14.925 33.095 15.175 34.105 ;
  LAYER M1 ;
        RECT 14.495 27.215 14.745 30.745 ;
  LAYER M1 ;
        RECT 14.065 27.215 14.315 30.745 ;
  LAYER M1 ;
        RECT 14.065 30.995 14.315 32.005 ;
  LAYER M1 ;
        RECT 14.065 33.095 14.315 34.105 ;
  LAYER M1 ;
        RECT 13.635 27.215 13.885 30.745 ;
  LAYER M1 ;
        RECT 13.205 27.215 13.455 30.745 ;
  LAYER M1 ;
        RECT 13.205 30.995 13.455 32.005 ;
  LAYER M1 ;
        RECT 13.205 33.095 13.455 34.105 ;
  LAYER M1 ;
        RECT 12.775 27.215 13.025 30.745 ;
  LAYER M2 ;
        RECT 13.16 33.46 22.96 33.74 ;
  LAYER M2 ;
        RECT 13.16 27.16 22.96 27.44 ;
  LAYER M2 ;
        RECT 13.16 31.36 22.96 31.64 ;
  LAYER M2 ;
        RECT 12.73 27.58 23.39 27.86 ;
  END 
END CURRENT_MIRROR_OTA
