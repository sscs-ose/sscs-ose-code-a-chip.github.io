MACRO DCL_NMOS_S_54772057_X32_Y3
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_S_54772057_X32_Y3 0 0 ;
  SIZE 29240 BY 19320 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 14480 260 14760 16540 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 14910 680 15190 18640 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 18985 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 18985 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 18985 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 18985 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 18985 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 18985 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 18985 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 18985 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 15625 ;
    LAYER M1 ;
      RECT 8045 15875 8295 16885 ;
    LAYER M1 ;
      RECT 8045 17975 8295 18985 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8475 12095 8725 15625 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 15625 ;
    LAYER M1 ;
      RECT 8905 15875 9155 16885 ;
    LAYER M1 ;
      RECT 8905 17975 9155 18985 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9335 12095 9585 15625 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 9745 ;
    LAYER M1 ;
      RECT 9765 9995 10015 11005 ;
    LAYER M1 ;
      RECT 9765 12095 10015 15625 ;
    LAYER M1 ;
      RECT 9765 15875 10015 16885 ;
    LAYER M1 ;
      RECT 9765 17975 10015 18985 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 6215 10445 9745 ;
    LAYER M1 ;
      RECT 10195 12095 10445 15625 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 9745 ;
    LAYER M1 ;
      RECT 10625 9995 10875 11005 ;
    LAYER M1 ;
      RECT 10625 12095 10875 15625 ;
    LAYER M1 ;
      RECT 10625 15875 10875 16885 ;
    LAYER M1 ;
      RECT 10625 17975 10875 18985 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11055 6215 11305 9745 ;
    LAYER M1 ;
      RECT 11055 12095 11305 15625 ;
    LAYER M1 ;
      RECT 11485 335 11735 3865 ;
    LAYER M1 ;
      RECT 11485 4115 11735 5125 ;
    LAYER M1 ;
      RECT 11485 6215 11735 9745 ;
    LAYER M1 ;
      RECT 11485 9995 11735 11005 ;
    LAYER M1 ;
      RECT 11485 12095 11735 15625 ;
    LAYER M1 ;
      RECT 11485 15875 11735 16885 ;
    LAYER M1 ;
      RECT 11485 17975 11735 18985 ;
    LAYER M1 ;
      RECT 11915 335 12165 3865 ;
    LAYER M1 ;
      RECT 11915 6215 12165 9745 ;
    LAYER M1 ;
      RECT 11915 12095 12165 15625 ;
    LAYER M1 ;
      RECT 12345 335 12595 3865 ;
    LAYER M1 ;
      RECT 12345 4115 12595 5125 ;
    LAYER M1 ;
      RECT 12345 6215 12595 9745 ;
    LAYER M1 ;
      RECT 12345 9995 12595 11005 ;
    LAYER M1 ;
      RECT 12345 12095 12595 15625 ;
    LAYER M1 ;
      RECT 12345 15875 12595 16885 ;
    LAYER M1 ;
      RECT 12345 17975 12595 18985 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M1 ;
      RECT 12775 6215 13025 9745 ;
    LAYER M1 ;
      RECT 12775 12095 13025 15625 ;
    LAYER M1 ;
      RECT 13205 335 13455 3865 ;
    LAYER M1 ;
      RECT 13205 4115 13455 5125 ;
    LAYER M1 ;
      RECT 13205 6215 13455 9745 ;
    LAYER M1 ;
      RECT 13205 9995 13455 11005 ;
    LAYER M1 ;
      RECT 13205 12095 13455 15625 ;
    LAYER M1 ;
      RECT 13205 15875 13455 16885 ;
    LAYER M1 ;
      RECT 13205 17975 13455 18985 ;
    LAYER M1 ;
      RECT 13635 335 13885 3865 ;
    LAYER M1 ;
      RECT 13635 6215 13885 9745 ;
    LAYER M1 ;
      RECT 13635 12095 13885 15625 ;
    LAYER M1 ;
      RECT 14065 335 14315 3865 ;
    LAYER M1 ;
      RECT 14065 4115 14315 5125 ;
    LAYER M1 ;
      RECT 14065 6215 14315 9745 ;
    LAYER M1 ;
      RECT 14065 9995 14315 11005 ;
    LAYER M1 ;
      RECT 14065 12095 14315 15625 ;
    LAYER M1 ;
      RECT 14065 15875 14315 16885 ;
    LAYER M1 ;
      RECT 14065 17975 14315 18985 ;
    LAYER M1 ;
      RECT 14495 335 14745 3865 ;
    LAYER M1 ;
      RECT 14495 6215 14745 9745 ;
    LAYER M1 ;
      RECT 14495 12095 14745 15625 ;
    LAYER M1 ;
      RECT 14925 335 15175 3865 ;
    LAYER M1 ;
      RECT 14925 4115 15175 5125 ;
    LAYER M1 ;
      RECT 14925 6215 15175 9745 ;
    LAYER M1 ;
      RECT 14925 9995 15175 11005 ;
    LAYER M1 ;
      RECT 14925 12095 15175 15625 ;
    LAYER M1 ;
      RECT 14925 15875 15175 16885 ;
    LAYER M1 ;
      RECT 14925 17975 15175 18985 ;
    LAYER M1 ;
      RECT 15355 335 15605 3865 ;
    LAYER M1 ;
      RECT 15355 6215 15605 9745 ;
    LAYER M1 ;
      RECT 15355 12095 15605 15625 ;
    LAYER M1 ;
      RECT 15785 335 16035 3865 ;
    LAYER M1 ;
      RECT 15785 4115 16035 5125 ;
    LAYER M1 ;
      RECT 15785 6215 16035 9745 ;
    LAYER M1 ;
      RECT 15785 9995 16035 11005 ;
    LAYER M1 ;
      RECT 15785 12095 16035 15625 ;
    LAYER M1 ;
      RECT 15785 15875 16035 16885 ;
    LAYER M1 ;
      RECT 15785 17975 16035 18985 ;
    LAYER M1 ;
      RECT 16215 335 16465 3865 ;
    LAYER M1 ;
      RECT 16215 6215 16465 9745 ;
    LAYER M1 ;
      RECT 16215 12095 16465 15625 ;
    LAYER M1 ;
      RECT 16645 335 16895 3865 ;
    LAYER M1 ;
      RECT 16645 4115 16895 5125 ;
    LAYER M1 ;
      RECT 16645 6215 16895 9745 ;
    LAYER M1 ;
      RECT 16645 9995 16895 11005 ;
    LAYER M1 ;
      RECT 16645 12095 16895 15625 ;
    LAYER M1 ;
      RECT 16645 15875 16895 16885 ;
    LAYER M1 ;
      RECT 16645 17975 16895 18985 ;
    LAYER M1 ;
      RECT 17075 335 17325 3865 ;
    LAYER M1 ;
      RECT 17075 6215 17325 9745 ;
    LAYER M1 ;
      RECT 17075 12095 17325 15625 ;
    LAYER M1 ;
      RECT 17505 335 17755 3865 ;
    LAYER M1 ;
      RECT 17505 4115 17755 5125 ;
    LAYER M1 ;
      RECT 17505 6215 17755 9745 ;
    LAYER M1 ;
      RECT 17505 9995 17755 11005 ;
    LAYER M1 ;
      RECT 17505 12095 17755 15625 ;
    LAYER M1 ;
      RECT 17505 15875 17755 16885 ;
    LAYER M1 ;
      RECT 17505 17975 17755 18985 ;
    LAYER M1 ;
      RECT 17935 335 18185 3865 ;
    LAYER M1 ;
      RECT 17935 6215 18185 9745 ;
    LAYER M1 ;
      RECT 17935 12095 18185 15625 ;
    LAYER M1 ;
      RECT 18365 335 18615 3865 ;
    LAYER M1 ;
      RECT 18365 4115 18615 5125 ;
    LAYER M1 ;
      RECT 18365 6215 18615 9745 ;
    LAYER M1 ;
      RECT 18365 9995 18615 11005 ;
    LAYER M1 ;
      RECT 18365 12095 18615 15625 ;
    LAYER M1 ;
      RECT 18365 15875 18615 16885 ;
    LAYER M1 ;
      RECT 18365 17975 18615 18985 ;
    LAYER M1 ;
      RECT 18795 335 19045 3865 ;
    LAYER M1 ;
      RECT 18795 6215 19045 9745 ;
    LAYER M1 ;
      RECT 18795 12095 19045 15625 ;
    LAYER M1 ;
      RECT 19225 335 19475 3865 ;
    LAYER M1 ;
      RECT 19225 4115 19475 5125 ;
    LAYER M1 ;
      RECT 19225 6215 19475 9745 ;
    LAYER M1 ;
      RECT 19225 9995 19475 11005 ;
    LAYER M1 ;
      RECT 19225 12095 19475 15625 ;
    LAYER M1 ;
      RECT 19225 15875 19475 16885 ;
    LAYER M1 ;
      RECT 19225 17975 19475 18985 ;
    LAYER M1 ;
      RECT 19655 335 19905 3865 ;
    LAYER M1 ;
      RECT 19655 6215 19905 9745 ;
    LAYER M1 ;
      RECT 19655 12095 19905 15625 ;
    LAYER M1 ;
      RECT 20085 335 20335 3865 ;
    LAYER M1 ;
      RECT 20085 4115 20335 5125 ;
    LAYER M1 ;
      RECT 20085 6215 20335 9745 ;
    LAYER M1 ;
      RECT 20085 9995 20335 11005 ;
    LAYER M1 ;
      RECT 20085 12095 20335 15625 ;
    LAYER M1 ;
      RECT 20085 15875 20335 16885 ;
    LAYER M1 ;
      RECT 20085 17975 20335 18985 ;
    LAYER M1 ;
      RECT 20515 335 20765 3865 ;
    LAYER M1 ;
      RECT 20515 6215 20765 9745 ;
    LAYER M1 ;
      RECT 20515 12095 20765 15625 ;
    LAYER M1 ;
      RECT 20945 335 21195 3865 ;
    LAYER M1 ;
      RECT 20945 4115 21195 5125 ;
    LAYER M1 ;
      RECT 20945 6215 21195 9745 ;
    LAYER M1 ;
      RECT 20945 9995 21195 11005 ;
    LAYER M1 ;
      RECT 20945 12095 21195 15625 ;
    LAYER M1 ;
      RECT 20945 15875 21195 16885 ;
    LAYER M1 ;
      RECT 20945 17975 21195 18985 ;
    LAYER M1 ;
      RECT 21375 335 21625 3865 ;
    LAYER M1 ;
      RECT 21375 6215 21625 9745 ;
    LAYER M1 ;
      RECT 21375 12095 21625 15625 ;
    LAYER M1 ;
      RECT 21805 335 22055 3865 ;
    LAYER M1 ;
      RECT 21805 4115 22055 5125 ;
    LAYER M1 ;
      RECT 21805 6215 22055 9745 ;
    LAYER M1 ;
      RECT 21805 9995 22055 11005 ;
    LAYER M1 ;
      RECT 21805 12095 22055 15625 ;
    LAYER M1 ;
      RECT 21805 15875 22055 16885 ;
    LAYER M1 ;
      RECT 21805 17975 22055 18985 ;
    LAYER M1 ;
      RECT 22235 335 22485 3865 ;
    LAYER M1 ;
      RECT 22235 6215 22485 9745 ;
    LAYER M1 ;
      RECT 22235 12095 22485 15625 ;
    LAYER M1 ;
      RECT 22665 335 22915 3865 ;
    LAYER M1 ;
      RECT 22665 4115 22915 5125 ;
    LAYER M1 ;
      RECT 22665 6215 22915 9745 ;
    LAYER M1 ;
      RECT 22665 9995 22915 11005 ;
    LAYER M1 ;
      RECT 22665 12095 22915 15625 ;
    LAYER M1 ;
      RECT 22665 15875 22915 16885 ;
    LAYER M1 ;
      RECT 22665 17975 22915 18985 ;
    LAYER M1 ;
      RECT 23095 335 23345 3865 ;
    LAYER M1 ;
      RECT 23095 6215 23345 9745 ;
    LAYER M1 ;
      RECT 23095 12095 23345 15625 ;
    LAYER M1 ;
      RECT 23525 335 23775 3865 ;
    LAYER M1 ;
      RECT 23525 4115 23775 5125 ;
    LAYER M1 ;
      RECT 23525 6215 23775 9745 ;
    LAYER M1 ;
      RECT 23525 9995 23775 11005 ;
    LAYER M1 ;
      RECT 23525 12095 23775 15625 ;
    LAYER M1 ;
      RECT 23525 15875 23775 16885 ;
    LAYER M1 ;
      RECT 23525 17975 23775 18985 ;
    LAYER M1 ;
      RECT 23955 335 24205 3865 ;
    LAYER M1 ;
      RECT 23955 6215 24205 9745 ;
    LAYER M1 ;
      RECT 23955 12095 24205 15625 ;
    LAYER M1 ;
      RECT 24385 335 24635 3865 ;
    LAYER M1 ;
      RECT 24385 4115 24635 5125 ;
    LAYER M1 ;
      RECT 24385 6215 24635 9745 ;
    LAYER M1 ;
      RECT 24385 9995 24635 11005 ;
    LAYER M1 ;
      RECT 24385 12095 24635 15625 ;
    LAYER M1 ;
      RECT 24385 15875 24635 16885 ;
    LAYER M1 ;
      RECT 24385 17975 24635 18985 ;
    LAYER M1 ;
      RECT 24815 335 25065 3865 ;
    LAYER M1 ;
      RECT 24815 6215 25065 9745 ;
    LAYER M1 ;
      RECT 24815 12095 25065 15625 ;
    LAYER M1 ;
      RECT 25245 335 25495 3865 ;
    LAYER M1 ;
      RECT 25245 4115 25495 5125 ;
    LAYER M1 ;
      RECT 25245 6215 25495 9745 ;
    LAYER M1 ;
      RECT 25245 9995 25495 11005 ;
    LAYER M1 ;
      RECT 25245 12095 25495 15625 ;
    LAYER M1 ;
      RECT 25245 15875 25495 16885 ;
    LAYER M1 ;
      RECT 25245 17975 25495 18985 ;
    LAYER M1 ;
      RECT 25675 335 25925 3865 ;
    LAYER M1 ;
      RECT 25675 6215 25925 9745 ;
    LAYER M1 ;
      RECT 25675 12095 25925 15625 ;
    LAYER M1 ;
      RECT 26105 335 26355 3865 ;
    LAYER M1 ;
      RECT 26105 4115 26355 5125 ;
    LAYER M1 ;
      RECT 26105 6215 26355 9745 ;
    LAYER M1 ;
      RECT 26105 9995 26355 11005 ;
    LAYER M1 ;
      RECT 26105 12095 26355 15625 ;
    LAYER M1 ;
      RECT 26105 15875 26355 16885 ;
    LAYER M1 ;
      RECT 26105 17975 26355 18985 ;
    LAYER M1 ;
      RECT 26535 335 26785 3865 ;
    LAYER M1 ;
      RECT 26535 6215 26785 9745 ;
    LAYER M1 ;
      RECT 26535 12095 26785 15625 ;
    LAYER M1 ;
      RECT 26965 335 27215 3865 ;
    LAYER M1 ;
      RECT 26965 4115 27215 5125 ;
    LAYER M1 ;
      RECT 26965 6215 27215 9745 ;
    LAYER M1 ;
      RECT 26965 9995 27215 11005 ;
    LAYER M1 ;
      RECT 26965 12095 27215 15625 ;
    LAYER M1 ;
      RECT 26965 15875 27215 16885 ;
    LAYER M1 ;
      RECT 26965 17975 27215 18985 ;
    LAYER M1 ;
      RECT 27395 335 27645 3865 ;
    LAYER M1 ;
      RECT 27395 6215 27645 9745 ;
    LAYER M1 ;
      RECT 27395 12095 27645 15625 ;
    LAYER M1 ;
      RECT 27825 335 28075 3865 ;
    LAYER M1 ;
      RECT 27825 4115 28075 5125 ;
    LAYER M1 ;
      RECT 27825 6215 28075 9745 ;
    LAYER M1 ;
      RECT 27825 9995 28075 11005 ;
    LAYER M1 ;
      RECT 27825 12095 28075 15625 ;
    LAYER M1 ;
      RECT 27825 15875 28075 16885 ;
    LAYER M1 ;
      RECT 27825 17975 28075 18985 ;
    LAYER M1 ;
      RECT 28255 335 28505 3865 ;
    LAYER M1 ;
      RECT 28255 6215 28505 9745 ;
    LAYER M1 ;
      RECT 28255 12095 28505 15625 ;
    LAYER M2 ;
      RECT 1120 280 28120 560 ;
    LAYER M2 ;
      RECT 1120 4480 28120 4760 ;
    LAYER M2 ;
      RECT 690 700 28550 980 ;
    LAYER M2 ;
      RECT 1120 6160 28120 6440 ;
    LAYER M2 ;
      RECT 1120 10360 28120 10640 ;
    LAYER M2 ;
      RECT 690 6580 28550 6860 ;
    LAYER M2 ;
      RECT 1120 12040 28120 12320 ;
    LAYER M2 ;
      RECT 1120 16240 28120 16520 ;
    LAYER M2 ;
      RECT 1120 18340 28120 18620 ;
    LAYER M2 ;
      RECT 690 12460 28550 12740 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 18395 1375 18565 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 18395 2235 18565 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 18395 3095 18565 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 18395 3955 18565 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 18395 4815 18565 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 18395 5675 18565 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 18395 6535 18565 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 18395 7395 18565 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12095 8255 12265 ;
    LAYER V1 ;
      RECT 8085 16295 8255 16465 ;
    LAYER V1 ;
      RECT 8085 18395 8255 18565 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12095 9115 12265 ;
    LAYER V1 ;
      RECT 8945 16295 9115 16465 ;
    LAYER V1 ;
      RECT 8945 18395 9115 18565 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6215 9975 6385 ;
    LAYER V1 ;
      RECT 9805 10415 9975 10585 ;
    LAYER V1 ;
      RECT 9805 12095 9975 12265 ;
    LAYER V1 ;
      RECT 9805 16295 9975 16465 ;
    LAYER V1 ;
      RECT 9805 18395 9975 18565 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6215 10835 6385 ;
    LAYER V1 ;
      RECT 10665 10415 10835 10585 ;
    LAYER V1 ;
      RECT 10665 12095 10835 12265 ;
    LAYER V1 ;
      RECT 10665 16295 10835 16465 ;
    LAYER V1 ;
      RECT 10665 18395 10835 18565 ;
    LAYER V1 ;
      RECT 11525 335 11695 505 ;
    LAYER V1 ;
      RECT 11525 4535 11695 4705 ;
    LAYER V1 ;
      RECT 11525 6215 11695 6385 ;
    LAYER V1 ;
      RECT 11525 10415 11695 10585 ;
    LAYER V1 ;
      RECT 11525 12095 11695 12265 ;
    LAYER V1 ;
      RECT 11525 16295 11695 16465 ;
    LAYER V1 ;
      RECT 11525 18395 11695 18565 ;
    LAYER V1 ;
      RECT 12385 335 12555 505 ;
    LAYER V1 ;
      RECT 12385 4535 12555 4705 ;
    LAYER V1 ;
      RECT 12385 6215 12555 6385 ;
    LAYER V1 ;
      RECT 12385 10415 12555 10585 ;
    LAYER V1 ;
      RECT 12385 12095 12555 12265 ;
    LAYER V1 ;
      RECT 12385 16295 12555 16465 ;
    LAYER V1 ;
      RECT 12385 18395 12555 18565 ;
    LAYER V1 ;
      RECT 13245 335 13415 505 ;
    LAYER V1 ;
      RECT 13245 4535 13415 4705 ;
    LAYER V1 ;
      RECT 13245 6215 13415 6385 ;
    LAYER V1 ;
      RECT 13245 10415 13415 10585 ;
    LAYER V1 ;
      RECT 13245 12095 13415 12265 ;
    LAYER V1 ;
      RECT 13245 16295 13415 16465 ;
    LAYER V1 ;
      RECT 13245 18395 13415 18565 ;
    LAYER V1 ;
      RECT 14105 335 14275 505 ;
    LAYER V1 ;
      RECT 14105 4535 14275 4705 ;
    LAYER V1 ;
      RECT 14105 6215 14275 6385 ;
    LAYER V1 ;
      RECT 14105 10415 14275 10585 ;
    LAYER V1 ;
      RECT 14105 12095 14275 12265 ;
    LAYER V1 ;
      RECT 14105 16295 14275 16465 ;
    LAYER V1 ;
      RECT 14105 18395 14275 18565 ;
    LAYER V1 ;
      RECT 14965 335 15135 505 ;
    LAYER V1 ;
      RECT 14965 4535 15135 4705 ;
    LAYER V1 ;
      RECT 14965 6215 15135 6385 ;
    LAYER V1 ;
      RECT 14965 10415 15135 10585 ;
    LAYER V1 ;
      RECT 14965 12095 15135 12265 ;
    LAYER V1 ;
      RECT 14965 16295 15135 16465 ;
    LAYER V1 ;
      RECT 14965 18395 15135 18565 ;
    LAYER V1 ;
      RECT 15825 335 15995 505 ;
    LAYER V1 ;
      RECT 15825 4535 15995 4705 ;
    LAYER V1 ;
      RECT 15825 6215 15995 6385 ;
    LAYER V1 ;
      RECT 15825 10415 15995 10585 ;
    LAYER V1 ;
      RECT 15825 12095 15995 12265 ;
    LAYER V1 ;
      RECT 15825 16295 15995 16465 ;
    LAYER V1 ;
      RECT 15825 18395 15995 18565 ;
    LAYER V1 ;
      RECT 16685 335 16855 505 ;
    LAYER V1 ;
      RECT 16685 4535 16855 4705 ;
    LAYER V1 ;
      RECT 16685 6215 16855 6385 ;
    LAYER V1 ;
      RECT 16685 10415 16855 10585 ;
    LAYER V1 ;
      RECT 16685 12095 16855 12265 ;
    LAYER V1 ;
      RECT 16685 16295 16855 16465 ;
    LAYER V1 ;
      RECT 16685 18395 16855 18565 ;
    LAYER V1 ;
      RECT 17545 335 17715 505 ;
    LAYER V1 ;
      RECT 17545 4535 17715 4705 ;
    LAYER V1 ;
      RECT 17545 6215 17715 6385 ;
    LAYER V1 ;
      RECT 17545 10415 17715 10585 ;
    LAYER V1 ;
      RECT 17545 12095 17715 12265 ;
    LAYER V1 ;
      RECT 17545 16295 17715 16465 ;
    LAYER V1 ;
      RECT 17545 18395 17715 18565 ;
    LAYER V1 ;
      RECT 18405 335 18575 505 ;
    LAYER V1 ;
      RECT 18405 4535 18575 4705 ;
    LAYER V1 ;
      RECT 18405 6215 18575 6385 ;
    LAYER V1 ;
      RECT 18405 10415 18575 10585 ;
    LAYER V1 ;
      RECT 18405 12095 18575 12265 ;
    LAYER V1 ;
      RECT 18405 16295 18575 16465 ;
    LAYER V1 ;
      RECT 18405 18395 18575 18565 ;
    LAYER V1 ;
      RECT 19265 335 19435 505 ;
    LAYER V1 ;
      RECT 19265 4535 19435 4705 ;
    LAYER V1 ;
      RECT 19265 6215 19435 6385 ;
    LAYER V1 ;
      RECT 19265 10415 19435 10585 ;
    LAYER V1 ;
      RECT 19265 12095 19435 12265 ;
    LAYER V1 ;
      RECT 19265 16295 19435 16465 ;
    LAYER V1 ;
      RECT 19265 18395 19435 18565 ;
    LAYER V1 ;
      RECT 20125 335 20295 505 ;
    LAYER V1 ;
      RECT 20125 4535 20295 4705 ;
    LAYER V1 ;
      RECT 20125 6215 20295 6385 ;
    LAYER V1 ;
      RECT 20125 10415 20295 10585 ;
    LAYER V1 ;
      RECT 20125 12095 20295 12265 ;
    LAYER V1 ;
      RECT 20125 16295 20295 16465 ;
    LAYER V1 ;
      RECT 20125 18395 20295 18565 ;
    LAYER V1 ;
      RECT 20985 335 21155 505 ;
    LAYER V1 ;
      RECT 20985 4535 21155 4705 ;
    LAYER V1 ;
      RECT 20985 6215 21155 6385 ;
    LAYER V1 ;
      RECT 20985 10415 21155 10585 ;
    LAYER V1 ;
      RECT 20985 12095 21155 12265 ;
    LAYER V1 ;
      RECT 20985 16295 21155 16465 ;
    LAYER V1 ;
      RECT 20985 18395 21155 18565 ;
    LAYER V1 ;
      RECT 21845 335 22015 505 ;
    LAYER V1 ;
      RECT 21845 4535 22015 4705 ;
    LAYER V1 ;
      RECT 21845 6215 22015 6385 ;
    LAYER V1 ;
      RECT 21845 10415 22015 10585 ;
    LAYER V1 ;
      RECT 21845 12095 22015 12265 ;
    LAYER V1 ;
      RECT 21845 16295 22015 16465 ;
    LAYER V1 ;
      RECT 21845 18395 22015 18565 ;
    LAYER V1 ;
      RECT 22705 335 22875 505 ;
    LAYER V1 ;
      RECT 22705 4535 22875 4705 ;
    LAYER V1 ;
      RECT 22705 6215 22875 6385 ;
    LAYER V1 ;
      RECT 22705 10415 22875 10585 ;
    LAYER V1 ;
      RECT 22705 12095 22875 12265 ;
    LAYER V1 ;
      RECT 22705 16295 22875 16465 ;
    LAYER V1 ;
      RECT 22705 18395 22875 18565 ;
    LAYER V1 ;
      RECT 23565 335 23735 505 ;
    LAYER V1 ;
      RECT 23565 4535 23735 4705 ;
    LAYER V1 ;
      RECT 23565 6215 23735 6385 ;
    LAYER V1 ;
      RECT 23565 10415 23735 10585 ;
    LAYER V1 ;
      RECT 23565 12095 23735 12265 ;
    LAYER V1 ;
      RECT 23565 16295 23735 16465 ;
    LAYER V1 ;
      RECT 23565 18395 23735 18565 ;
    LAYER V1 ;
      RECT 24425 335 24595 505 ;
    LAYER V1 ;
      RECT 24425 4535 24595 4705 ;
    LAYER V1 ;
      RECT 24425 6215 24595 6385 ;
    LAYER V1 ;
      RECT 24425 10415 24595 10585 ;
    LAYER V1 ;
      RECT 24425 12095 24595 12265 ;
    LAYER V1 ;
      RECT 24425 16295 24595 16465 ;
    LAYER V1 ;
      RECT 24425 18395 24595 18565 ;
    LAYER V1 ;
      RECT 25285 335 25455 505 ;
    LAYER V1 ;
      RECT 25285 4535 25455 4705 ;
    LAYER V1 ;
      RECT 25285 6215 25455 6385 ;
    LAYER V1 ;
      RECT 25285 10415 25455 10585 ;
    LAYER V1 ;
      RECT 25285 12095 25455 12265 ;
    LAYER V1 ;
      RECT 25285 16295 25455 16465 ;
    LAYER V1 ;
      RECT 25285 18395 25455 18565 ;
    LAYER V1 ;
      RECT 26145 335 26315 505 ;
    LAYER V1 ;
      RECT 26145 4535 26315 4705 ;
    LAYER V1 ;
      RECT 26145 6215 26315 6385 ;
    LAYER V1 ;
      RECT 26145 10415 26315 10585 ;
    LAYER V1 ;
      RECT 26145 12095 26315 12265 ;
    LAYER V1 ;
      RECT 26145 16295 26315 16465 ;
    LAYER V1 ;
      RECT 26145 18395 26315 18565 ;
    LAYER V1 ;
      RECT 27005 335 27175 505 ;
    LAYER V1 ;
      RECT 27005 4535 27175 4705 ;
    LAYER V1 ;
      RECT 27005 6215 27175 6385 ;
    LAYER V1 ;
      RECT 27005 10415 27175 10585 ;
    LAYER V1 ;
      RECT 27005 12095 27175 12265 ;
    LAYER V1 ;
      RECT 27005 16295 27175 16465 ;
    LAYER V1 ;
      RECT 27005 18395 27175 18565 ;
    LAYER V1 ;
      RECT 27865 335 28035 505 ;
    LAYER V1 ;
      RECT 27865 4535 28035 4705 ;
    LAYER V1 ;
      RECT 27865 6215 28035 6385 ;
    LAYER V1 ;
      RECT 27865 10415 28035 10585 ;
    LAYER V1 ;
      RECT 27865 12095 28035 12265 ;
    LAYER V1 ;
      RECT 27865 16295 28035 16465 ;
    LAYER V1 ;
      RECT 27865 18395 28035 18565 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 8515 12515 8685 12685 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 9375 6635 9545 6805 ;
    LAYER V1 ;
      RECT 9375 12515 9545 12685 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 10235 6635 10405 6805 ;
    LAYER V1 ;
      RECT 10235 12515 10405 12685 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11095 6635 11265 6805 ;
    LAYER V1 ;
      RECT 11095 12515 11265 12685 ;
    LAYER V1 ;
      RECT 11955 755 12125 925 ;
    LAYER V1 ;
      RECT 11955 6635 12125 6805 ;
    LAYER V1 ;
      RECT 11955 12515 12125 12685 ;
    LAYER V1 ;
      RECT 12815 755 12985 925 ;
    LAYER V1 ;
      RECT 12815 6635 12985 6805 ;
    LAYER V1 ;
      RECT 12815 12515 12985 12685 ;
    LAYER V1 ;
      RECT 13675 755 13845 925 ;
    LAYER V1 ;
      RECT 13675 6635 13845 6805 ;
    LAYER V1 ;
      RECT 13675 12515 13845 12685 ;
    LAYER V1 ;
      RECT 14535 755 14705 925 ;
    LAYER V1 ;
      RECT 14535 6635 14705 6805 ;
    LAYER V1 ;
      RECT 14535 12515 14705 12685 ;
    LAYER V1 ;
      RECT 15395 755 15565 925 ;
    LAYER V1 ;
      RECT 15395 6635 15565 6805 ;
    LAYER V1 ;
      RECT 15395 12515 15565 12685 ;
    LAYER V1 ;
      RECT 16255 755 16425 925 ;
    LAYER V1 ;
      RECT 16255 6635 16425 6805 ;
    LAYER V1 ;
      RECT 16255 12515 16425 12685 ;
    LAYER V1 ;
      RECT 17115 755 17285 925 ;
    LAYER V1 ;
      RECT 17115 6635 17285 6805 ;
    LAYER V1 ;
      RECT 17115 12515 17285 12685 ;
    LAYER V1 ;
      RECT 17975 755 18145 925 ;
    LAYER V1 ;
      RECT 17975 6635 18145 6805 ;
    LAYER V1 ;
      RECT 17975 12515 18145 12685 ;
    LAYER V1 ;
      RECT 18835 755 19005 925 ;
    LAYER V1 ;
      RECT 18835 6635 19005 6805 ;
    LAYER V1 ;
      RECT 18835 12515 19005 12685 ;
    LAYER V1 ;
      RECT 19695 755 19865 925 ;
    LAYER V1 ;
      RECT 19695 6635 19865 6805 ;
    LAYER V1 ;
      RECT 19695 12515 19865 12685 ;
    LAYER V1 ;
      RECT 20555 755 20725 925 ;
    LAYER V1 ;
      RECT 20555 6635 20725 6805 ;
    LAYER V1 ;
      RECT 20555 12515 20725 12685 ;
    LAYER V1 ;
      RECT 21415 755 21585 925 ;
    LAYER V1 ;
      RECT 21415 6635 21585 6805 ;
    LAYER V1 ;
      RECT 21415 12515 21585 12685 ;
    LAYER V1 ;
      RECT 22275 755 22445 925 ;
    LAYER V1 ;
      RECT 22275 6635 22445 6805 ;
    LAYER V1 ;
      RECT 22275 12515 22445 12685 ;
    LAYER V1 ;
      RECT 23135 755 23305 925 ;
    LAYER V1 ;
      RECT 23135 6635 23305 6805 ;
    LAYER V1 ;
      RECT 23135 12515 23305 12685 ;
    LAYER V1 ;
      RECT 23995 755 24165 925 ;
    LAYER V1 ;
      RECT 23995 6635 24165 6805 ;
    LAYER V1 ;
      RECT 23995 12515 24165 12685 ;
    LAYER V1 ;
      RECT 24855 755 25025 925 ;
    LAYER V1 ;
      RECT 24855 6635 25025 6805 ;
    LAYER V1 ;
      RECT 24855 12515 25025 12685 ;
    LAYER V1 ;
      RECT 25715 755 25885 925 ;
    LAYER V1 ;
      RECT 25715 6635 25885 6805 ;
    LAYER V1 ;
      RECT 25715 12515 25885 12685 ;
    LAYER V1 ;
      RECT 26575 755 26745 925 ;
    LAYER V1 ;
      RECT 26575 6635 26745 6805 ;
    LAYER V1 ;
      RECT 26575 12515 26745 12685 ;
    LAYER V1 ;
      RECT 27435 755 27605 925 ;
    LAYER V1 ;
      RECT 27435 6635 27605 6805 ;
    LAYER V1 ;
      RECT 27435 12515 27605 12685 ;
    LAYER V1 ;
      RECT 28295 755 28465 925 ;
    LAYER V1 ;
      RECT 28295 6635 28465 6805 ;
    LAYER V1 ;
      RECT 28295 12515 28465 12685 ;
    LAYER V2 ;
      RECT 14545 345 14695 495 ;
    LAYER V2 ;
      RECT 14545 4545 14695 4695 ;
    LAYER V2 ;
      RECT 14545 6225 14695 6375 ;
    LAYER V2 ;
      RECT 14545 10425 14695 10575 ;
    LAYER V2 ;
      RECT 14545 12105 14695 12255 ;
    LAYER V2 ;
      RECT 14545 16305 14695 16455 ;
    LAYER V2 ;
      RECT 14975 765 15125 915 ;
    LAYER V2 ;
      RECT 14975 6645 15125 6795 ;
    LAYER V2 ;
      RECT 14975 12525 15125 12675 ;
    LAYER V2 ;
      RECT 14975 18405 15125 18555 ;
  END
END DCL_NMOS_S_54772057_X32_Y3
