MACRO NMOS_S_12565100_X1_Y148
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_12565100_X1_Y148 0 0 ;
  SIZE 2580 BY 871920 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720 260 1000 864940 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 4460 1430 869140 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 871240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 68545 ;
    LAYER M1 ;
      RECT 1165 68795 1415 69805 ;
    LAYER M1 ;
      RECT 1165 70895 1415 74425 ;
    LAYER M1 ;
      RECT 1165 74675 1415 75685 ;
    LAYER M1 ;
      RECT 1165 76775 1415 80305 ;
    LAYER M1 ;
      RECT 1165 80555 1415 81565 ;
    LAYER M1 ;
      RECT 1165 82655 1415 86185 ;
    LAYER M1 ;
      RECT 1165 86435 1415 87445 ;
    LAYER M1 ;
      RECT 1165 88535 1415 92065 ;
    LAYER M1 ;
      RECT 1165 92315 1415 93325 ;
    LAYER M1 ;
      RECT 1165 94415 1415 97945 ;
    LAYER M1 ;
      RECT 1165 98195 1415 99205 ;
    LAYER M1 ;
      RECT 1165 100295 1415 103825 ;
    LAYER M1 ;
      RECT 1165 104075 1415 105085 ;
    LAYER M1 ;
      RECT 1165 106175 1415 109705 ;
    LAYER M1 ;
      RECT 1165 109955 1415 110965 ;
    LAYER M1 ;
      RECT 1165 112055 1415 115585 ;
    LAYER M1 ;
      RECT 1165 115835 1415 116845 ;
    LAYER M1 ;
      RECT 1165 117935 1415 121465 ;
    LAYER M1 ;
      RECT 1165 121715 1415 122725 ;
    LAYER M1 ;
      RECT 1165 123815 1415 127345 ;
    LAYER M1 ;
      RECT 1165 127595 1415 128605 ;
    LAYER M1 ;
      RECT 1165 129695 1415 133225 ;
    LAYER M1 ;
      RECT 1165 133475 1415 134485 ;
    LAYER M1 ;
      RECT 1165 135575 1415 139105 ;
    LAYER M1 ;
      RECT 1165 139355 1415 140365 ;
    LAYER M1 ;
      RECT 1165 141455 1415 144985 ;
    LAYER M1 ;
      RECT 1165 145235 1415 146245 ;
    LAYER M1 ;
      RECT 1165 147335 1415 150865 ;
    LAYER M1 ;
      RECT 1165 151115 1415 152125 ;
    LAYER M1 ;
      RECT 1165 153215 1415 156745 ;
    LAYER M1 ;
      RECT 1165 156995 1415 158005 ;
    LAYER M1 ;
      RECT 1165 159095 1415 162625 ;
    LAYER M1 ;
      RECT 1165 162875 1415 163885 ;
    LAYER M1 ;
      RECT 1165 164975 1415 168505 ;
    LAYER M1 ;
      RECT 1165 168755 1415 169765 ;
    LAYER M1 ;
      RECT 1165 170855 1415 174385 ;
    LAYER M1 ;
      RECT 1165 174635 1415 175645 ;
    LAYER M1 ;
      RECT 1165 176735 1415 180265 ;
    LAYER M1 ;
      RECT 1165 180515 1415 181525 ;
    LAYER M1 ;
      RECT 1165 182615 1415 186145 ;
    LAYER M1 ;
      RECT 1165 186395 1415 187405 ;
    LAYER M1 ;
      RECT 1165 188495 1415 192025 ;
    LAYER M1 ;
      RECT 1165 192275 1415 193285 ;
    LAYER M1 ;
      RECT 1165 194375 1415 197905 ;
    LAYER M1 ;
      RECT 1165 198155 1415 199165 ;
    LAYER M1 ;
      RECT 1165 200255 1415 203785 ;
    LAYER M1 ;
      RECT 1165 204035 1415 205045 ;
    LAYER M1 ;
      RECT 1165 206135 1415 209665 ;
    LAYER M1 ;
      RECT 1165 209915 1415 210925 ;
    LAYER M1 ;
      RECT 1165 212015 1415 215545 ;
    LAYER M1 ;
      RECT 1165 215795 1415 216805 ;
    LAYER M1 ;
      RECT 1165 217895 1415 221425 ;
    LAYER M1 ;
      RECT 1165 221675 1415 222685 ;
    LAYER M1 ;
      RECT 1165 223775 1415 227305 ;
    LAYER M1 ;
      RECT 1165 227555 1415 228565 ;
    LAYER M1 ;
      RECT 1165 229655 1415 233185 ;
    LAYER M1 ;
      RECT 1165 233435 1415 234445 ;
    LAYER M1 ;
      RECT 1165 235535 1415 239065 ;
    LAYER M1 ;
      RECT 1165 239315 1415 240325 ;
    LAYER M1 ;
      RECT 1165 241415 1415 244945 ;
    LAYER M1 ;
      RECT 1165 245195 1415 246205 ;
    LAYER M1 ;
      RECT 1165 247295 1415 250825 ;
    LAYER M1 ;
      RECT 1165 251075 1415 252085 ;
    LAYER M1 ;
      RECT 1165 253175 1415 256705 ;
    LAYER M1 ;
      RECT 1165 256955 1415 257965 ;
    LAYER M1 ;
      RECT 1165 259055 1415 262585 ;
    LAYER M1 ;
      RECT 1165 262835 1415 263845 ;
    LAYER M1 ;
      RECT 1165 264935 1415 268465 ;
    LAYER M1 ;
      RECT 1165 268715 1415 269725 ;
    LAYER M1 ;
      RECT 1165 270815 1415 274345 ;
    LAYER M1 ;
      RECT 1165 274595 1415 275605 ;
    LAYER M1 ;
      RECT 1165 276695 1415 280225 ;
    LAYER M1 ;
      RECT 1165 280475 1415 281485 ;
    LAYER M1 ;
      RECT 1165 282575 1415 286105 ;
    LAYER M1 ;
      RECT 1165 286355 1415 287365 ;
    LAYER M1 ;
      RECT 1165 288455 1415 291985 ;
    LAYER M1 ;
      RECT 1165 292235 1415 293245 ;
    LAYER M1 ;
      RECT 1165 294335 1415 297865 ;
    LAYER M1 ;
      RECT 1165 298115 1415 299125 ;
    LAYER M1 ;
      RECT 1165 300215 1415 303745 ;
    LAYER M1 ;
      RECT 1165 303995 1415 305005 ;
    LAYER M1 ;
      RECT 1165 306095 1415 309625 ;
    LAYER M1 ;
      RECT 1165 309875 1415 310885 ;
    LAYER M1 ;
      RECT 1165 311975 1415 315505 ;
    LAYER M1 ;
      RECT 1165 315755 1415 316765 ;
    LAYER M1 ;
      RECT 1165 317855 1415 321385 ;
    LAYER M1 ;
      RECT 1165 321635 1415 322645 ;
    LAYER M1 ;
      RECT 1165 323735 1415 327265 ;
    LAYER M1 ;
      RECT 1165 327515 1415 328525 ;
    LAYER M1 ;
      RECT 1165 329615 1415 333145 ;
    LAYER M1 ;
      RECT 1165 333395 1415 334405 ;
    LAYER M1 ;
      RECT 1165 335495 1415 339025 ;
    LAYER M1 ;
      RECT 1165 339275 1415 340285 ;
    LAYER M1 ;
      RECT 1165 341375 1415 344905 ;
    LAYER M1 ;
      RECT 1165 345155 1415 346165 ;
    LAYER M1 ;
      RECT 1165 347255 1415 350785 ;
    LAYER M1 ;
      RECT 1165 351035 1415 352045 ;
    LAYER M1 ;
      RECT 1165 353135 1415 356665 ;
    LAYER M1 ;
      RECT 1165 356915 1415 357925 ;
    LAYER M1 ;
      RECT 1165 359015 1415 362545 ;
    LAYER M1 ;
      RECT 1165 362795 1415 363805 ;
    LAYER M1 ;
      RECT 1165 364895 1415 368425 ;
    LAYER M1 ;
      RECT 1165 368675 1415 369685 ;
    LAYER M1 ;
      RECT 1165 370775 1415 374305 ;
    LAYER M1 ;
      RECT 1165 374555 1415 375565 ;
    LAYER M1 ;
      RECT 1165 376655 1415 380185 ;
    LAYER M1 ;
      RECT 1165 380435 1415 381445 ;
    LAYER M1 ;
      RECT 1165 382535 1415 386065 ;
    LAYER M1 ;
      RECT 1165 386315 1415 387325 ;
    LAYER M1 ;
      RECT 1165 388415 1415 391945 ;
    LAYER M1 ;
      RECT 1165 392195 1415 393205 ;
    LAYER M1 ;
      RECT 1165 394295 1415 397825 ;
    LAYER M1 ;
      RECT 1165 398075 1415 399085 ;
    LAYER M1 ;
      RECT 1165 400175 1415 403705 ;
    LAYER M1 ;
      RECT 1165 403955 1415 404965 ;
    LAYER M1 ;
      RECT 1165 406055 1415 409585 ;
    LAYER M1 ;
      RECT 1165 409835 1415 410845 ;
    LAYER M1 ;
      RECT 1165 411935 1415 415465 ;
    LAYER M1 ;
      RECT 1165 415715 1415 416725 ;
    LAYER M1 ;
      RECT 1165 417815 1415 421345 ;
    LAYER M1 ;
      RECT 1165 421595 1415 422605 ;
    LAYER M1 ;
      RECT 1165 423695 1415 427225 ;
    LAYER M1 ;
      RECT 1165 427475 1415 428485 ;
    LAYER M1 ;
      RECT 1165 429575 1415 433105 ;
    LAYER M1 ;
      RECT 1165 433355 1415 434365 ;
    LAYER M1 ;
      RECT 1165 435455 1415 438985 ;
    LAYER M1 ;
      RECT 1165 439235 1415 440245 ;
    LAYER M1 ;
      RECT 1165 441335 1415 444865 ;
    LAYER M1 ;
      RECT 1165 445115 1415 446125 ;
    LAYER M1 ;
      RECT 1165 447215 1415 450745 ;
    LAYER M1 ;
      RECT 1165 450995 1415 452005 ;
    LAYER M1 ;
      RECT 1165 453095 1415 456625 ;
    LAYER M1 ;
      RECT 1165 456875 1415 457885 ;
    LAYER M1 ;
      RECT 1165 458975 1415 462505 ;
    LAYER M1 ;
      RECT 1165 462755 1415 463765 ;
    LAYER M1 ;
      RECT 1165 464855 1415 468385 ;
    LAYER M1 ;
      RECT 1165 468635 1415 469645 ;
    LAYER M1 ;
      RECT 1165 470735 1415 474265 ;
    LAYER M1 ;
      RECT 1165 474515 1415 475525 ;
    LAYER M1 ;
      RECT 1165 476615 1415 480145 ;
    LAYER M1 ;
      RECT 1165 480395 1415 481405 ;
    LAYER M1 ;
      RECT 1165 482495 1415 486025 ;
    LAYER M1 ;
      RECT 1165 486275 1415 487285 ;
    LAYER M1 ;
      RECT 1165 488375 1415 491905 ;
    LAYER M1 ;
      RECT 1165 492155 1415 493165 ;
    LAYER M1 ;
      RECT 1165 494255 1415 497785 ;
    LAYER M1 ;
      RECT 1165 498035 1415 499045 ;
    LAYER M1 ;
      RECT 1165 500135 1415 503665 ;
    LAYER M1 ;
      RECT 1165 503915 1415 504925 ;
    LAYER M1 ;
      RECT 1165 506015 1415 509545 ;
    LAYER M1 ;
      RECT 1165 509795 1415 510805 ;
    LAYER M1 ;
      RECT 1165 511895 1415 515425 ;
    LAYER M1 ;
      RECT 1165 515675 1415 516685 ;
    LAYER M1 ;
      RECT 1165 517775 1415 521305 ;
    LAYER M1 ;
      RECT 1165 521555 1415 522565 ;
    LAYER M1 ;
      RECT 1165 523655 1415 527185 ;
    LAYER M1 ;
      RECT 1165 527435 1415 528445 ;
    LAYER M1 ;
      RECT 1165 529535 1415 533065 ;
    LAYER M1 ;
      RECT 1165 533315 1415 534325 ;
    LAYER M1 ;
      RECT 1165 535415 1415 538945 ;
    LAYER M1 ;
      RECT 1165 539195 1415 540205 ;
    LAYER M1 ;
      RECT 1165 541295 1415 544825 ;
    LAYER M1 ;
      RECT 1165 545075 1415 546085 ;
    LAYER M1 ;
      RECT 1165 547175 1415 550705 ;
    LAYER M1 ;
      RECT 1165 550955 1415 551965 ;
    LAYER M1 ;
      RECT 1165 553055 1415 556585 ;
    LAYER M1 ;
      RECT 1165 556835 1415 557845 ;
    LAYER M1 ;
      RECT 1165 558935 1415 562465 ;
    LAYER M1 ;
      RECT 1165 562715 1415 563725 ;
    LAYER M1 ;
      RECT 1165 564815 1415 568345 ;
    LAYER M1 ;
      RECT 1165 568595 1415 569605 ;
    LAYER M1 ;
      RECT 1165 570695 1415 574225 ;
    LAYER M1 ;
      RECT 1165 574475 1415 575485 ;
    LAYER M1 ;
      RECT 1165 576575 1415 580105 ;
    LAYER M1 ;
      RECT 1165 580355 1415 581365 ;
    LAYER M1 ;
      RECT 1165 582455 1415 585985 ;
    LAYER M1 ;
      RECT 1165 586235 1415 587245 ;
    LAYER M1 ;
      RECT 1165 588335 1415 591865 ;
    LAYER M1 ;
      RECT 1165 592115 1415 593125 ;
    LAYER M1 ;
      RECT 1165 594215 1415 597745 ;
    LAYER M1 ;
      RECT 1165 597995 1415 599005 ;
    LAYER M1 ;
      RECT 1165 600095 1415 603625 ;
    LAYER M1 ;
      RECT 1165 603875 1415 604885 ;
    LAYER M1 ;
      RECT 1165 605975 1415 609505 ;
    LAYER M1 ;
      RECT 1165 609755 1415 610765 ;
    LAYER M1 ;
      RECT 1165 611855 1415 615385 ;
    LAYER M1 ;
      RECT 1165 615635 1415 616645 ;
    LAYER M1 ;
      RECT 1165 617735 1415 621265 ;
    LAYER M1 ;
      RECT 1165 621515 1415 622525 ;
    LAYER M1 ;
      RECT 1165 623615 1415 627145 ;
    LAYER M1 ;
      RECT 1165 627395 1415 628405 ;
    LAYER M1 ;
      RECT 1165 629495 1415 633025 ;
    LAYER M1 ;
      RECT 1165 633275 1415 634285 ;
    LAYER M1 ;
      RECT 1165 635375 1415 638905 ;
    LAYER M1 ;
      RECT 1165 639155 1415 640165 ;
    LAYER M1 ;
      RECT 1165 641255 1415 644785 ;
    LAYER M1 ;
      RECT 1165 645035 1415 646045 ;
    LAYER M1 ;
      RECT 1165 647135 1415 650665 ;
    LAYER M1 ;
      RECT 1165 650915 1415 651925 ;
    LAYER M1 ;
      RECT 1165 653015 1415 656545 ;
    LAYER M1 ;
      RECT 1165 656795 1415 657805 ;
    LAYER M1 ;
      RECT 1165 658895 1415 662425 ;
    LAYER M1 ;
      RECT 1165 662675 1415 663685 ;
    LAYER M1 ;
      RECT 1165 664775 1415 668305 ;
    LAYER M1 ;
      RECT 1165 668555 1415 669565 ;
    LAYER M1 ;
      RECT 1165 670655 1415 674185 ;
    LAYER M1 ;
      RECT 1165 674435 1415 675445 ;
    LAYER M1 ;
      RECT 1165 676535 1415 680065 ;
    LAYER M1 ;
      RECT 1165 680315 1415 681325 ;
    LAYER M1 ;
      RECT 1165 682415 1415 685945 ;
    LAYER M1 ;
      RECT 1165 686195 1415 687205 ;
    LAYER M1 ;
      RECT 1165 688295 1415 691825 ;
    LAYER M1 ;
      RECT 1165 692075 1415 693085 ;
    LAYER M1 ;
      RECT 1165 694175 1415 697705 ;
    LAYER M1 ;
      RECT 1165 697955 1415 698965 ;
    LAYER M1 ;
      RECT 1165 700055 1415 703585 ;
    LAYER M1 ;
      RECT 1165 703835 1415 704845 ;
    LAYER M1 ;
      RECT 1165 705935 1415 709465 ;
    LAYER M1 ;
      RECT 1165 709715 1415 710725 ;
    LAYER M1 ;
      RECT 1165 711815 1415 715345 ;
    LAYER M1 ;
      RECT 1165 715595 1415 716605 ;
    LAYER M1 ;
      RECT 1165 717695 1415 721225 ;
    LAYER M1 ;
      RECT 1165 721475 1415 722485 ;
    LAYER M1 ;
      RECT 1165 723575 1415 727105 ;
    LAYER M1 ;
      RECT 1165 727355 1415 728365 ;
    LAYER M1 ;
      RECT 1165 729455 1415 732985 ;
    LAYER M1 ;
      RECT 1165 733235 1415 734245 ;
    LAYER M1 ;
      RECT 1165 735335 1415 738865 ;
    LAYER M1 ;
      RECT 1165 739115 1415 740125 ;
    LAYER M1 ;
      RECT 1165 741215 1415 744745 ;
    LAYER M1 ;
      RECT 1165 744995 1415 746005 ;
    LAYER M1 ;
      RECT 1165 747095 1415 750625 ;
    LAYER M1 ;
      RECT 1165 750875 1415 751885 ;
    LAYER M1 ;
      RECT 1165 752975 1415 756505 ;
    LAYER M1 ;
      RECT 1165 756755 1415 757765 ;
    LAYER M1 ;
      RECT 1165 758855 1415 762385 ;
    LAYER M1 ;
      RECT 1165 762635 1415 763645 ;
    LAYER M1 ;
      RECT 1165 764735 1415 768265 ;
    LAYER M1 ;
      RECT 1165 768515 1415 769525 ;
    LAYER M1 ;
      RECT 1165 770615 1415 774145 ;
    LAYER M1 ;
      RECT 1165 774395 1415 775405 ;
    LAYER M1 ;
      RECT 1165 776495 1415 780025 ;
    LAYER M1 ;
      RECT 1165 780275 1415 781285 ;
    LAYER M1 ;
      RECT 1165 782375 1415 785905 ;
    LAYER M1 ;
      RECT 1165 786155 1415 787165 ;
    LAYER M1 ;
      RECT 1165 788255 1415 791785 ;
    LAYER M1 ;
      RECT 1165 792035 1415 793045 ;
    LAYER M1 ;
      RECT 1165 794135 1415 797665 ;
    LAYER M1 ;
      RECT 1165 797915 1415 798925 ;
    LAYER M1 ;
      RECT 1165 800015 1415 803545 ;
    LAYER M1 ;
      RECT 1165 803795 1415 804805 ;
    LAYER M1 ;
      RECT 1165 805895 1415 809425 ;
    LAYER M1 ;
      RECT 1165 809675 1415 810685 ;
    LAYER M1 ;
      RECT 1165 811775 1415 815305 ;
    LAYER M1 ;
      RECT 1165 815555 1415 816565 ;
    LAYER M1 ;
      RECT 1165 817655 1415 821185 ;
    LAYER M1 ;
      RECT 1165 821435 1415 822445 ;
    LAYER M1 ;
      RECT 1165 823535 1415 827065 ;
    LAYER M1 ;
      RECT 1165 827315 1415 828325 ;
    LAYER M1 ;
      RECT 1165 829415 1415 832945 ;
    LAYER M1 ;
      RECT 1165 833195 1415 834205 ;
    LAYER M1 ;
      RECT 1165 835295 1415 838825 ;
    LAYER M1 ;
      RECT 1165 839075 1415 840085 ;
    LAYER M1 ;
      RECT 1165 841175 1415 844705 ;
    LAYER M1 ;
      RECT 1165 844955 1415 845965 ;
    LAYER M1 ;
      RECT 1165 847055 1415 850585 ;
    LAYER M1 ;
      RECT 1165 850835 1415 851845 ;
    LAYER M1 ;
      RECT 1165 852935 1415 856465 ;
    LAYER M1 ;
      RECT 1165 856715 1415 857725 ;
    LAYER M1 ;
      RECT 1165 858815 1415 862345 ;
    LAYER M1 ;
      RECT 1165 862595 1415 863605 ;
    LAYER M1 ;
      RECT 1165 864695 1415 868225 ;
    LAYER M1 ;
      RECT 1165 868475 1415 869485 ;
    LAYER M1 ;
      RECT 1165 870575 1415 871585 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 735 65015 985 68545 ;
    LAYER M1 ;
      RECT 735 70895 985 74425 ;
    LAYER M1 ;
      RECT 735 76775 985 80305 ;
    LAYER M1 ;
      RECT 735 82655 985 86185 ;
    LAYER M1 ;
      RECT 735 88535 985 92065 ;
    LAYER M1 ;
      RECT 735 94415 985 97945 ;
    LAYER M1 ;
      RECT 735 100295 985 103825 ;
    LAYER M1 ;
      RECT 735 106175 985 109705 ;
    LAYER M1 ;
      RECT 735 112055 985 115585 ;
    LAYER M1 ;
      RECT 735 117935 985 121465 ;
    LAYER M1 ;
      RECT 735 123815 985 127345 ;
    LAYER M1 ;
      RECT 735 129695 985 133225 ;
    LAYER M1 ;
      RECT 735 135575 985 139105 ;
    LAYER M1 ;
      RECT 735 141455 985 144985 ;
    LAYER M1 ;
      RECT 735 147335 985 150865 ;
    LAYER M1 ;
      RECT 735 153215 985 156745 ;
    LAYER M1 ;
      RECT 735 159095 985 162625 ;
    LAYER M1 ;
      RECT 735 164975 985 168505 ;
    LAYER M1 ;
      RECT 735 170855 985 174385 ;
    LAYER M1 ;
      RECT 735 176735 985 180265 ;
    LAYER M1 ;
      RECT 735 182615 985 186145 ;
    LAYER M1 ;
      RECT 735 188495 985 192025 ;
    LAYER M1 ;
      RECT 735 194375 985 197905 ;
    LAYER M1 ;
      RECT 735 200255 985 203785 ;
    LAYER M1 ;
      RECT 735 206135 985 209665 ;
    LAYER M1 ;
      RECT 735 212015 985 215545 ;
    LAYER M1 ;
      RECT 735 217895 985 221425 ;
    LAYER M1 ;
      RECT 735 223775 985 227305 ;
    LAYER M1 ;
      RECT 735 229655 985 233185 ;
    LAYER M1 ;
      RECT 735 235535 985 239065 ;
    LAYER M1 ;
      RECT 735 241415 985 244945 ;
    LAYER M1 ;
      RECT 735 247295 985 250825 ;
    LAYER M1 ;
      RECT 735 253175 985 256705 ;
    LAYER M1 ;
      RECT 735 259055 985 262585 ;
    LAYER M1 ;
      RECT 735 264935 985 268465 ;
    LAYER M1 ;
      RECT 735 270815 985 274345 ;
    LAYER M1 ;
      RECT 735 276695 985 280225 ;
    LAYER M1 ;
      RECT 735 282575 985 286105 ;
    LAYER M1 ;
      RECT 735 288455 985 291985 ;
    LAYER M1 ;
      RECT 735 294335 985 297865 ;
    LAYER M1 ;
      RECT 735 300215 985 303745 ;
    LAYER M1 ;
      RECT 735 306095 985 309625 ;
    LAYER M1 ;
      RECT 735 311975 985 315505 ;
    LAYER M1 ;
      RECT 735 317855 985 321385 ;
    LAYER M1 ;
      RECT 735 323735 985 327265 ;
    LAYER M1 ;
      RECT 735 329615 985 333145 ;
    LAYER M1 ;
      RECT 735 335495 985 339025 ;
    LAYER M1 ;
      RECT 735 341375 985 344905 ;
    LAYER M1 ;
      RECT 735 347255 985 350785 ;
    LAYER M1 ;
      RECT 735 353135 985 356665 ;
    LAYER M1 ;
      RECT 735 359015 985 362545 ;
    LAYER M1 ;
      RECT 735 364895 985 368425 ;
    LAYER M1 ;
      RECT 735 370775 985 374305 ;
    LAYER M1 ;
      RECT 735 376655 985 380185 ;
    LAYER M1 ;
      RECT 735 382535 985 386065 ;
    LAYER M1 ;
      RECT 735 388415 985 391945 ;
    LAYER M1 ;
      RECT 735 394295 985 397825 ;
    LAYER M1 ;
      RECT 735 400175 985 403705 ;
    LAYER M1 ;
      RECT 735 406055 985 409585 ;
    LAYER M1 ;
      RECT 735 411935 985 415465 ;
    LAYER M1 ;
      RECT 735 417815 985 421345 ;
    LAYER M1 ;
      RECT 735 423695 985 427225 ;
    LAYER M1 ;
      RECT 735 429575 985 433105 ;
    LAYER M1 ;
      RECT 735 435455 985 438985 ;
    LAYER M1 ;
      RECT 735 441335 985 444865 ;
    LAYER M1 ;
      RECT 735 447215 985 450745 ;
    LAYER M1 ;
      RECT 735 453095 985 456625 ;
    LAYER M1 ;
      RECT 735 458975 985 462505 ;
    LAYER M1 ;
      RECT 735 464855 985 468385 ;
    LAYER M1 ;
      RECT 735 470735 985 474265 ;
    LAYER M1 ;
      RECT 735 476615 985 480145 ;
    LAYER M1 ;
      RECT 735 482495 985 486025 ;
    LAYER M1 ;
      RECT 735 488375 985 491905 ;
    LAYER M1 ;
      RECT 735 494255 985 497785 ;
    LAYER M1 ;
      RECT 735 500135 985 503665 ;
    LAYER M1 ;
      RECT 735 506015 985 509545 ;
    LAYER M1 ;
      RECT 735 511895 985 515425 ;
    LAYER M1 ;
      RECT 735 517775 985 521305 ;
    LAYER M1 ;
      RECT 735 523655 985 527185 ;
    LAYER M1 ;
      RECT 735 529535 985 533065 ;
    LAYER M1 ;
      RECT 735 535415 985 538945 ;
    LAYER M1 ;
      RECT 735 541295 985 544825 ;
    LAYER M1 ;
      RECT 735 547175 985 550705 ;
    LAYER M1 ;
      RECT 735 553055 985 556585 ;
    LAYER M1 ;
      RECT 735 558935 985 562465 ;
    LAYER M1 ;
      RECT 735 564815 985 568345 ;
    LAYER M1 ;
      RECT 735 570695 985 574225 ;
    LAYER M1 ;
      RECT 735 576575 985 580105 ;
    LAYER M1 ;
      RECT 735 582455 985 585985 ;
    LAYER M1 ;
      RECT 735 588335 985 591865 ;
    LAYER M1 ;
      RECT 735 594215 985 597745 ;
    LAYER M1 ;
      RECT 735 600095 985 603625 ;
    LAYER M1 ;
      RECT 735 605975 985 609505 ;
    LAYER M1 ;
      RECT 735 611855 985 615385 ;
    LAYER M1 ;
      RECT 735 617735 985 621265 ;
    LAYER M1 ;
      RECT 735 623615 985 627145 ;
    LAYER M1 ;
      RECT 735 629495 985 633025 ;
    LAYER M1 ;
      RECT 735 635375 985 638905 ;
    LAYER M1 ;
      RECT 735 641255 985 644785 ;
    LAYER M1 ;
      RECT 735 647135 985 650665 ;
    LAYER M1 ;
      RECT 735 653015 985 656545 ;
    LAYER M1 ;
      RECT 735 658895 985 662425 ;
    LAYER M1 ;
      RECT 735 664775 985 668305 ;
    LAYER M1 ;
      RECT 735 670655 985 674185 ;
    LAYER M1 ;
      RECT 735 676535 985 680065 ;
    LAYER M1 ;
      RECT 735 682415 985 685945 ;
    LAYER M1 ;
      RECT 735 688295 985 691825 ;
    LAYER M1 ;
      RECT 735 694175 985 697705 ;
    LAYER M1 ;
      RECT 735 700055 985 703585 ;
    LAYER M1 ;
      RECT 735 705935 985 709465 ;
    LAYER M1 ;
      RECT 735 711815 985 715345 ;
    LAYER M1 ;
      RECT 735 717695 985 721225 ;
    LAYER M1 ;
      RECT 735 723575 985 727105 ;
    LAYER M1 ;
      RECT 735 729455 985 732985 ;
    LAYER M1 ;
      RECT 735 735335 985 738865 ;
    LAYER M1 ;
      RECT 735 741215 985 744745 ;
    LAYER M1 ;
      RECT 735 747095 985 750625 ;
    LAYER M1 ;
      RECT 735 752975 985 756505 ;
    LAYER M1 ;
      RECT 735 758855 985 762385 ;
    LAYER M1 ;
      RECT 735 764735 985 768265 ;
    LAYER M1 ;
      RECT 735 770615 985 774145 ;
    LAYER M1 ;
      RECT 735 776495 985 780025 ;
    LAYER M1 ;
      RECT 735 782375 985 785905 ;
    LAYER M1 ;
      RECT 735 788255 985 791785 ;
    LAYER M1 ;
      RECT 735 794135 985 797665 ;
    LAYER M1 ;
      RECT 735 800015 985 803545 ;
    LAYER M1 ;
      RECT 735 805895 985 809425 ;
    LAYER M1 ;
      RECT 735 811775 985 815305 ;
    LAYER M1 ;
      RECT 735 817655 985 821185 ;
    LAYER M1 ;
      RECT 735 823535 985 827065 ;
    LAYER M1 ;
      RECT 735 829415 985 832945 ;
    LAYER M1 ;
      RECT 735 835295 985 838825 ;
    LAYER M1 ;
      RECT 735 841175 985 844705 ;
    LAYER M1 ;
      RECT 735 847055 985 850585 ;
    LAYER M1 ;
      RECT 735 852935 985 856465 ;
    LAYER M1 ;
      RECT 735 858815 985 862345 ;
    LAYER M1 ;
      RECT 735 864695 985 868225 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 1595 65015 1845 68545 ;
    LAYER M1 ;
      RECT 1595 70895 1845 74425 ;
    LAYER M1 ;
      RECT 1595 76775 1845 80305 ;
    LAYER M1 ;
      RECT 1595 82655 1845 86185 ;
    LAYER M1 ;
      RECT 1595 88535 1845 92065 ;
    LAYER M1 ;
      RECT 1595 94415 1845 97945 ;
    LAYER M1 ;
      RECT 1595 100295 1845 103825 ;
    LAYER M1 ;
      RECT 1595 106175 1845 109705 ;
    LAYER M1 ;
      RECT 1595 112055 1845 115585 ;
    LAYER M1 ;
      RECT 1595 117935 1845 121465 ;
    LAYER M1 ;
      RECT 1595 123815 1845 127345 ;
    LAYER M1 ;
      RECT 1595 129695 1845 133225 ;
    LAYER M1 ;
      RECT 1595 135575 1845 139105 ;
    LAYER M1 ;
      RECT 1595 141455 1845 144985 ;
    LAYER M1 ;
      RECT 1595 147335 1845 150865 ;
    LAYER M1 ;
      RECT 1595 153215 1845 156745 ;
    LAYER M1 ;
      RECT 1595 159095 1845 162625 ;
    LAYER M1 ;
      RECT 1595 164975 1845 168505 ;
    LAYER M1 ;
      RECT 1595 170855 1845 174385 ;
    LAYER M1 ;
      RECT 1595 176735 1845 180265 ;
    LAYER M1 ;
      RECT 1595 182615 1845 186145 ;
    LAYER M1 ;
      RECT 1595 188495 1845 192025 ;
    LAYER M1 ;
      RECT 1595 194375 1845 197905 ;
    LAYER M1 ;
      RECT 1595 200255 1845 203785 ;
    LAYER M1 ;
      RECT 1595 206135 1845 209665 ;
    LAYER M1 ;
      RECT 1595 212015 1845 215545 ;
    LAYER M1 ;
      RECT 1595 217895 1845 221425 ;
    LAYER M1 ;
      RECT 1595 223775 1845 227305 ;
    LAYER M1 ;
      RECT 1595 229655 1845 233185 ;
    LAYER M1 ;
      RECT 1595 235535 1845 239065 ;
    LAYER M1 ;
      RECT 1595 241415 1845 244945 ;
    LAYER M1 ;
      RECT 1595 247295 1845 250825 ;
    LAYER M1 ;
      RECT 1595 253175 1845 256705 ;
    LAYER M1 ;
      RECT 1595 259055 1845 262585 ;
    LAYER M1 ;
      RECT 1595 264935 1845 268465 ;
    LAYER M1 ;
      RECT 1595 270815 1845 274345 ;
    LAYER M1 ;
      RECT 1595 276695 1845 280225 ;
    LAYER M1 ;
      RECT 1595 282575 1845 286105 ;
    LAYER M1 ;
      RECT 1595 288455 1845 291985 ;
    LAYER M1 ;
      RECT 1595 294335 1845 297865 ;
    LAYER M1 ;
      RECT 1595 300215 1845 303745 ;
    LAYER M1 ;
      RECT 1595 306095 1845 309625 ;
    LAYER M1 ;
      RECT 1595 311975 1845 315505 ;
    LAYER M1 ;
      RECT 1595 317855 1845 321385 ;
    LAYER M1 ;
      RECT 1595 323735 1845 327265 ;
    LAYER M1 ;
      RECT 1595 329615 1845 333145 ;
    LAYER M1 ;
      RECT 1595 335495 1845 339025 ;
    LAYER M1 ;
      RECT 1595 341375 1845 344905 ;
    LAYER M1 ;
      RECT 1595 347255 1845 350785 ;
    LAYER M1 ;
      RECT 1595 353135 1845 356665 ;
    LAYER M1 ;
      RECT 1595 359015 1845 362545 ;
    LAYER M1 ;
      RECT 1595 364895 1845 368425 ;
    LAYER M1 ;
      RECT 1595 370775 1845 374305 ;
    LAYER M1 ;
      RECT 1595 376655 1845 380185 ;
    LAYER M1 ;
      RECT 1595 382535 1845 386065 ;
    LAYER M1 ;
      RECT 1595 388415 1845 391945 ;
    LAYER M1 ;
      RECT 1595 394295 1845 397825 ;
    LAYER M1 ;
      RECT 1595 400175 1845 403705 ;
    LAYER M1 ;
      RECT 1595 406055 1845 409585 ;
    LAYER M1 ;
      RECT 1595 411935 1845 415465 ;
    LAYER M1 ;
      RECT 1595 417815 1845 421345 ;
    LAYER M1 ;
      RECT 1595 423695 1845 427225 ;
    LAYER M1 ;
      RECT 1595 429575 1845 433105 ;
    LAYER M1 ;
      RECT 1595 435455 1845 438985 ;
    LAYER M1 ;
      RECT 1595 441335 1845 444865 ;
    LAYER M1 ;
      RECT 1595 447215 1845 450745 ;
    LAYER M1 ;
      RECT 1595 453095 1845 456625 ;
    LAYER M1 ;
      RECT 1595 458975 1845 462505 ;
    LAYER M1 ;
      RECT 1595 464855 1845 468385 ;
    LAYER M1 ;
      RECT 1595 470735 1845 474265 ;
    LAYER M1 ;
      RECT 1595 476615 1845 480145 ;
    LAYER M1 ;
      RECT 1595 482495 1845 486025 ;
    LAYER M1 ;
      RECT 1595 488375 1845 491905 ;
    LAYER M1 ;
      RECT 1595 494255 1845 497785 ;
    LAYER M1 ;
      RECT 1595 500135 1845 503665 ;
    LAYER M1 ;
      RECT 1595 506015 1845 509545 ;
    LAYER M1 ;
      RECT 1595 511895 1845 515425 ;
    LAYER M1 ;
      RECT 1595 517775 1845 521305 ;
    LAYER M1 ;
      RECT 1595 523655 1845 527185 ;
    LAYER M1 ;
      RECT 1595 529535 1845 533065 ;
    LAYER M1 ;
      RECT 1595 535415 1845 538945 ;
    LAYER M1 ;
      RECT 1595 541295 1845 544825 ;
    LAYER M1 ;
      RECT 1595 547175 1845 550705 ;
    LAYER M1 ;
      RECT 1595 553055 1845 556585 ;
    LAYER M1 ;
      RECT 1595 558935 1845 562465 ;
    LAYER M1 ;
      RECT 1595 564815 1845 568345 ;
    LAYER M1 ;
      RECT 1595 570695 1845 574225 ;
    LAYER M1 ;
      RECT 1595 576575 1845 580105 ;
    LAYER M1 ;
      RECT 1595 582455 1845 585985 ;
    LAYER M1 ;
      RECT 1595 588335 1845 591865 ;
    LAYER M1 ;
      RECT 1595 594215 1845 597745 ;
    LAYER M1 ;
      RECT 1595 600095 1845 603625 ;
    LAYER M1 ;
      RECT 1595 605975 1845 609505 ;
    LAYER M1 ;
      RECT 1595 611855 1845 615385 ;
    LAYER M1 ;
      RECT 1595 617735 1845 621265 ;
    LAYER M1 ;
      RECT 1595 623615 1845 627145 ;
    LAYER M1 ;
      RECT 1595 629495 1845 633025 ;
    LAYER M1 ;
      RECT 1595 635375 1845 638905 ;
    LAYER M1 ;
      RECT 1595 641255 1845 644785 ;
    LAYER M1 ;
      RECT 1595 647135 1845 650665 ;
    LAYER M1 ;
      RECT 1595 653015 1845 656545 ;
    LAYER M1 ;
      RECT 1595 658895 1845 662425 ;
    LAYER M1 ;
      RECT 1595 664775 1845 668305 ;
    LAYER M1 ;
      RECT 1595 670655 1845 674185 ;
    LAYER M1 ;
      RECT 1595 676535 1845 680065 ;
    LAYER M1 ;
      RECT 1595 682415 1845 685945 ;
    LAYER M1 ;
      RECT 1595 688295 1845 691825 ;
    LAYER M1 ;
      RECT 1595 694175 1845 697705 ;
    LAYER M1 ;
      RECT 1595 700055 1845 703585 ;
    LAYER M1 ;
      RECT 1595 705935 1845 709465 ;
    LAYER M1 ;
      RECT 1595 711815 1845 715345 ;
    LAYER M1 ;
      RECT 1595 717695 1845 721225 ;
    LAYER M1 ;
      RECT 1595 723575 1845 727105 ;
    LAYER M1 ;
      RECT 1595 729455 1845 732985 ;
    LAYER M1 ;
      RECT 1595 735335 1845 738865 ;
    LAYER M1 ;
      RECT 1595 741215 1845 744745 ;
    LAYER M1 ;
      RECT 1595 747095 1845 750625 ;
    LAYER M1 ;
      RECT 1595 752975 1845 756505 ;
    LAYER M1 ;
      RECT 1595 758855 1845 762385 ;
    LAYER M1 ;
      RECT 1595 764735 1845 768265 ;
    LAYER M1 ;
      RECT 1595 770615 1845 774145 ;
    LAYER M1 ;
      RECT 1595 776495 1845 780025 ;
    LAYER M1 ;
      RECT 1595 782375 1845 785905 ;
    LAYER M1 ;
      RECT 1595 788255 1845 791785 ;
    LAYER M1 ;
      RECT 1595 794135 1845 797665 ;
    LAYER M1 ;
      RECT 1595 800015 1845 803545 ;
    LAYER M1 ;
      RECT 1595 805895 1845 809425 ;
    LAYER M1 ;
      RECT 1595 811775 1845 815305 ;
    LAYER M1 ;
      RECT 1595 817655 1845 821185 ;
    LAYER M1 ;
      RECT 1595 823535 1845 827065 ;
    LAYER M1 ;
      RECT 1595 829415 1845 832945 ;
    LAYER M1 ;
      RECT 1595 835295 1845 838825 ;
    LAYER M1 ;
      RECT 1595 841175 1845 844705 ;
    LAYER M1 ;
      RECT 1595 847055 1845 850585 ;
    LAYER M1 ;
      RECT 1595 852935 1845 856465 ;
    LAYER M1 ;
      RECT 1595 858815 1845 862345 ;
    LAYER M1 ;
      RECT 1595 864695 1845 868225 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 260 4480 1460 4760 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER M2 ;
      RECT 260 6160 1460 6440 ;
    LAYER M2 ;
      RECT 260 10360 1460 10640 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 260 12040 1460 12320 ;
    LAYER M2 ;
      RECT 260 16240 1460 16520 ;
    LAYER M2 ;
      RECT 690 12460 1890 12740 ;
    LAYER M2 ;
      RECT 260 17920 1460 18200 ;
    LAYER M2 ;
      RECT 260 22120 1460 22400 ;
    LAYER M2 ;
      RECT 690 18340 1890 18620 ;
    LAYER M2 ;
      RECT 260 23800 1460 24080 ;
    LAYER M2 ;
      RECT 260 28000 1460 28280 ;
    LAYER M2 ;
      RECT 690 24220 1890 24500 ;
    LAYER M2 ;
      RECT 260 29680 1460 29960 ;
    LAYER M2 ;
      RECT 260 33880 1460 34160 ;
    LAYER M2 ;
      RECT 690 30100 1890 30380 ;
    LAYER M2 ;
      RECT 260 35560 1460 35840 ;
    LAYER M2 ;
      RECT 260 39760 1460 40040 ;
    LAYER M2 ;
      RECT 690 35980 1890 36260 ;
    LAYER M2 ;
      RECT 260 41440 1460 41720 ;
    LAYER M2 ;
      RECT 260 45640 1460 45920 ;
    LAYER M2 ;
      RECT 690 41860 1890 42140 ;
    LAYER M2 ;
      RECT 260 47320 1460 47600 ;
    LAYER M2 ;
      RECT 260 51520 1460 51800 ;
    LAYER M2 ;
      RECT 690 47740 1890 48020 ;
    LAYER M2 ;
      RECT 260 53200 1460 53480 ;
    LAYER M2 ;
      RECT 260 57400 1460 57680 ;
    LAYER M2 ;
      RECT 690 53620 1890 53900 ;
    LAYER M2 ;
      RECT 260 59080 1460 59360 ;
    LAYER M2 ;
      RECT 260 63280 1460 63560 ;
    LAYER M2 ;
      RECT 690 59500 1890 59780 ;
    LAYER M2 ;
      RECT 260 64960 1460 65240 ;
    LAYER M2 ;
      RECT 260 69160 1460 69440 ;
    LAYER M2 ;
      RECT 690 65380 1890 65660 ;
    LAYER M2 ;
      RECT 260 70840 1460 71120 ;
    LAYER M2 ;
      RECT 260 75040 1460 75320 ;
    LAYER M2 ;
      RECT 690 71260 1890 71540 ;
    LAYER M2 ;
      RECT 260 76720 1460 77000 ;
    LAYER M2 ;
      RECT 260 80920 1460 81200 ;
    LAYER M2 ;
      RECT 690 77140 1890 77420 ;
    LAYER M2 ;
      RECT 260 82600 1460 82880 ;
    LAYER M2 ;
      RECT 260 86800 1460 87080 ;
    LAYER M2 ;
      RECT 690 83020 1890 83300 ;
    LAYER M2 ;
      RECT 260 88480 1460 88760 ;
    LAYER M2 ;
      RECT 260 92680 1460 92960 ;
    LAYER M2 ;
      RECT 690 88900 1890 89180 ;
    LAYER M2 ;
      RECT 260 94360 1460 94640 ;
    LAYER M2 ;
      RECT 260 98560 1460 98840 ;
    LAYER M2 ;
      RECT 690 94780 1890 95060 ;
    LAYER M2 ;
      RECT 260 100240 1460 100520 ;
    LAYER M2 ;
      RECT 260 104440 1460 104720 ;
    LAYER M2 ;
      RECT 690 100660 1890 100940 ;
    LAYER M2 ;
      RECT 260 106120 1460 106400 ;
    LAYER M2 ;
      RECT 260 110320 1460 110600 ;
    LAYER M2 ;
      RECT 690 106540 1890 106820 ;
    LAYER M2 ;
      RECT 260 112000 1460 112280 ;
    LAYER M2 ;
      RECT 260 116200 1460 116480 ;
    LAYER M2 ;
      RECT 690 112420 1890 112700 ;
    LAYER M2 ;
      RECT 260 117880 1460 118160 ;
    LAYER M2 ;
      RECT 260 122080 1460 122360 ;
    LAYER M2 ;
      RECT 690 118300 1890 118580 ;
    LAYER M2 ;
      RECT 260 123760 1460 124040 ;
    LAYER M2 ;
      RECT 260 127960 1460 128240 ;
    LAYER M2 ;
      RECT 690 124180 1890 124460 ;
    LAYER M2 ;
      RECT 260 129640 1460 129920 ;
    LAYER M2 ;
      RECT 260 133840 1460 134120 ;
    LAYER M2 ;
      RECT 690 130060 1890 130340 ;
    LAYER M2 ;
      RECT 260 135520 1460 135800 ;
    LAYER M2 ;
      RECT 260 139720 1460 140000 ;
    LAYER M2 ;
      RECT 690 135940 1890 136220 ;
    LAYER M2 ;
      RECT 260 141400 1460 141680 ;
    LAYER M2 ;
      RECT 260 145600 1460 145880 ;
    LAYER M2 ;
      RECT 690 141820 1890 142100 ;
    LAYER M2 ;
      RECT 260 147280 1460 147560 ;
    LAYER M2 ;
      RECT 260 151480 1460 151760 ;
    LAYER M2 ;
      RECT 690 147700 1890 147980 ;
    LAYER M2 ;
      RECT 260 153160 1460 153440 ;
    LAYER M2 ;
      RECT 260 157360 1460 157640 ;
    LAYER M2 ;
      RECT 690 153580 1890 153860 ;
    LAYER M2 ;
      RECT 260 159040 1460 159320 ;
    LAYER M2 ;
      RECT 260 163240 1460 163520 ;
    LAYER M2 ;
      RECT 690 159460 1890 159740 ;
    LAYER M2 ;
      RECT 260 164920 1460 165200 ;
    LAYER M2 ;
      RECT 260 169120 1460 169400 ;
    LAYER M2 ;
      RECT 690 165340 1890 165620 ;
    LAYER M2 ;
      RECT 260 170800 1460 171080 ;
    LAYER M2 ;
      RECT 260 175000 1460 175280 ;
    LAYER M2 ;
      RECT 690 171220 1890 171500 ;
    LAYER M2 ;
      RECT 260 176680 1460 176960 ;
    LAYER M2 ;
      RECT 260 180880 1460 181160 ;
    LAYER M2 ;
      RECT 690 177100 1890 177380 ;
    LAYER M2 ;
      RECT 260 182560 1460 182840 ;
    LAYER M2 ;
      RECT 260 186760 1460 187040 ;
    LAYER M2 ;
      RECT 690 182980 1890 183260 ;
    LAYER M2 ;
      RECT 260 188440 1460 188720 ;
    LAYER M2 ;
      RECT 260 192640 1460 192920 ;
    LAYER M2 ;
      RECT 690 188860 1890 189140 ;
    LAYER M2 ;
      RECT 260 194320 1460 194600 ;
    LAYER M2 ;
      RECT 260 198520 1460 198800 ;
    LAYER M2 ;
      RECT 690 194740 1890 195020 ;
    LAYER M2 ;
      RECT 260 200200 1460 200480 ;
    LAYER M2 ;
      RECT 260 204400 1460 204680 ;
    LAYER M2 ;
      RECT 690 200620 1890 200900 ;
    LAYER M2 ;
      RECT 260 206080 1460 206360 ;
    LAYER M2 ;
      RECT 260 210280 1460 210560 ;
    LAYER M2 ;
      RECT 690 206500 1890 206780 ;
    LAYER M2 ;
      RECT 260 211960 1460 212240 ;
    LAYER M2 ;
      RECT 260 216160 1460 216440 ;
    LAYER M2 ;
      RECT 690 212380 1890 212660 ;
    LAYER M2 ;
      RECT 260 217840 1460 218120 ;
    LAYER M2 ;
      RECT 260 222040 1460 222320 ;
    LAYER M2 ;
      RECT 690 218260 1890 218540 ;
    LAYER M2 ;
      RECT 260 223720 1460 224000 ;
    LAYER M2 ;
      RECT 260 227920 1460 228200 ;
    LAYER M2 ;
      RECT 690 224140 1890 224420 ;
    LAYER M2 ;
      RECT 260 229600 1460 229880 ;
    LAYER M2 ;
      RECT 260 233800 1460 234080 ;
    LAYER M2 ;
      RECT 690 230020 1890 230300 ;
    LAYER M2 ;
      RECT 260 235480 1460 235760 ;
    LAYER M2 ;
      RECT 260 239680 1460 239960 ;
    LAYER M2 ;
      RECT 690 235900 1890 236180 ;
    LAYER M2 ;
      RECT 260 241360 1460 241640 ;
    LAYER M2 ;
      RECT 260 245560 1460 245840 ;
    LAYER M2 ;
      RECT 690 241780 1890 242060 ;
    LAYER M2 ;
      RECT 260 247240 1460 247520 ;
    LAYER M2 ;
      RECT 260 251440 1460 251720 ;
    LAYER M2 ;
      RECT 690 247660 1890 247940 ;
    LAYER M2 ;
      RECT 260 253120 1460 253400 ;
    LAYER M2 ;
      RECT 260 257320 1460 257600 ;
    LAYER M2 ;
      RECT 690 253540 1890 253820 ;
    LAYER M2 ;
      RECT 260 259000 1460 259280 ;
    LAYER M2 ;
      RECT 260 263200 1460 263480 ;
    LAYER M2 ;
      RECT 690 259420 1890 259700 ;
    LAYER M2 ;
      RECT 260 264880 1460 265160 ;
    LAYER M2 ;
      RECT 260 269080 1460 269360 ;
    LAYER M2 ;
      RECT 690 265300 1890 265580 ;
    LAYER M2 ;
      RECT 260 270760 1460 271040 ;
    LAYER M2 ;
      RECT 260 274960 1460 275240 ;
    LAYER M2 ;
      RECT 690 271180 1890 271460 ;
    LAYER M2 ;
      RECT 260 276640 1460 276920 ;
    LAYER M2 ;
      RECT 260 280840 1460 281120 ;
    LAYER M2 ;
      RECT 690 277060 1890 277340 ;
    LAYER M2 ;
      RECT 260 282520 1460 282800 ;
    LAYER M2 ;
      RECT 260 286720 1460 287000 ;
    LAYER M2 ;
      RECT 690 282940 1890 283220 ;
    LAYER M2 ;
      RECT 260 288400 1460 288680 ;
    LAYER M2 ;
      RECT 260 292600 1460 292880 ;
    LAYER M2 ;
      RECT 690 288820 1890 289100 ;
    LAYER M2 ;
      RECT 260 294280 1460 294560 ;
    LAYER M2 ;
      RECT 260 298480 1460 298760 ;
    LAYER M2 ;
      RECT 690 294700 1890 294980 ;
    LAYER M2 ;
      RECT 260 300160 1460 300440 ;
    LAYER M2 ;
      RECT 260 304360 1460 304640 ;
    LAYER M2 ;
      RECT 690 300580 1890 300860 ;
    LAYER M2 ;
      RECT 260 306040 1460 306320 ;
    LAYER M2 ;
      RECT 260 310240 1460 310520 ;
    LAYER M2 ;
      RECT 690 306460 1890 306740 ;
    LAYER M2 ;
      RECT 260 311920 1460 312200 ;
    LAYER M2 ;
      RECT 260 316120 1460 316400 ;
    LAYER M2 ;
      RECT 690 312340 1890 312620 ;
    LAYER M2 ;
      RECT 260 317800 1460 318080 ;
    LAYER M2 ;
      RECT 260 322000 1460 322280 ;
    LAYER M2 ;
      RECT 690 318220 1890 318500 ;
    LAYER M2 ;
      RECT 260 323680 1460 323960 ;
    LAYER M2 ;
      RECT 260 327880 1460 328160 ;
    LAYER M2 ;
      RECT 690 324100 1890 324380 ;
    LAYER M2 ;
      RECT 260 329560 1460 329840 ;
    LAYER M2 ;
      RECT 260 333760 1460 334040 ;
    LAYER M2 ;
      RECT 690 329980 1890 330260 ;
    LAYER M2 ;
      RECT 260 335440 1460 335720 ;
    LAYER M2 ;
      RECT 260 339640 1460 339920 ;
    LAYER M2 ;
      RECT 690 335860 1890 336140 ;
    LAYER M2 ;
      RECT 260 341320 1460 341600 ;
    LAYER M2 ;
      RECT 260 345520 1460 345800 ;
    LAYER M2 ;
      RECT 690 341740 1890 342020 ;
    LAYER M2 ;
      RECT 260 347200 1460 347480 ;
    LAYER M2 ;
      RECT 260 351400 1460 351680 ;
    LAYER M2 ;
      RECT 690 347620 1890 347900 ;
    LAYER M2 ;
      RECT 260 353080 1460 353360 ;
    LAYER M2 ;
      RECT 260 357280 1460 357560 ;
    LAYER M2 ;
      RECT 690 353500 1890 353780 ;
    LAYER M2 ;
      RECT 260 358960 1460 359240 ;
    LAYER M2 ;
      RECT 260 363160 1460 363440 ;
    LAYER M2 ;
      RECT 690 359380 1890 359660 ;
    LAYER M2 ;
      RECT 260 364840 1460 365120 ;
    LAYER M2 ;
      RECT 260 369040 1460 369320 ;
    LAYER M2 ;
      RECT 690 365260 1890 365540 ;
    LAYER M2 ;
      RECT 260 370720 1460 371000 ;
    LAYER M2 ;
      RECT 260 374920 1460 375200 ;
    LAYER M2 ;
      RECT 690 371140 1890 371420 ;
    LAYER M2 ;
      RECT 260 376600 1460 376880 ;
    LAYER M2 ;
      RECT 260 380800 1460 381080 ;
    LAYER M2 ;
      RECT 690 377020 1890 377300 ;
    LAYER M2 ;
      RECT 260 382480 1460 382760 ;
    LAYER M2 ;
      RECT 260 386680 1460 386960 ;
    LAYER M2 ;
      RECT 690 382900 1890 383180 ;
    LAYER M2 ;
      RECT 260 388360 1460 388640 ;
    LAYER M2 ;
      RECT 260 392560 1460 392840 ;
    LAYER M2 ;
      RECT 690 388780 1890 389060 ;
    LAYER M2 ;
      RECT 260 394240 1460 394520 ;
    LAYER M2 ;
      RECT 260 398440 1460 398720 ;
    LAYER M2 ;
      RECT 690 394660 1890 394940 ;
    LAYER M2 ;
      RECT 260 400120 1460 400400 ;
    LAYER M2 ;
      RECT 260 404320 1460 404600 ;
    LAYER M2 ;
      RECT 690 400540 1890 400820 ;
    LAYER M2 ;
      RECT 260 406000 1460 406280 ;
    LAYER M2 ;
      RECT 260 410200 1460 410480 ;
    LAYER M2 ;
      RECT 690 406420 1890 406700 ;
    LAYER M2 ;
      RECT 260 411880 1460 412160 ;
    LAYER M2 ;
      RECT 260 416080 1460 416360 ;
    LAYER M2 ;
      RECT 690 412300 1890 412580 ;
    LAYER M2 ;
      RECT 260 417760 1460 418040 ;
    LAYER M2 ;
      RECT 260 421960 1460 422240 ;
    LAYER M2 ;
      RECT 690 418180 1890 418460 ;
    LAYER M2 ;
      RECT 260 423640 1460 423920 ;
    LAYER M2 ;
      RECT 260 427840 1460 428120 ;
    LAYER M2 ;
      RECT 690 424060 1890 424340 ;
    LAYER M2 ;
      RECT 260 429520 1460 429800 ;
    LAYER M2 ;
      RECT 260 433720 1460 434000 ;
    LAYER M2 ;
      RECT 690 429940 1890 430220 ;
    LAYER M2 ;
      RECT 260 435400 1460 435680 ;
    LAYER M2 ;
      RECT 260 439600 1460 439880 ;
    LAYER M2 ;
      RECT 690 435820 1890 436100 ;
    LAYER M2 ;
      RECT 260 441280 1460 441560 ;
    LAYER M2 ;
      RECT 260 445480 1460 445760 ;
    LAYER M2 ;
      RECT 690 441700 1890 441980 ;
    LAYER M2 ;
      RECT 260 447160 1460 447440 ;
    LAYER M2 ;
      RECT 260 451360 1460 451640 ;
    LAYER M2 ;
      RECT 690 447580 1890 447860 ;
    LAYER M2 ;
      RECT 260 453040 1460 453320 ;
    LAYER M2 ;
      RECT 260 457240 1460 457520 ;
    LAYER M2 ;
      RECT 690 453460 1890 453740 ;
    LAYER M2 ;
      RECT 260 458920 1460 459200 ;
    LAYER M2 ;
      RECT 260 463120 1460 463400 ;
    LAYER M2 ;
      RECT 690 459340 1890 459620 ;
    LAYER M2 ;
      RECT 260 464800 1460 465080 ;
    LAYER M2 ;
      RECT 260 469000 1460 469280 ;
    LAYER M2 ;
      RECT 690 465220 1890 465500 ;
    LAYER M2 ;
      RECT 260 470680 1460 470960 ;
    LAYER M2 ;
      RECT 260 474880 1460 475160 ;
    LAYER M2 ;
      RECT 690 471100 1890 471380 ;
    LAYER M2 ;
      RECT 260 476560 1460 476840 ;
    LAYER M2 ;
      RECT 260 480760 1460 481040 ;
    LAYER M2 ;
      RECT 690 476980 1890 477260 ;
    LAYER M2 ;
      RECT 260 482440 1460 482720 ;
    LAYER M2 ;
      RECT 260 486640 1460 486920 ;
    LAYER M2 ;
      RECT 690 482860 1890 483140 ;
    LAYER M2 ;
      RECT 260 488320 1460 488600 ;
    LAYER M2 ;
      RECT 260 492520 1460 492800 ;
    LAYER M2 ;
      RECT 690 488740 1890 489020 ;
    LAYER M2 ;
      RECT 260 494200 1460 494480 ;
    LAYER M2 ;
      RECT 260 498400 1460 498680 ;
    LAYER M2 ;
      RECT 690 494620 1890 494900 ;
    LAYER M2 ;
      RECT 260 500080 1460 500360 ;
    LAYER M2 ;
      RECT 260 504280 1460 504560 ;
    LAYER M2 ;
      RECT 690 500500 1890 500780 ;
    LAYER M2 ;
      RECT 260 505960 1460 506240 ;
    LAYER M2 ;
      RECT 260 510160 1460 510440 ;
    LAYER M2 ;
      RECT 690 506380 1890 506660 ;
    LAYER M2 ;
      RECT 260 511840 1460 512120 ;
    LAYER M2 ;
      RECT 260 516040 1460 516320 ;
    LAYER M2 ;
      RECT 690 512260 1890 512540 ;
    LAYER M2 ;
      RECT 260 517720 1460 518000 ;
    LAYER M2 ;
      RECT 260 521920 1460 522200 ;
    LAYER M2 ;
      RECT 690 518140 1890 518420 ;
    LAYER M2 ;
      RECT 260 523600 1460 523880 ;
    LAYER M2 ;
      RECT 260 527800 1460 528080 ;
    LAYER M2 ;
      RECT 690 524020 1890 524300 ;
    LAYER M2 ;
      RECT 260 529480 1460 529760 ;
    LAYER M2 ;
      RECT 260 533680 1460 533960 ;
    LAYER M2 ;
      RECT 690 529900 1890 530180 ;
    LAYER M2 ;
      RECT 260 535360 1460 535640 ;
    LAYER M2 ;
      RECT 260 539560 1460 539840 ;
    LAYER M2 ;
      RECT 690 535780 1890 536060 ;
    LAYER M2 ;
      RECT 260 541240 1460 541520 ;
    LAYER M2 ;
      RECT 260 545440 1460 545720 ;
    LAYER M2 ;
      RECT 690 541660 1890 541940 ;
    LAYER M2 ;
      RECT 260 547120 1460 547400 ;
    LAYER M2 ;
      RECT 260 551320 1460 551600 ;
    LAYER M2 ;
      RECT 690 547540 1890 547820 ;
    LAYER M2 ;
      RECT 260 553000 1460 553280 ;
    LAYER M2 ;
      RECT 260 557200 1460 557480 ;
    LAYER M2 ;
      RECT 690 553420 1890 553700 ;
    LAYER M2 ;
      RECT 260 558880 1460 559160 ;
    LAYER M2 ;
      RECT 260 563080 1460 563360 ;
    LAYER M2 ;
      RECT 690 559300 1890 559580 ;
    LAYER M2 ;
      RECT 260 564760 1460 565040 ;
    LAYER M2 ;
      RECT 260 568960 1460 569240 ;
    LAYER M2 ;
      RECT 690 565180 1890 565460 ;
    LAYER M2 ;
      RECT 260 570640 1460 570920 ;
    LAYER M2 ;
      RECT 260 574840 1460 575120 ;
    LAYER M2 ;
      RECT 690 571060 1890 571340 ;
    LAYER M2 ;
      RECT 260 576520 1460 576800 ;
    LAYER M2 ;
      RECT 260 580720 1460 581000 ;
    LAYER M2 ;
      RECT 690 576940 1890 577220 ;
    LAYER M2 ;
      RECT 260 582400 1460 582680 ;
    LAYER M2 ;
      RECT 260 586600 1460 586880 ;
    LAYER M2 ;
      RECT 690 582820 1890 583100 ;
    LAYER M2 ;
      RECT 260 588280 1460 588560 ;
    LAYER M2 ;
      RECT 260 592480 1460 592760 ;
    LAYER M2 ;
      RECT 690 588700 1890 588980 ;
    LAYER M2 ;
      RECT 260 594160 1460 594440 ;
    LAYER M2 ;
      RECT 260 598360 1460 598640 ;
    LAYER M2 ;
      RECT 690 594580 1890 594860 ;
    LAYER M2 ;
      RECT 260 600040 1460 600320 ;
    LAYER M2 ;
      RECT 260 604240 1460 604520 ;
    LAYER M2 ;
      RECT 690 600460 1890 600740 ;
    LAYER M2 ;
      RECT 260 605920 1460 606200 ;
    LAYER M2 ;
      RECT 260 610120 1460 610400 ;
    LAYER M2 ;
      RECT 690 606340 1890 606620 ;
    LAYER M2 ;
      RECT 260 611800 1460 612080 ;
    LAYER M2 ;
      RECT 260 616000 1460 616280 ;
    LAYER M2 ;
      RECT 690 612220 1890 612500 ;
    LAYER M2 ;
      RECT 260 617680 1460 617960 ;
    LAYER M2 ;
      RECT 260 621880 1460 622160 ;
    LAYER M2 ;
      RECT 690 618100 1890 618380 ;
    LAYER M2 ;
      RECT 260 623560 1460 623840 ;
    LAYER M2 ;
      RECT 260 627760 1460 628040 ;
    LAYER M2 ;
      RECT 690 623980 1890 624260 ;
    LAYER M2 ;
      RECT 260 629440 1460 629720 ;
    LAYER M2 ;
      RECT 260 633640 1460 633920 ;
    LAYER M2 ;
      RECT 690 629860 1890 630140 ;
    LAYER M2 ;
      RECT 260 635320 1460 635600 ;
    LAYER M2 ;
      RECT 260 639520 1460 639800 ;
    LAYER M2 ;
      RECT 690 635740 1890 636020 ;
    LAYER M2 ;
      RECT 260 641200 1460 641480 ;
    LAYER M2 ;
      RECT 260 645400 1460 645680 ;
    LAYER M2 ;
      RECT 690 641620 1890 641900 ;
    LAYER M2 ;
      RECT 260 647080 1460 647360 ;
    LAYER M2 ;
      RECT 260 651280 1460 651560 ;
    LAYER M2 ;
      RECT 690 647500 1890 647780 ;
    LAYER M2 ;
      RECT 260 652960 1460 653240 ;
    LAYER M2 ;
      RECT 260 657160 1460 657440 ;
    LAYER M2 ;
      RECT 690 653380 1890 653660 ;
    LAYER M2 ;
      RECT 260 658840 1460 659120 ;
    LAYER M2 ;
      RECT 260 663040 1460 663320 ;
    LAYER M2 ;
      RECT 690 659260 1890 659540 ;
    LAYER M2 ;
      RECT 260 664720 1460 665000 ;
    LAYER M2 ;
      RECT 260 668920 1460 669200 ;
    LAYER M2 ;
      RECT 690 665140 1890 665420 ;
    LAYER M2 ;
      RECT 260 670600 1460 670880 ;
    LAYER M2 ;
      RECT 260 674800 1460 675080 ;
    LAYER M2 ;
      RECT 690 671020 1890 671300 ;
    LAYER M2 ;
      RECT 260 676480 1460 676760 ;
    LAYER M2 ;
      RECT 260 680680 1460 680960 ;
    LAYER M2 ;
      RECT 690 676900 1890 677180 ;
    LAYER M2 ;
      RECT 260 682360 1460 682640 ;
    LAYER M2 ;
      RECT 260 686560 1460 686840 ;
    LAYER M2 ;
      RECT 690 682780 1890 683060 ;
    LAYER M2 ;
      RECT 260 688240 1460 688520 ;
    LAYER M2 ;
      RECT 260 692440 1460 692720 ;
    LAYER M2 ;
      RECT 690 688660 1890 688940 ;
    LAYER M2 ;
      RECT 260 694120 1460 694400 ;
    LAYER M2 ;
      RECT 260 698320 1460 698600 ;
    LAYER M2 ;
      RECT 690 694540 1890 694820 ;
    LAYER M2 ;
      RECT 260 700000 1460 700280 ;
    LAYER M2 ;
      RECT 260 704200 1460 704480 ;
    LAYER M2 ;
      RECT 690 700420 1890 700700 ;
    LAYER M2 ;
      RECT 260 705880 1460 706160 ;
    LAYER M2 ;
      RECT 260 710080 1460 710360 ;
    LAYER M2 ;
      RECT 690 706300 1890 706580 ;
    LAYER M2 ;
      RECT 260 711760 1460 712040 ;
    LAYER M2 ;
      RECT 260 715960 1460 716240 ;
    LAYER M2 ;
      RECT 690 712180 1890 712460 ;
    LAYER M2 ;
      RECT 260 717640 1460 717920 ;
    LAYER M2 ;
      RECT 260 721840 1460 722120 ;
    LAYER M2 ;
      RECT 690 718060 1890 718340 ;
    LAYER M2 ;
      RECT 260 723520 1460 723800 ;
    LAYER M2 ;
      RECT 260 727720 1460 728000 ;
    LAYER M2 ;
      RECT 690 723940 1890 724220 ;
    LAYER M2 ;
      RECT 260 729400 1460 729680 ;
    LAYER M2 ;
      RECT 260 733600 1460 733880 ;
    LAYER M2 ;
      RECT 690 729820 1890 730100 ;
    LAYER M2 ;
      RECT 260 735280 1460 735560 ;
    LAYER M2 ;
      RECT 260 739480 1460 739760 ;
    LAYER M2 ;
      RECT 690 735700 1890 735980 ;
    LAYER M2 ;
      RECT 260 741160 1460 741440 ;
    LAYER M2 ;
      RECT 260 745360 1460 745640 ;
    LAYER M2 ;
      RECT 690 741580 1890 741860 ;
    LAYER M2 ;
      RECT 260 747040 1460 747320 ;
    LAYER M2 ;
      RECT 260 751240 1460 751520 ;
    LAYER M2 ;
      RECT 690 747460 1890 747740 ;
    LAYER M2 ;
      RECT 260 752920 1460 753200 ;
    LAYER M2 ;
      RECT 260 757120 1460 757400 ;
    LAYER M2 ;
      RECT 690 753340 1890 753620 ;
    LAYER M2 ;
      RECT 260 758800 1460 759080 ;
    LAYER M2 ;
      RECT 260 763000 1460 763280 ;
    LAYER M2 ;
      RECT 690 759220 1890 759500 ;
    LAYER M2 ;
      RECT 260 764680 1460 764960 ;
    LAYER M2 ;
      RECT 260 768880 1460 769160 ;
    LAYER M2 ;
      RECT 690 765100 1890 765380 ;
    LAYER M2 ;
      RECT 260 770560 1460 770840 ;
    LAYER M2 ;
      RECT 260 774760 1460 775040 ;
    LAYER M2 ;
      RECT 690 770980 1890 771260 ;
    LAYER M2 ;
      RECT 260 776440 1460 776720 ;
    LAYER M2 ;
      RECT 260 780640 1460 780920 ;
    LAYER M2 ;
      RECT 690 776860 1890 777140 ;
    LAYER M2 ;
      RECT 260 782320 1460 782600 ;
    LAYER M2 ;
      RECT 260 786520 1460 786800 ;
    LAYER M2 ;
      RECT 690 782740 1890 783020 ;
    LAYER M2 ;
      RECT 260 788200 1460 788480 ;
    LAYER M2 ;
      RECT 260 792400 1460 792680 ;
    LAYER M2 ;
      RECT 690 788620 1890 788900 ;
    LAYER M2 ;
      RECT 260 794080 1460 794360 ;
    LAYER M2 ;
      RECT 260 798280 1460 798560 ;
    LAYER M2 ;
      RECT 690 794500 1890 794780 ;
    LAYER M2 ;
      RECT 260 799960 1460 800240 ;
    LAYER M2 ;
      RECT 260 804160 1460 804440 ;
    LAYER M2 ;
      RECT 690 800380 1890 800660 ;
    LAYER M2 ;
      RECT 260 805840 1460 806120 ;
    LAYER M2 ;
      RECT 260 810040 1460 810320 ;
    LAYER M2 ;
      RECT 690 806260 1890 806540 ;
    LAYER M2 ;
      RECT 260 811720 1460 812000 ;
    LAYER M2 ;
      RECT 260 815920 1460 816200 ;
    LAYER M2 ;
      RECT 690 812140 1890 812420 ;
    LAYER M2 ;
      RECT 260 817600 1460 817880 ;
    LAYER M2 ;
      RECT 260 821800 1460 822080 ;
    LAYER M2 ;
      RECT 690 818020 1890 818300 ;
    LAYER M2 ;
      RECT 260 823480 1460 823760 ;
    LAYER M2 ;
      RECT 260 827680 1460 827960 ;
    LAYER M2 ;
      RECT 690 823900 1890 824180 ;
    LAYER M2 ;
      RECT 260 829360 1460 829640 ;
    LAYER M2 ;
      RECT 260 833560 1460 833840 ;
    LAYER M2 ;
      RECT 690 829780 1890 830060 ;
    LAYER M2 ;
      RECT 260 835240 1460 835520 ;
    LAYER M2 ;
      RECT 260 839440 1460 839720 ;
    LAYER M2 ;
      RECT 690 835660 1890 835940 ;
    LAYER M2 ;
      RECT 260 841120 1460 841400 ;
    LAYER M2 ;
      RECT 260 845320 1460 845600 ;
    LAYER M2 ;
      RECT 690 841540 1890 841820 ;
    LAYER M2 ;
      RECT 260 847000 1460 847280 ;
    LAYER M2 ;
      RECT 260 851200 1460 851480 ;
    LAYER M2 ;
      RECT 690 847420 1890 847700 ;
    LAYER M2 ;
      RECT 260 852880 1460 853160 ;
    LAYER M2 ;
      RECT 260 857080 1460 857360 ;
    LAYER M2 ;
      RECT 690 853300 1890 853580 ;
    LAYER M2 ;
      RECT 260 858760 1460 859040 ;
    LAYER M2 ;
      RECT 260 862960 1460 863240 ;
    LAYER M2 ;
      RECT 690 859180 1890 859460 ;
    LAYER M2 ;
      RECT 260 864640 1460 864920 ;
    LAYER M2 ;
      RECT 260 868840 1460 869120 ;
    LAYER M2 ;
      RECT 690 870940 1890 871220 ;
    LAYER M2 ;
      RECT 690 865060 1890 865340 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53255 1375 53425 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65015 1375 65185 ;
    LAYER V1 ;
      RECT 1205 69215 1375 69385 ;
    LAYER V1 ;
      RECT 1205 70895 1375 71065 ;
    LAYER V1 ;
      RECT 1205 75095 1375 75265 ;
    LAYER V1 ;
      RECT 1205 76775 1375 76945 ;
    LAYER V1 ;
      RECT 1205 80975 1375 81145 ;
    LAYER V1 ;
      RECT 1205 82655 1375 82825 ;
    LAYER V1 ;
      RECT 1205 86855 1375 87025 ;
    LAYER V1 ;
      RECT 1205 88535 1375 88705 ;
    LAYER V1 ;
      RECT 1205 92735 1375 92905 ;
    LAYER V1 ;
      RECT 1205 94415 1375 94585 ;
    LAYER V1 ;
      RECT 1205 98615 1375 98785 ;
    LAYER V1 ;
      RECT 1205 100295 1375 100465 ;
    LAYER V1 ;
      RECT 1205 104495 1375 104665 ;
    LAYER V1 ;
      RECT 1205 106175 1375 106345 ;
    LAYER V1 ;
      RECT 1205 110375 1375 110545 ;
    LAYER V1 ;
      RECT 1205 112055 1375 112225 ;
    LAYER V1 ;
      RECT 1205 116255 1375 116425 ;
    LAYER V1 ;
      RECT 1205 117935 1375 118105 ;
    LAYER V1 ;
      RECT 1205 122135 1375 122305 ;
    LAYER V1 ;
      RECT 1205 123815 1375 123985 ;
    LAYER V1 ;
      RECT 1205 128015 1375 128185 ;
    LAYER V1 ;
      RECT 1205 129695 1375 129865 ;
    LAYER V1 ;
      RECT 1205 133895 1375 134065 ;
    LAYER V1 ;
      RECT 1205 135575 1375 135745 ;
    LAYER V1 ;
      RECT 1205 139775 1375 139945 ;
    LAYER V1 ;
      RECT 1205 141455 1375 141625 ;
    LAYER V1 ;
      RECT 1205 145655 1375 145825 ;
    LAYER V1 ;
      RECT 1205 147335 1375 147505 ;
    LAYER V1 ;
      RECT 1205 151535 1375 151705 ;
    LAYER V1 ;
      RECT 1205 153215 1375 153385 ;
    LAYER V1 ;
      RECT 1205 157415 1375 157585 ;
    LAYER V1 ;
      RECT 1205 159095 1375 159265 ;
    LAYER V1 ;
      RECT 1205 163295 1375 163465 ;
    LAYER V1 ;
      RECT 1205 164975 1375 165145 ;
    LAYER V1 ;
      RECT 1205 169175 1375 169345 ;
    LAYER V1 ;
      RECT 1205 170855 1375 171025 ;
    LAYER V1 ;
      RECT 1205 175055 1375 175225 ;
    LAYER V1 ;
      RECT 1205 176735 1375 176905 ;
    LAYER V1 ;
      RECT 1205 180935 1375 181105 ;
    LAYER V1 ;
      RECT 1205 182615 1375 182785 ;
    LAYER V1 ;
      RECT 1205 186815 1375 186985 ;
    LAYER V1 ;
      RECT 1205 188495 1375 188665 ;
    LAYER V1 ;
      RECT 1205 192695 1375 192865 ;
    LAYER V1 ;
      RECT 1205 194375 1375 194545 ;
    LAYER V1 ;
      RECT 1205 198575 1375 198745 ;
    LAYER V1 ;
      RECT 1205 200255 1375 200425 ;
    LAYER V1 ;
      RECT 1205 204455 1375 204625 ;
    LAYER V1 ;
      RECT 1205 206135 1375 206305 ;
    LAYER V1 ;
      RECT 1205 210335 1375 210505 ;
    LAYER V1 ;
      RECT 1205 212015 1375 212185 ;
    LAYER V1 ;
      RECT 1205 216215 1375 216385 ;
    LAYER V1 ;
      RECT 1205 217895 1375 218065 ;
    LAYER V1 ;
      RECT 1205 222095 1375 222265 ;
    LAYER V1 ;
      RECT 1205 223775 1375 223945 ;
    LAYER V1 ;
      RECT 1205 227975 1375 228145 ;
    LAYER V1 ;
      RECT 1205 229655 1375 229825 ;
    LAYER V1 ;
      RECT 1205 233855 1375 234025 ;
    LAYER V1 ;
      RECT 1205 235535 1375 235705 ;
    LAYER V1 ;
      RECT 1205 239735 1375 239905 ;
    LAYER V1 ;
      RECT 1205 241415 1375 241585 ;
    LAYER V1 ;
      RECT 1205 245615 1375 245785 ;
    LAYER V1 ;
      RECT 1205 247295 1375 247465 ;
    LAYER V1 ;
      RECT 1205 251495 1375 251665 ;
    LAYER V1 ;
      RECT 1205 253175 1375 253345 ;
    LAYER V1 ;
      RECT 1205 257375 1375 257545 ;
    LAYER V1 ;
      RECT 1205 259055 1375 259225 ;
    LAYER V1 ;
      RECT 1205 263255 1375 263425 ;
    LAYER V1 ;
      RECT 1205 264935 1375 265105 ;
    LAYER V1 ;
      RECT 1205 269135 1375 269305 ;
    LAYER V1 ;
      RECT 1205 270815 1375 270985 ;
    LAYER V1 ;
      RECT 1205 275015 1375 275185 ;
    LAYER V1 ;
      RECT 1205 276695 1375 276865 ;
    LAYER V1 ;
      RECT 1205 280895 1375 281065 ;
    LAYER V1 ;
      RECT 1205 282575 1375 282745 ;
    LAYER V1 ;
      RECT 1205 286775 1375 286945 ;
    LAYER V1 ;
      RECT 1205 288455 1375 288625 ;
    LAYER V1 ;
      RECT 1205 292655 1375 292825 ;
    LAYER V1 ;
      RECT 1205 294335 1375 294505 ;
    LAYER V1 ;
      RECT 1205 298535 1375 298705 ;
    LAYER V1 ;
      RECT 1205 300215 1375 300385 ;
    LAYER V1 ;
      RECT 1205 304415 1375 304585 ;
    LAYER V1 ;
      RECT 1205 306095 1375 306265 ;
    LAYER V1 ;
      RECT 1205 310295 1375 310465 ;
    LAYER V1 ;
      RECT 1205 311975 1375 312145 ;
    LAYER V1 ;
      RECT 1205 316175 1375 316345 ;
    LAYER V1 ;
      RECT 1205 317855 1375 318025 ;
    LAYER V1 ;
      RECT 1205 322055 1375 322225 ;
    LAYER V1 ;
      RECT 1205 323735 1375 323905 ;
    LAYER V1 ;
      RECT 1205 327935 1375 328105 ;
    LAYER V1 ;
      RECT 1205 329615 1375 329785 ;
    LAYER V1 ;
      RECT 1205 333815 1375 333985 ;
    LAYER V1 ;
      RECT 1205 335495 1375 335665 ;
    LAYER V1 ;
      RECT 1205 339695 1375 339865 ;
    LAYER V1 ;
      RECT 1205 341375 1375 341545 ;
    LAYER V1 ;
      RECT 1205 345575 1375 345745 ;
    LAYER V1 ;
      RECT 1205 347255 1375 347425 ;
    LAYER V1 ;
      RECT 1205 351455 1375 351625 ;
    LAYER V1 ;
      RECT 1205 353135 1375 353305 ;
    LAYER V1 ;
      RECT 1205 357335 1375 357505 ;
    LAYER V1 ;
      RECT 1205 359015 1375 359185 ;
    LAYER V1 ;
      RECT 1205 363215 1375 363385 ;
    LAYER V1 ;
      RECT 1205 364895 1375 365065 ;
    LAYER V1 ;
      RECT 1205 369095 1375 369265 ;
    LAYER V1 ;
      RECT 1205 370775 1375 370945 ;
    LAYER V1 ;
      RECT 1205 374975 1375 375145 ;
    LAYER V1 ;
      RECT 1205 376655 1375 376825 ;
    LAYER V1 ;
      RECT 1205 380855 1375 381025 ;
    LAYER V1 ;
      RECT 1205 382535 1375 382705 ;
    LAYER V1 ;
      RECT 1205 386735 1375 386905 ;
    LAYER V1 ;
      RECT 1205 388415 1375 388585 ;
    LAYER V1 ;
      RECT 1205 392615 1375 392785 ;
    LAYER V1 ;
      RECT 1205 394295 1375 394465 ;
    LAYER V1 ;
      RECT 1205 398495 1375 398665 ;
    LAYER V1 ;
      RECT 1205 400175 1375 400345 ;
    LAYER V1 ;
      RECT 1205 404375 1375 404545 ;
    LAYER V1 ;
      RECT 1205 406055 1375 406225 ;
    LAYER V1 ;
      RECT 1205 410255 1375 410425 ;
    LAYER V1 ;
      RECT 1205 411935 1375 412105 ;
    LAYER V1 ;
      RECT 1205 416135 1375 416305 ;
    LAYER V1 ;
      RECT 1205 417815 1375 417985 ;
    LAYER V1 ;
      RECT 1205 422015 1375 422185 ;
    LAYER V1 ;
      RECT 1205 423695 1375 423865 ;
    LAYER V1 ;
      RECT 1205 427895 1375 428065 ;
    LAYER V1 ;
      RECT 1205 429575 1375 429745 ;
    LAYER V1 ;
      RECT 1205 433775 1375 433945 ;
    LAYER V1 ;
      RECT 1205 435455 1375 435625 ;
    LAYER V1 ;
      RECT 1205 439655 1375 439825 ;
    LAYER V1 ;
      RECT 1205 441335 1375 441505 ;
    LAYER V1 ;
      RECT 1205 445535 1375 445705 ;
    LAYER V1 ;
      RECT 1205 447215 1375 447385 ;
    LAYER V1 ;
      RECT 1205 451415 1375 451585 ;
    LAYER V1 ;
      RECT 1205 453095 1375 453265 ;
    LAYER V1 ;
      RECT 1205 457295 1375 457465 ;
    LAYER V1 ;
      RECT 1205 458975 1375 459145 ;
    LAYER V1 ;
      RECT 1205 463175 1375 463345 ;
    LAYER V1 ;
      RECT 1205 464855 1375 465025 ;
    LAYER V1 ;
      RECT 1205 469055 1375 469225 ;
    LAYER V1 ;
      RECT 1205 470735 1375 470905 ;
    LAYER V1 ;
      RECT 1205 474935 1375 475105 ;
    LAYER V1 ;
      RECT 1205 476615 1375 476785 ;
    LAYER V1 ;
      RECT 1205 480815 1375 480985 ;
    LAYER V1 ;
      RECT 1205 482495 1375 482665 ;
    LAYER V1 ;
      RECT 1205 486695 1375 486865 ;
    LAYER V1 ;
      RECT 1205 488375 1375 488545 ;
    LAYER V1 ;
      RECT 1205 492575 1375 492745 ;
    LAYER V1 ;
      RECT 1205 494255 1375 494425 ;
    LAYER V1 ;
      RECT 1205 498455 1375 498625 ;
    LAYER V1 ;
      RECT 1205 500135 1375 500305 ;
    LAYER V1 ;
      RECT 1205 504335 1375 504505 ;
    LAYER V1 ;
      RECT 1205 506015 1375 506185 ;
    LAYER V1 ;
      RECT 1205 510215 1375 510385 ;
    LAYER V1 ;
      RECT 1205 511895 1375 512065 ;
    LAYER V1 ;
      RECT 1205 516095 1375 516265 ;
    LAYER V1 ;
      RECT 1205 517775 1375 517945 ;
    LAYER V1 ;
      RECT 1205 521975 1375 522145 ;
    LAYER V1 ;
      RECT 1205 523655 1375 523825 ;
    LAYER V1 ;
      RECT 1205 527855 1375 528025 ;
    LAYER V1 ;
      RECT 1205 529535 1375 529705 ;
    LAYER V1 ;
      RECT 1205 533735 1375 533905 ;
    LAYER V1 ;
      RECT 1205 535415 1375 535585 ;
    LAYER V1 ;
      RECT 1205 539615 1375 539785 ;
    LAYER V1 ;
      RECT 1205 541295 1375 541465 ;
    LAYER V1 ;
      RECT 1205 545495 1375 545665 ;
    LAYER V1 ;
      RECT 1205 547175 1375 547345 ;
    LAYER V1 ;
      RECT 1205 551375 1375 551545 ;
    LAYER V1 ;
      RECT 1205 553055 1375 553225 ;
    LAYER V1 ;
      RECT 1205 557255 1375 557425 ;
    LAYER V1 ;
      RECT 1205 558935 1375 559105 ;
    LAYER V1 ;
      RECT 1205 563135 1375 563305 ;
    LAYER V1 ;
      RECT 1205 564815 1375 564985 ;
    LAYER V1 ;
      RECT 1205 569015 1375 569185 ;
    LAYER V1 ;
      RECT 1205 570695 1375 570865 ;
    LAYER V1 ;
      RECT 1205 574895 1375 575065 ;
    LAYER V1 ;
      RECT 1205 576575 1375 576745 ;
    LAYER V1 ;
      RECT 1205 580775 1375 580945 ;
    LAYER V1 ;
      RECT 1205 582455 1375 582625 ;
    LAYER V1 ;
      RECT 1205 586655 1375 586825 ;
    LAYER V1 ;
      RECT 1205 588335 1375 588505 ;
    LAYER V1 ;
      RECT 1205 592535 1375 592705 ;
    LAYER V1 ;
      RECT 1205 594215 1375 594385 ;
    LAYER V1 ;
      RECT 1205 598415 1375 598585 ;
    LAYER V1 ;
      RECT 1205 600095 1375 600265 ;
    LAYER V1 ;
      RECT 1205 604295 1375 604465 ;
    LAYER V1 ;
      RECT 1205 605975 1375 606145 ;
    LAYER V1 ;
      RECT 1205 610175 1375 610345 ;
    LAYER V1 ;
      RECT 1205 611855 1375 612025 ;
    LAYER V1 ;
      RECT 1205 616055 1375 616225 ;
    LAYER V1 ;
      RECT 1205 617735 1375 617905 ;
    LAYER V1 ;
      RECT 1205 621935 1375 622105 ;
    LAYER V1 ;
      RECT 1205 623615 1375 623785 ;
    LAYER V1 ;
      RECT 1205 627815 1375 627985 ;
    LAYER V1 ;
      RECT 1205 629495 1375 629665 ;
    LAYER V1 ;
      RECT 1205 633695 1375 633865 ;
    LAYER V1 ;
      RECT 1205 635375 1375 635545 ;
    LAYER V1 ;
      RECT 1205 639575 1375 639745 ;
    LAYER V1 ;
      RECT 1205 641255 1375 641425 ;
    LAYER V1 ;
      RECT 1205 645455 1375 645625 ;
    LAYER V1 ;
      RECT 1205 647135 1375 647305 ;
    LAYER V1 ;
      RECT 1205 651335 1375 651505 ;
    LAYER V1 ;
      RECT 1205 653015 1375 653185 ;
    LAYER V1 ;
      RECT 1205 657215 1375 657385 ;
    LAYER V1 ;
      RECT 1205 658895 1375 659065 ;
    LAYER V1 ;
      RECT 1205 663095 1375 663265 ;
    LAYER V1 ;
      RECT 1205 664775 1375 664945 ;
    LAYER V1 ;
      RECT 1205 668975 1375 669145 ;
    LAYER V1 ;
      RECT 1205 670655 1375 670825 ;
    LAYER V1 ;
      RECT 1205 674855 1375 675025 ;
    LAYER V1 ;
      RECT 1205 676535 1375 676705 ;
    LAYER V1 ;
      RECT 1205 680735 1375 680905 ;
    LAYER V1 ;
      RECT 1205 682415 1375 682585 ;
    LAYER V1 ;
      RECT 1205 686615 1375 686785 ;
    LAYER V1 ;
      RECT 1205 688295 1375 688465 ;
    LAYER V1 ;
      RECT 1205 692495 1375 692665 ;
    LAYER V1 ;
      RECT 1205 694175 1375 694345 ;
    LAYER V1 ;
      RECT 1205 698375 1375 698545 ;
    LAYER V1 ;
      RECT 1205 700055 1375 700225 ;
    LAYER V1 ;
      RECT 1205 704255 1375 704425 ;
    LAYER V1 ;
      RECT 1205 705935 1375 706105 ;
    LAYER V1 ;
      RECT 1205 710135 1375 710305 ;
    LAYER V1 ;
      RECT 1205 711815 1375 711985 ;
    LAYER V1 ;
      RECT 1205 716015 1375 716185 ;
    LAYER V1 ;
      RECT 1205 717695 1375 717865 ;
    LAYER V1 ;
      RECT 1205 721895 1375 722065 ;
    LAYER V1 ;
      RECT 1205 723575 1375 723745 ;
    LAYER V1 ;
      RECT 1205 727775 1375 727945 ;
    LAYER V1 ;
      RECT 1205 729455 1375 729625 ;
    LAYER V1 ;
      RECT 1205 733655 1375 733825 ;
    LAYER V1 ;
      RECT 1205 735335 1375 735505 ;
    LAYER V1 ;
      RECT 1205 739535 1375 739705 ;
    LAYER V1 ;
      RECT 1205 741215 1375 741385 ;
    LAYER V1 ;
      RECT 1205 745415 1375 745585 ;
    LAYER V1 ;
      RECT 1205 747095 1375 747265 ;
    LAYER V1 ;
      RECT 1205 751295 1375 751465 ;
    LAYER V1 ;
      RECT 1205 752975 1375 753145 ;
    LAYER V1 ;
      RECT 1205 757175 1375 757345 ;
    LAYER V1 ;
      RECT 1205 758855 1375 759025 ;
    LAYER V1 ;
      RECT 1205 763055 1375 763225 ;
    LAYER V1 ;
      RECT 1205 764735 1375 764905 ;
    LAYER V1 ;
      RECT 1205 768935 1375 769105 ;
    LAYER V1 ;
      RECT 1205 770615 1375 770785 ;
    LAYER V1 ;
      RECT 1205 774815 1375 774985 ;
    LAYER V1 ;
      RECT 1205 776495 1375 776665 ;
    LAYER V1 ;
      RECT 1205 780695 1375 780865 ;
    LAYER V1 ;
      RECT 1205 782375 1375 782545 ;
    LAYER V1 ;
      RECT 1205 786575 1375 786745 ;
    LAYER V1 ;
      RECT 1205 788255 1375 788425 ;
    LAYER V1 ;
      RECT 1205 792455 1375 792625 ;
    LAYER V1 ;
      RECT 1205 794135 1375 794305 ;
    LAYER V1 ;
      RECT 1205 798335 1375 798505 ;
    LAYER V1 ;
      RECT 1205 800015 1375 800185 ;
    LAYER V1 ;
      RECT 1205 804215 1375 804385 ;
    LAYER V1 ;
      RECT 1205 805895 1375 806065 ;
    LAYER V1 ;
      RECT 1205 810095 1375 810265 ;
    LAYER V1 ;
      RECT 1205 811775 1375 811945 ;
    LAYER V1 ;
      RECT 1205 815975 1375 816145 ;
    LAYER V1 ;
      RECT 1205 817655 1375 817825 ;
    LAYER V1 ;
      RECT 1205 821855 1375 822025 ;
    LAYER V1 ;
      RECT 1205 823535 1375 823705 ;
    LAYER V1 ;
      RECT 1205 827735 1375 827905 ;
    LAYER V1 ;
      RECT 1205 829415 1375 829585 ;
    LAYER V1 ;
      RECT 1205 833615 1375 833785 ;
    LAYER V1 ;
      RECT 1205 835295 1375 835465 ;
    LAYER V1 ;
      RECT 1205 839495 1375 839665 ;
    LAYER V1 ;
      RECT 1205 841175 1375 841345 ;
    LAYER V1 ;
      RECT 1205 845375 1375 845545 ;
    LAYER V1 ;
      RECT 1205 847055 1375 847225 ;
    LAYER V1 ;
      RECT 1205 851255 1375 851425 ;
    LAYER V1 ;
      RECT 1205 852935 1375 853105 ;
    LAYER V1 ;
      RECT 1205 857135 1375 857305 ;
    LAYER V1 ;
      RECT 1205 858815 1375 858985 ;
    LAYER V1 ;
      RECT 1205 863015 1375 863185 ;
    LAYER V1 ;
      RECT 1205 864695 1375 864865 ;
    LAYER V1 ;
      RECT 1205 868895 1375 869065 ;
    LAYER V1 ;
      RECT 1205 870995 1375 871165 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 775 53675 945 53845 ;
    LAYER V1 ;
      RECT 775 59555 945 59725 ;
    LAYER V1 ;
      RECT 775 65435 945 65605 ;
    LAYER V1 ;
      RECT 775 71315 945 71485 ;
    LAYER V1 ;
      RECT 775 77195 945 77365 ;
    LAYER V1 ;
      RECT 775 83075 945 83245 ;
    LAYER V1 ;
      RECT 775 88955 945 89125 ;
    LAYER V1 ;
      RECT 775 94835 945 95005 ;
    LAYER V1 ;
      RECT 775 100715 945 100885 ;
    LAYER V1 ;
      RECT 775 106595 945 106765 ;
    LAYER V1 ;
      RECT 775 112475 945 112645 ;
    LAYER V1 ;
      RECT 775 118355 945 118525 ;
    LAYER V1 ;
      RECT 775 124235 945 124405 ;
    LAYER V1 ;
      RECT 775 130115 945 130285 ;
    LAYER V1 ;
      RECT 775 135995 945 136165 ;
    LAYER V1 ;
      RECT 775 141875 945 142045 ;
    LAYER V1 ;
      RECT 775 147755 945 147925 ;
    LAYER V1 ;
      RECT 775 153635 945 153805 ;
    LAYER V1 ;
      RECT 775 159515 945 159685 ;
    LAYER V1 ;
      RECT 775 165395 945 165565 ;
    LAYER V1 ;
      RECT 775 171275 945 171445 ;
    LAYER V1 ;
      RECT 775 177155 945 177325 ;
    LAYER V1 ;
      RECT 775 183035 945 183205 ;
    LAYER V1 ;
      RECT 775 188915 945 189085 ;
    LAYER V1 ;
      RECT 775 194795 945 194965 ;
    LAYER V1 ;
      RECT 775 200675 945 200845 ;
    LAYER V1 ;
      RECT 775 206555 945 206725 ;
    LAYER V1 ;
      RECT 775 212435 945 212605 ;
    LAYER V1 ;
      RECT 775 218315 945 218485 ;
    LAYER V1 ;
      RECT 775 224195 945 224365 ;
    LAYER V1 ;
      RECT 775 230075 945 230245 ;
    LAYER V1 ;
      RECT 775 235955 945 236125 ;
    LAYER V1 ;
      RECT 775 241835 945 242005 ;
    LAYER V1 ;
      RECT 775 247715 945 247885 ;
    LAYER V1 ;
      RECT 775 253595 945 253765 ;
    LAYER V1 ;
      RECT 775 259475 945 259645 ;
    LAYER V1 ;
      RECT 775 265355 945 265525 ;
    LAYER V1 ;
      RECT 775 271235 945 271405 ;
    LAYER V1 ;
      RECT 775 277115 945 277285 ;
    LAYER V1 ;
      RECT 775 282995 945 283165 ;
    LAYER V1 ;
      RECT 775 288875 945 289045 ;
    LAYER V1 ;
      RECT 775 294755 945 294925 ;
    LAYER V1 ;
      RECT 775 300635 945 300805 ;
    LAYER V1 ;
      RECT 775 306515 945 306685 ;
    LAYER V1 ;
      RECT 775 312395 945 312565 ;
    LAYER V1 ;
      RECT 775 318275 945 318445 ;
    LAYER V1 ;
      RECT 775 324155 945 324325 ;
    LAYER V1 ;
      RECT 775 330035 945 330205 ;
    LAYER V1 ;
      RECT 775 335915 945 336085 ;
    LAYER V1 ;
      RECT 775 341795 945 341965 ;
    LAYER V1 ;
      RECT 775 347675 945 347845 ;
    LAYER V1 ;
      RECT 775 353555 945 353725 ;
    LAYER V1 ;
      RECT 775 359435 945 359605 ;
    LAYER V1 ;
      RECT 775 365315 945 365485 ;
    LAYER V1 ;
      RECT 775 371195 945 371365 ;
    LAYER V1 ;
      RECT 775 377075 945 377245 ;
    LAYER V1 ;
      RECT 775 382955 945 383125 ;
    LAYER V1 ;
      RECT 775 388835 945 389005 ;
    LAYER V1 ;
      RECT 775 394715 945 394885 ;
    LAYER V1 ;
      RECT 775 400595 945 400765 ;
    LAYER V1 ;
      RECT 775 406475 945 406645 ;
    LAYER V1 ;
      RECT 775 412355 945 412525 ;
    LAYER V1 ;
      RECT 775 418235 945 418405 ;
    LAYER V1 ;
      RECT 775 424115 945 424285 ;
    LAYER V1 ;
      RECT 775 429995 945 430165 ;
    LAYER V1 ;
      RECT 775 435875 945 436045 ;
    LAYER V1 ;
      RECT 775 441755 945 441925 ;
    LAYER V1 ;
      RECT 775 447635 945 447805 ;
    LAYER V1 ;
      RECT 775 453515 945 453685 ;
    LAYER V1 ;
      RECT 775 459395 945 459565 ;
    LAYER V1 ;
      RECT 775 465275 945 465445 ;
    LAYER V1 ;
      RECT 775 471155 945 471325 ;
    LAYER V1 ;
      RECT 775 477035 945 477205 ;
    LAYER V1 ;
      RECT 775 482915 945 483085 ;
    LAYER V1 ;
      RECT 775 488795 945 488965 ;
    LAYER V1 ;
      RECT 775 494675 945 494845 ;
    LAYER V1 ;
      RECT 775 500555 945 500725 ;
    LAYER V1 ;
      RECT 775 506435 945 506605 ;
    LAYER V1 ;
      RECT 775 512315 945 512485 ;
    LAYER V1 ;
      RECT 775 518195 945 518365 ;
    LAYER V1 ;
      RECT 775 524075 945 524245 ;
    LAYER V1 ;
      RECT 775 529955 945 530125 ;
    LAYER V1 ;
      RECT 775 535835 945 536005 ;
    LAYER V1 ;
      RECT 775 541715 945 541885 ;
    LAYER V1 ;
      RECT 775 547595 945 547765 ;
    LAYER V1 ;
      RECT 775 553475 945 553645 ;
    LAYER V1 ;
      RECT 775 559355 945 559525 ;
    LAYER V1 ;
      RECT 775 565235 945 565405 ;
    LAYER V1 ;
      RECT 775 571115 945 571285 ;
    LAYER V1 ;
      RECT 775 576995 945 577165 ;
    LAYER V1 ;
      RECT 775 582875 945 583045 ;
    LAYER V1 ;
      RECT 775 588755 945 588925 ;
    LAYER V1 ;
      RECT 775 594635 945 594805 ;
    LAYER V1 ;
      RECT 775 600515 945 600685 ;
    LAYER V1 ;
      RECT 775 606395 945 606565 ;
    LAYER V1 ;
      RECT 775 612275 945 612445 ;
    LAYER V1 ;
      RECT 775 618155 945 618325 ;
    LAYER V1 ;
      RECT 775 624035 945 624205 ;
    LAYER V1 ;
      RECT 775 629915 945 630085 ;
    LAYER V1 ;
      RECT 775 635795 945 635965 ;
    LAYER V1 ;
      RECT 775 641675 945 641845 ;
    LAYER V1 ;
      RECT 775 647555 945 647725 ;
    LAYER V1 ;
      RECT 775 653435 945 653605 ;
    LAYER V1 ;
      RECT 775 659315 945 659485 ;
    LAYER V1 ;
      RECT 775 665195 945 665365 ;
    LAYER V1 ;
      RECT 775 671075 945 671245 ;
    LAYER V1 ;
      RECT 775 676955 945 677125 ;
    LAYER V1 ;
      RECT 775 682835 945 683005 ;
    LAYER V1 ;
      RECT 775 688715 945 688885 ;
    LAYER V1 ;
      RECT 775 694595 945 694765 ;
    LAYER V1 ;
      RECT 775 700475 945 700645 ;
    LAYER V1 ;
      RECT 775 706355 945 706525 ;
    LAYER V1 ;
      RECT 775 712235 945 712405 ;
    LAYER V1 ;
      RECT 775 718115 945 718285 ;
    LAYER V1 ;
      RECT 775 723995 945 724165 ;
    LAYER V1 ;
      RECT 775 729875 945 730045 ;
    LAYER V1 ;
      RECT 775 735755 945 735925 ;
    LAYER V1 ;
      RECT 775 741635 945 741805 ;
    LAYER V1 ;
      RECT 775 747515 945 747685 ;
    LAYER V1 ;
      RECT 775 753395 945 753565 ;
    LAYER V1 ;
      RECT 775 759275 945 759445 ;
    LAYER V1 ;
      RECT 775 765155 945 765325 ;
    LAYER V1 ;
      RECT 775 771035 945 771205 ;
    LAYER V1 ;
      RECT 775 776915 945 777085 ;
    LAYER V1 ;
      RECT 775 782795 945 782965 ;
    LAYER V1 ;
      RECT 775 788675 945 788845 ;
    LAYER V1 ;
      RECT 775 794555 945 794725 ;
    LAYER V1 ;
      RECT 775 800435 945 800605 ;
    LAYER V1 ;
      RECT 775 806315 945 806485 ;
    LAYER V1 ;
      RECT 775 812195 945 812365 ;
    LAYER V1 ;
      RECT 775 818075 945 818245 ;
    LAYER V1 ;
      RECT 775 823955 945 824125 ;
    LAYER V1 ;
      RECT 775 829835 945 830005 ;
    LAYER V1 ;
      RECT 775 835715 945 835885 ;
    LAYER V1 ;
      RECT 775 841595 945 841765 ;
    LAYER V1 ;
      RECT 775 847475 945 847645 ;
    LAYER V1 ;
      RECT 775 853355 945 853525 ;
    LAYER V1 ;
      RECT 775 859235 945 859405 ;
    LAYER V1 ;
      RECT 775 865115 945 865285 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 1635 53675 1805 53845 ;
    LAYER V1 ;
      RECT 1635 59555 1805 59725 ;
    LAYER V1 ;
      RECT 1635 65435 1805 65605 ;
    LAYER V1 ;
      RECT 1635 71315 1805 71485 ;
    LAYER V1 ;
      RECT 1635 77195 1805 77365 ;
    LAYER V1 ;
      RECT 1635 83075 1805 83245 ;
    LAYER V1 ;
      RECT 1635 88955 1805 89125 ;
    LAYER V1 ;
      RECT 1635 94835 1805 95005 ;
    LAYER V1 ;
      RECT 1635 100715 1805 100885 ;
    LAYER V1 ;
      RECT 1635 106595 1805 106765 ;
    LAYER V1 ;
      RECT 1635 112475 1805 112645 ;
    LAYER V1 ;
      RECT 1635 118355 1805 118525 ;
    LAYER V1 ;
      RECT 1635 124235 1805 124405 ;
    LAYER V1 ;
      RECT 1635 130115 1805 130285 ;
    LAYER V1 ;
      RECT 1635 135995 1805 136165 ;
    LAYER V1 ;
      RECT 1635 141875 1805 142045 ;
    LAYER V1 ;
      RECT 1635 147755 1805 147925 ;
    LAYER V1 ;
      RECT 1635 153635 1805 153805 ;
    LAYER V1 ;
      RECT 1635 159515 1805 159685 ;
    LAYER V1 ;
      RECT 1635 165395 1805 165565 ;
    LAYER V1 ;
      RECT 1635 171275 1805 171445 ;
    LAYER V1 ;
      RECT 1635 177155 1805 177325 ;
    LAYER V1 ;
      RECT 1635 183035 1805 183205 ;
    LAYER V1 ;
      RECT 1635 188915 1805 189085 ;
    LAYER V1 ;
      RECT 1635 194795 1805 194965 ;
    LAYER V1 ;
      RECT 1635 200675 1805 200845 ;
    LAYER V1 ;
      RECT 1635 206555 1805 206725 ;
    LAYER V1 ;
      RECT 1635 212435 1805 212605 ;
    LAYER V1 ;
      RECT 1635 218315 1805 218485 ;
    LAYER V1 ;
      RECT 1635 224195 1805 224365 ;
    LAYER V1 ;
      RECT 1635 230075 1805 230245 ;
    LAYER V1 ;
      RECT 1635 235955 1805 236125 ;
    LAYER V1 ;
      RECT 1635 241835 1805 242005 ;
    LAYER V1 ;
      RECT 1635 247715 1805 247885 ;
    LAYER V1 ;
      RECT 1635 253595 1805 253765 ;
    LAYER V1 ;
      RECT 1635 259475 1805 259645 ;
    LAYER V1 ;
      RECT 1635 265355 1805 265525 ;
    LAYER V1 ;
      RECT 1635 271235 1805 271405 ;
    LAYER V1 ;
      RECT 1635 277115 1805 277285 ;
    LAYER V1 ;
      RECT 1635 282995 1805 283165 ;
    LAYER V1 ;
      RECT 1635 288875 1805 289045 ;
    LAYER V1 ;
      RECT 1635 294755 1805 294925 ;
    LAYER V1 ;
      RECT 1635 300635 1805 300805 ;
    LAYER V1 ;
      RECT 1635 306515 1805 306685 ;
    LAYER V1 ;
      RECT 1635 312395 1805 312565 ;
    LAYER V1 ;
      RECT 1635 318275 1805 318445 ;
    LAYER V1 ;
      RECT 1635 324155 1805 324325 ;
    LAYER V1 ;
      RECT 1635 330035 1805 330205 ;
    LAYER V1 ;
      RECT 1635 335915 1805 336085 ;
    LAYER V1 ;
      RECT 1635 341795 1805 341965 ;
    LAYER V1 ;
      RECT 1635 347675 1805 347845 ;
    LAYER V1 ;
      RECT 1635 353555 1805 353725 ;
    LAYER V1 ;
      RECT 1635 359435 1805 359605 ;
    LAYER V1 ;
      RECT 1635 365315 1805 365485 ;
    LAYER V1 ;
      RECT 1635 371195 1805 371365 ;
    LAYER V1 ;
      RECT 1635 377075 1805 377245 ;
    LAYER V1 ;
      RECT 1635 382955 1805 383125 ;
    LAYER V1 ;
      RECT 1635 388835 1805 389005 ;
    LAYER V1 ;
      RECT 1635 394715 1805 394885 ;
    LAYER V1 ;
      RECT 1635 400595 1805 400765 ;
    LAYER V1 ;
      RECT 1635 406475 1805 406645 ;
    LAYER V1 ;
      RECT 1635 412355 1805 412525 ;
    LAYER V1 ;
      RECT 1635 418235 1805 418405 ;
    LAYER V1 ;
      RECT 1635 424115 1805 424285 ;
    LAYER V1 ;
      RECT 1635 429995 1805 430165 ;
    LAYER V1 ;
      RECT 1635 435875 1805 436045 ;
    LAYER V1 ;
      RECT 1635 441755 1805 441925 ;
    LAYER V1 ;
      RECT 1635 447635 1805 447805 ;
    LAYER V1 ;
      RECT 1635 453515 1805 453685 ;
    LAYER V1 ;
      RECT 1635 459395 1805 459565 ;
    LAYER V1 ;
      RECT 1635 465275 1805 465445 ;
    LAYER V1 ;
      RECT 1635 471155 1805 471325 ;
    LAYER V1 ;
      RECT 1635 477035 1805 477205 ;
    LAYER V1 ;
      RECT 1635 482915 1805 483085 ;
    LAYER V1 ;
      RECT 1635 488795 1805 488965 ;
    LAYER V1 ;
      RECT 1635 494675 1805 494845 ;
    LAYER V1 ;
      RECT 1635 500555 1805 500725 ;
    LAYER V1 ;
      RECT 1635 506435 1805 506605 ;
    LAYER V1 ;
      RECT 1635 512315 1805 512485 ;
    LAYER V1 ;
      RECT 1635 518195 1805 518365 ;
    LAYER V1 ;
      RECT 1635 524075 1805 524245 ;
    LAYER V1 ;
      RECT 1635 529955 1805 530125 ;
    LAYER V1 ;
      RECT 1635 535835 1805 536005 ;
    LAYER V1 ;
      RECT 1635 541715 1805 541885 ;
    LAYER V1 ;
      RECT 1635 547595 1805 547765 ;
    LAYER V1 ;
      RECT 1635 553475 1805 553645 ;
    LAYER V1 ;
      RECT 1635 559355 1805 559525 ;
    LAYER V1 ;
      RECT 1635 565235 1805 565405 ;
    LAYER V1 ;
      RECT 1635 571115 1805 571285 ;
    LAYER V1 ;
      RECT 1635 576995 1805 577165 ;
    LAYER V1 ;
      RECT 1635 582875 1805 583045 ;
    LAYER V1 ;
      RECT 1635 588755 1805 588925 ;
    LAYER V1 ;
      RECT 1635 594635 1805 594805 ;
    LAYER V1 ;
      RECT 1635 600515 1805 600685 ;
    LAYER V1 ;
      RECT 1635 606395 1805 606565 ;
    LAYER V1 ;
      RECT 1635 612275 1805 612445 ;
    LAYER V1 ;
      RECT 1635 618155 1805 618325 ;
    LAYER V1 ;
      RECT 1635 624035 1805 624205 ;
    LAYER V1 ;
      RECT 1635 629915 1805 630085 ;
    LAYER V1 ;
      RECT 1635 635795 1805 635965 ;
    LAYER V1 ;
      RECT 1635 641675 1805 641845 ;
    LAYER V1 ;
      RECT 1635 647555 1805 647725 ;
    LAYER V1 ;
      RECT 1635 653435 1805 653605 ;
    LAYER V1 ;
      RECT 1635 659315 1805 659485 ;
    LAYER V1 ;
      RECT 1635 665195 1805 665365 ;
    LAYER V1 ;
      RECT 1635 671075 1805 671245 ;
    LAYER V1 ;
      RECT 1635 676955 1805 677125 ;
    LAYER V1 ;
      RECT 1635 682835 1805 683005 ;
    LAYER V1 ;
      RECT 1635 688715 1805 688885 ;
    LAYER V1 ;
      RECT 1635 694595 1805 694765 ;
    LAYER V1 ;
      RECT 1635 700475 1805 700645 ;
    LAYER V1 ;
      RECT 1635 706355 1805 706525 ;
    LAYER V1 ;
      RECT 1635 712235 1805 712405 ;
    LAYER V1 ;
      RECT 1635 718115 1805 718285 ;
    LAYER V1 ;
      RECT 1635 723995 1805 724165 ;
    LAYER V1 ;
      RECT 1635 729875 1805 730045 ;
    LAYER V1 ;
      RECT 1635 735755 1805 735925 ;
    LAYER V1 ;
      RECT 1635 741635 1805 741805 ;
    LAYER V1 ;
      RECT 1635 747515 1805 747685 ;
    LAYER V1 ;
      RECT 1635 753395 1805 753565 ;
    LAYER V1 ;
      RECT 1635 759275 1805 759445 ;
    LAYER V1 ;
      RECT 1635 765155 1805 765325 ;
    LAYER V1 ;
      RECT 1635 771035 1805 771205 ;
    LAYER V1 ;
      RECT 1635 776915 1805 777085 ;
    LAYER V1 ;
      RECT 1635 782795 1805 782965 ;
    LAYER V1 ;
      RECT 1635 788675 1805 788845 ;
    LAYER V1 ;
      RECT 1635 794555 1805 794725 ;
    LAYER V1 ;
      RECT 1635 800435 1805 800605 ;
    LAYER V1 ;
      RECT 1635 806315 1805 806485 ;
    LAYER V1 ;
      RECT 1635 812195 1805 812365 ;
    LAYER V1 ;
      RECT 1635 818075 1805 818245 ;
    LAYER V1 ;
      RECT 1635 823955 1805 824125 ;
    LAYER V1 ;
      RECT 1635 829835 1805 830005 ;
    LAYER V1 ;
      RECT 1635 835715 1805 835885 ;
    LAYER V1 ;
      RECT 1635 841595 1805 841765 ;
    LAYER V1 ;
      RECT 1635 847475 1805 847645 ;
    LAYER V1 ;
      RECT 1635 853355 1805 853525 ;
    LAYER V1 ;
      RECT 1635 859235 1805 859405 ;
    LAYER V1 ;
      RECT 1635 865115 1805 865285 ;
    LAYER V2 ;
      RECT 785 345 935 495 ;
    LAYER V2 ;
      RECT 785 6225 935 6375 ;
    LAYER V2 ;
      RECT 785 12105 935 12255 ;
    LAYER V2 ;
      RECT 785 17985 935 18135 ;
    LAYER V2 ;
      RECT 785 23865 935 24015 ;
    LAYER V2 ;
      RECT 785 29745 935 29895 ;
    LAYER V2 ;
      RECT 785 35625 935 35775 ;
    LAYER V2 ;
      RECT 785 41505 935 41655 ;
    LAYER V2 ;
      RECT 785 47385 935 47535 ;
    LAYER V2 ;
      RECT 785 53265 935 53415 ;
    LAYER V2 ;
      RECT 785 59145 935 59295 ;
    LAYER V2 ;
      RECT 785 65025 935 65175 ;
    LAYER V2 ;
      RECT 785 70905 935 71055 ;
    LAYER V2 ;
      RECT 785 76785 935 76935 ;
    LAYER V2 ;
      RECT 785 82665 935 82815 ;
    LAYER V2 ;
      RECT 785 88545 935 88695 ;
    LAYER V2 ;
      RECT 785 94425 935 94575 ;
    LAYER V2 ;
      RECT 785 100305 935 100455 ;
    LAYER V2 ;
      RECT 785 106185 935 106335 ;
    LAYER V2 ;
      RECT 785 112065 935 112215 ;
    LAYER V2 ;
      RECT 785 117945 935 118095 ;
    LAYER V2 ;
      RECT 785 123825 935 123975 ;
    LAYER V2 ;
      RECT 785 129705 935 129855 ;
    LAYER V2 ;
      RECT 785 135585 935 135735 ;
    LAYER V2 ;
      RECT 785 141465 935 141615 ;
    LAYER V2 ;
      RECT 785 147345 935 147495 ;
    LAYER V2 ;
      RECT 785 153225 935 153375 ;
    LAYER V2 ;
      RECT 785 159105 935 159255 ;
    LAYER V2 ;
      RECT 785 164985 935 165135 ;
    LAYER V2 ;
      RECT 785 170865 935 171015 ;
    LAYER V2 ;
      RECT 785 176745 935 176895 ;
    LAYER V2 ;
      RECT 785 182625 935 182775 ;
    LAYER V2 ;
      RECT 785 188505 935 188655 ;
    LAYER V2 ;
      RECT 785 194385 935 194535 ;
    LAYER V2 ;
      RECT 785 200265 935 200415 ;
    LAYER V2 ;
      RECT 785 206145 935 206295 ;
    LAYER V2 ;
      RECT 785 212025 935 212175 ;
    LAYER V2 ;
      RECT 785 217905 935 218055 ;
    LAYER V2 ;
      RECT 785 223785 935 223935 ;
    LAYER V2 ;
      RECT 785 229665 935 229815 ;
    LAYER V2 ;
      RECT 785 235545 935 235695 ;
    LAYER V2 ;
      RECT 785 241425 935 241575 ;
    LAYER V2 ;
      RECT 785 247305 935 247455 ;
    LAYER V2 ;
      RECT 785 253185 935 253335 ;
    LAYER V2 ;
      RECT 785 259065 935 259215 ;
    LAYER V2 ;
      RECT 785 264945 935 265095 ;
    LAYER V2 ;
      RECT 785 270825 935 270975 ;
    LAYER V2 ;
      RECT 785 276705 935 276855 ;
    LAYER V2 ;
      RECT 785 282585 935 282735 ;
    LAYER V2 ;
      RECT 785 288465 935 288615 ;
    LAYER V2 ;
      RECT 785 294345 935 294495 ;
    LAYER V2 ;
      RECT 785 300225 935 300375 ;
    LAYER V2 ;
      RECT 785 306105 935 306255 ;
    LAYER V2 ;
      RECT 785 311985 935 312135 ;
    LAYER V2 ;
      RECT 785 317865 935 318015 ;
    LAYER V2 ;
      RECT 785 323745 935 323895 ;
    LAYER V2 ;
      RECT 785 329625 935 329775 ;
    LAYER V2 ;
      RECT 785 335505 935 335655 ;
    LAYER V2 ;
      RECT 785 341385 935 341535 ;
    LAYER V2 ;
      RECT 785 347265 935 347415 ;
    LAYER V2 ;
      RECT 785 353145 935 353295 ;
    LAYER V2 ;
      RECT 785 359025 935 359175 ;
    LAYER V2 ;
      RECT 785 364905 935 365055 ;
    LAYER V2 ;
      RECT 785 370785 935 370935 ;
    LAYER V2 ;
      RECT 785 376665 935 376815 ;
    LAYER V2 ;
      RECT 785 382545 935 382695 ;
    LAYER V2 ;
      RECT 785 388425 935 388575 ;
    LAYER V2 ;
      RECT 785 394305 935 394455 ;
    LAYER V2 ;
      RECT 785 400185 935 400335 ;
    LAYER V2 ;
      RECT 785 406065 935 406215 ;
    LAYER V2 ;
      RECT 785 411945 935 412095 ;
    LAYER V2 ;
      RECT 785 417825 935 417975 ;
    LAYER V2 ;
      RECT 785 423705 935 423855 ;
    LAYER V2 ;
      RECT 785 429585 935 429735 ;
    LAYER V2 ;
      RECT 785 435465 935 435615 ;
    LAYER V2 ;
      RECT 785 441345 935 441495 ;
    LAYER V2 ;
      RECT 785 447225 935 447375 ;
    LAYER V2 ;
      RECT 785 453105 935 453255 ;
    LAYER V2 ;
      RECT 785 458985 935 459135 ;
    LAYER V2 ;
      RECT 785 464865 935 465015 ;
    LAYER V2 ;
      RECT 785 470745 935 470895 ;
    LAYER V2 ;
      RECT 785 476625 935 476775 ;
    LAYER V2 ;
      RECT 785 482505 935 482655 ;
    LAYER V2 ;
      RECT 785 488385 935 488535 ;
    LAYER V2 ;
      RECT 785 494265 935 494415 ;
    LAYER V2 ;
      RECT 785 500145 935 500295 ;
    LAYER V2 ;
      RECT 785 506025 935 506175 ;
    LAYER V2 ;
      RECT 785 511905 935 512055 ;
    LAYER V2 ;
      RECT 785 517785 935 517935 ;
    LAYER V2 ;
      RECT 785 523665 935 523815 ;
    LAYER V2 ;
      RECT 785 529545 935 529695 ;
    LAYER V2 ;
      RECT 785 535425 935 535575 ;
    LAYER V2 ;
      RECT 785 541305 935 541455 ;
    LAYER V2 ;
      RECT 785 547185 935 547335 ;
    LAYER V2 ;
      RECT 785 553065 935 553215 ;
    LAYER V2 ;
      RECT 785 558945 935 559095 ;
    LAYER V2 ;
      RECT 785 564825 935 564975 ;
    LAYER V2 ;
      RECT 785 570705 935 570855 ;
    LAYER V2 ;
      RECT 785 576585 935 576735 ;
    LAYER V2 ;
      RECT 785 582465 935 582615 ;
    LAYER V2 ;
      RECT 785 588345 935 588495 ;
    LAYER V2 ;
      RECT 785 594225 935 594375 ;
    LAYER V2 ;
      RECT 785 600105 935 600255 ;
    LAYER V2 ;
      RECT 785 605985 935 606135 ;
    LAYER V2 ;
      RECT 785 611865 935 612015 ;
    LAYER V2 ;
      RECT 785 617745 935 617895 ;
    LAYER V2 ;
      RECT 785 623625 935 623775 ;
    LAYER V2 ;
      RECT 785 629505 935 629655 ;
    LAYER V2 ;
      RECT 785 635385 935 635535 ;
    LAYER V2 ;
      RECT 785 641265 935 641415 ;
    LAYER V2 ;
      RECT 785 647145 935 647295 ;
    LAYER V2 ;
      RECT 785 653025 935 653175 ;
    LAYER V2 ;
      RECT 785 658905 935 659055 ;
    LAYER V2 ;
      RECT 785 664785 935 664935 ;
    LAYER V2 ;
      RECT 785 670665 935 670815 ;
    LAYER V2 ;
      RECT 785 676545 935 676695 ;
    LAYER V2 ;
      RECT 785 682425 935 682575 ;
    LAYER V2 ;
      RECT 785 688305 935 688455 ;
    LAYER V2 ;
      RECT 785 694185 935 694335 ;
    LAYER V2 ;
      RECT 785 700065 935 700215 ;
    LAYER V2 ;
      RECT 785 705945 935 706095 ;
    LAYER V2 ;
      RECT 785 711825 935 711975 ;
    LAYER V2 ;
      RECT 785 717705 935 717855 ;
    LAYER V2 ;
      RECT 785 723585 935 723735 ;
    LAYER V2 ;
      RECT 785 729465 935 729615 ;
    LAYER V2 ;
      RECT 785 735345 935 735495 ;
    LAYER V2 ;
      RECT 785 741225 935 741375 ;
    LAYER V2 ;
      RECT 785 747105 935 747255 ;
    LAYER V2 ;
      RECT 785 752985 935 753135 ;
    LAYER V2 ;
      RECT 785 758865 935 759015 ;
    LAYER V2 ;
      RECT 785 764745 935 764895 ;
    LAYER V2 ;
      RECT 785 770625 935 770775 ;
    LAYER V2 ;
      RECT 785 776505 935 776655 ;
    LAYER V2 ;
      RECT 785 782385 935 782535 ;
    LAYER V2 ;
      RECT 785 788265 935 788415 ;
    LAYER V2 ;
      RECT 785 794145 935 794295 ;
    LAYER V2 ;
      RECT 785 800025 935 800175 ;
    LAYER V2 ;
      RECT 785 805905 935 806055 ;
    LAYER V2 ;
      RECT 785 811785 935 811935 ;
    LAYER V2 ;
      RECT 785 817665 935 817815 ;
    LAYER V2 ;
      RECT 785 823545 935 823695 ;
    LAYER V2 ;
      RECT 785 829425 935 829575 ;
    LAYER V2 ;
      RECT 785 835305 935 835455 ;
    LAYER V2 ;
      RECT 785 841185 935 841335 ;
    LAYER V2 ;
      RECT 785 847065 935 847215 ;
    LAYER V2 ;
      RECT 785 852945 935 853095 ;
    LAYER V2 ;
      RECT 785 858825 935 858975 ;
    LAYER V2 ;
      RECT 785 864705 935 864855 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1215 10425 1365 10575 ;
    LAYER V2 ;
      RECT 1215 16305 1365 16455 ;
    LAYER V2 ;
      RECT 1215 22185 1365 22335 ;
    LAYER V2 ;
      RECT 1215 28065 1365 28215 ;
    LAYER V2 ;
      RECT 1215 33945 1365 34095 ;
    LAYER V2 ;
      RECT 1215 39825 1365 39975 ;
    LAYER V2 ;
      RECT 1215 45705 1365 45855 ;
    LAYER V2 ;
      RECT 1215 51585 1365 51735 ;
    LAYER V2 ;
      RECT 1215 57465 1365 57615 ;
    LAYER V2 ;
      RECT 1215 63345 1365 63495 ;
    LAYER V2 ;
      RECT 1215 69225 1365 69375 ;
    LAYER V2 ;
      RECT 1215 75105 1365 75255 ;
    LAYER V2 ;
      RECT 1215 80985 1365 81135 ;
    LAYER V2 ;
      RECT 1215 86865 1365 87015 ;
    LAYER V2 ;
      RECT 1215 92745 1365 92895 ;
    LAYER V2 ;
      RECT 1215 98625 1365 98775 ;
    LAYER V2 ;
      RECT 1215 104505 1365 104655 ;
    LAYER V2 ;
      RECT 1215 110385 1365 110535 ;
    LAYER V2 ;
      RECT 1215 116265 1365 116415 ;
    LAYER V2 ;
      RECT 1215 122145 1365 122295 ;
    LAYER V2 ;
      RECT 1215 128025 1365 128175 ;
    LAYER V2 ;
      RECT 1215 133905 1365 134055 ;
    LAYER V2 ;
      RECT 1215 139785 1365 139935 ;
    LAYER V2 ;
      RECT 1215 145665 1365 145815 ;
    LAYER V2 ;
      RECT 1215 151545 1365 151695 ;
    LAYER V2 ;
      RECT 1215 157425 1365 157575 ;
    LAYER V2 ;
      RECT 1215 163305 1365 163455 ;
    LAYER V2 ;
      RECT 1215 169185 1365 169335 ;
    LAYER V2 ;
      RECT 1215 175065 1365 175215 ;
    LAYER V2 ;
      RECT 1215 180945 1365 181095 ;
    LAYER V2 ;
      RECT 1215 186825 1365 186975 ;
    LAYER V2 ;
      RECT 1215 192705 1365 192855 ;
    LAYER V2 ;
      RECT 1215 198585 1365 198735 ;
    LAYER V2 ;
      RECT 1215 204465 1365 204615 ;
    LAYER V2 ;
      RECT 1215 210345 1365 210495 ;
    LAYER V2 ;
      RECT 1215 216225 1365 216375 ;
    LAYER V2 ;
      RECT 1215 222105 1365 222255 ;
    LAYER V2 ;
      RECT 1215 227985 1365 228135 ;
    LAYER V2 ;
      RECT 1215 233865 1365 234015 ;
    LAYER V2 ;
      RECT 1215 239745 1365 239895 ;
    LAYER V2 ;
      RECT 1215 245625 1365 245775 ;
    LAYER V2 ;
      RECT 1215 251505 1365 251655 ;
    LAYER V2 ;
      RECT 1215 257385 1365 257535 ;
    LAYER V2 ;
      RECT 1215 263265 1365 263415 ;
    LAYER V2 ;
      RECT 1215 269145 1365 269295 ;
    LAYER V2 ;
      RECT 1215 275025 1365 275175 ;
    LAYER V2 ;
      RECT 1215 280905 1365 281055 ;
    LAYER V2 ;
      RECT 1215 286785 1365 286935 ;
    LAYER V2 ;
      RECT 1215 292665 1365 292815 ;
    LAYER V2 ;
      RECT 1215 298545 1365 298695 ;
    LAYER V2 ;
      RECT 1215 304425 1365 304575 ;
    LAYER V2 ;
      RECT 1215 310305 1365 310455 ;
    LAYER V2 ;
      RECT 1215 316185 1365 316335 ;
    LAYER V2 ;
      RECT 1215 322065 1365 322215 ;
    LAYER V2 ;
      RECT 1215 327945 1365 328095 ;
    LAYER V2 ;
      RECT 1215 333825 1365 333975 ;
    LAYER V2 ;
      RECT 1215 339705 1365 339855 ;
    LAYER V2 ;
      RECT 1215 345585 1365 345735 ;
    LAYER V2 ;
      RECT 1215 351465 1365 351615 ;
    LAYER V2 ;
      RECT 1215 357345 1365 357495 ;
    LAYER V2 ;
      RECT 1215 363225 1365 363375 ;
    LAYER V2 ;
      RECT 1215 369105 1365 369255 ;
    LAYER V2 ;
      RECT 1215 374985 1365 375135 ;
    LAYER V2 ;
      RECT 1215 380865 1365 381015 ;
    LAYER V2 ;
      RECT 1215 386745 1365 386895 ;
    LAYER V2 ;
      RECT 1215 392625 1365 392775 ;
    LAYER V2 ;
      RECT 1215 398505 1365 398655 ;
    LAYER V2 ;
      RECT 1215 404385 1365 404535 ;
    LAYER V2 ;
      RECT 1215 410265 1365 410415 ;
    LAYER V2 ;
      RECT 1215 416145 1365 416295 ;
    LAYER V2 ;
      RECT 1215 422025 1365 422175 ;
    LAYER V2 ;
      RECT 1215 427905 1365 428055 ;
    LAYER V2 ;
      RECT 1215 433785 1365 433935 ;
    LAYER V2 ;
      RECT 1215 439665 1365 439815 ;
    LAYER V2 ;
      RECT 1215 445545 1365 445695 ;
    LAYER V2 ;
      RECT 1215 451425 1365 451575 ;
    LAYER V2 ;
      RECT 1215 457305 1365 457455 ;
    LAYER V2 ;
      RECT 1215 463185 1365 463335 ;
    LAYER V2 ;
      RECT 1215 469065 1365 469215 ;
    LAYER V2 ;
      RECT 1215 474945 1365 475095 ;
    LAYER V2 ;
      RECT 1215 480825 1365 480975 ;
    LAYER V2 ;
      RECT 1215 486705 1365 486855 ;
    LAYER V2 ;
      RECT 1215 492585 1365 492735 ;
    LAYER V2 ;
      RECT 1215 498465 1365 498615 ;
    LAYER V2 ;
      RECT 1215 504345 1365 504495 ;
    LAYER V2 ;
      RECT 1215 510225 1365 510375 ;
    LAYER V2 ;
      RECT 1215 516105 1365 516255 ;
    LAYER V2 ;
      RECT 1215 521985 1365 522135 ;
    LAYER V2 ;
      RECT 1215 527865 1365 528015 ;
    LAYER V2 ;
      RECT 1215 533745 1365 533895 ;
    LAYER V2 ;
      RECT 1215 539625 1365 539775 ;
    LAYER V2 ;
      RECT 1215 545505 1365 545655 ;
    LAYER V2 ;
      RECT 1215 551385 1365 551535 ;
    LAYER V2 ;
      RECT 1215 557265 1365 557415 ;
    LAYER V2 ;
      RECT 1215 563145 1365 563295 ;
    LAYER V2 ;
      RECT 1215 569025 1365 569175 ;
    LAYER V2 ;
      RECT 1215 574905 1365 575055 ;
    LAYER V2 ;
      RECT 1215 580785 1365 580935 ;
    LAYER V2 ;
      RECT 1215 586665 1365 586815 ;
    LAYER V2 ;
      RECT 1215 592545 1365 592695 ;
    LAYER V2 ;
      RECT 1215 598425 1365 598575 ;
    LAYER V2 ;
      RECT 1215 604305 1365 604455 ;
    LAYER V2 ;
      RECT 1215 610185 1365 610335 ;
    LAYER V2 ;
      RECT 1215 616065 1365 616215 ;
    LAYER V2 ;
      RECT 1215 621945 1365 622095 ;
    LAYER V2 ;
      RECT 1215 627825 1365 627975 ;
    LAYER V2 ;
      RECT 1215 633705 1365 633855 ;
    LAYER V2 ;
      RECT 1215 639585 1365 639735 ;
    LAYER V2 ;
      RECT 1215 645465 1365 645615 ;
    LAYER V2 ;
      RECT 1215 651345 1365 651495 ;
    LAYER V2 ;
      RECT 1215 657225 1365 657375 ;
    LAYER V2 ;
      RECT 1215 663105 1365 663255 ;
    LAYER V2 ;
      RECT 1215 668985 1365 669135 ;
    LAYER V2 ;
      RECT 1215 674865 1365 675015 ;
    LAYER V2 ;
      RECT 1215 680745 1365 680895 ;
    LAYER V2 ;
      RECT 1215 686625 1365 686775 ;
    LAYER V2 ;
      RECT 1215 692505 1365 692655 ;
    LAYER V2 ;
      RECT 1215 698385 1365 698535 ;
    LAYER V2 ;
      RECT 1215 704265 1365 704415 ;
    LAYER V2 ;
      RECT 1215 710145 1365 710295 ;
    LAYER V2 ;
      RECT 1215 716025 1365 716175 ;
    LAYER V2 ;
      RECT 1215 721905 1365 722055 ;
    LAYER V2 ;
      RECT 1215 727785 1365 727935 ;
    LAYER V2 ;
      RECT 1215 733665 1365 733815 ;
    LAYER V2 ;
      RECT 1215 739545 1365 739695 ;
    LAYER V2 ;
      RECT 1215 745425 1365 745575 ;
    LAYER V2 ;
      RECT 1215 751305 1365 751455 ;
    LAYER V2 ;
      RECT 1215 757185 1365 757335 ;
    LAYER V2 ;
      RECT 1215 763065 1365 763215 ;
    LAYER V2 ;
      RECT 1215 768945 1365 769095 ;
    LAYER V2 ;
      RECT 1215 774825 1365 774975 ;
    LAYER V2 ;
      RECT 1215 780705 1365 780855 ;
    LAYER V2 ;
      RECT 1215 786585 1365 786735 ;
    LAYER V2 ;
      RECT 1215 792465 1365 792615 ;
    LAYER V2 ;
      RECT 1215 798345 1365 798495 ;
    LAYER V2 ;
      RECT 1215 804225 1365 804375 ;
    LAYER V2 ;
      RECT 1215 810105 1365 810255 ;
    LAYER V2 ;
      RECT 1215 815985 1365 816135 ;
    LAYER V2 ;
      RECT 1215 821865 1365 822015 ;
    LAYER V2 ;
      RECT 1215 827745 1365 827895 ;
    LAYER V2 ;
      RECT 1215 833625 1365 833775 ;
    LAYER V2 ;
      RECT 1215 839505 1365 839655 ;
    LAYER V2 ;
      RECT 1215 845385 1365 845535 ;
    LAYER V2 ;
      RECT 1215 851265 1365 851415 ;
    LAYER V2 ;
      RECT 1215 857145 1365 857295 ;
    LAYER V2 ;
      RECT 1215 863025 1365 863175 ;
    LAYER V2 ;
      RECT 1215 868905 1365 869055 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V2 ;
      RECT 1645 12525 1795 12675 ;
    LAYER V2 ;
      RECT 1645 18405 1795 18555 ;
    LAYER V2 ;
      RECT 1645 24285 1795 24435 ;
    LAYER V2 ;
      RECT 1645 30165 1795 30315 ;
    LAYER V2 ;
      RECT 1645 36045 1795 36195 ;
    LAYER V2 ;
      RECT 1645 41925 1795 42075 ;
    LAYER V2 ;
      RECT 1645 47805 1795 47955 ;
    LAYER V2 ;
      RECT 1645 53685 1795 53835 ;
    LAYER V2 ;
      RECT 1645 59565 1795 59715 ;
    LAYER V2 ;
      RECT 1645 65445 1795 65595 ;
    LAYER V2 ;
      RECT 1645 71325 1795 71475 ;
    LAYER V2 ;
      RECT 1645 77205 1795 77355 ;
    LAYER V2 ;
      RECT 1645 83085 1795 83235 ;
    LAYER V2 ;
      RECT 1645 88965 1795 89115 ;
    LAYER V2 ;
      RECT 1645 94845 1795 94995 ;
    LAYER V2 ;
      RECT 1645 100725 1795 100875 ;
    LAYER V2 ;
      RECT 1645 106605 1795 106755 ;
    LAYER V2 ;
      RECT 1645 112485 1795 112635 ;
    LAYER V2 ;
      RECT 1645 118365 1795 118515 ;
    LAYER V2 ;
      RECT 1645 124245 1795 124395 ;
    LAYER V2 ;
      RECT 1645 130125 1795 130275 ;
    LAYER V2 ;
      RECT 1645 136005 1795 136155 ;
    LAYER V2 ;
      RECT 1645 141885 1795 142035 ;
    LAYER V2 ;
      RECT 1645 147765 1795 147915 ;
    LAYER V2 ;
      RECT 1645 153645 1795 153795 ;
    LAYER V2 ;
      RECT 1645 159525 1795 159675 ;
    LAYER V2 ;
      RECT 1645 165405 1795 165555 ;
    LAYER V2 ;
      RECT 1645 171285 1795 171435 ;
    LAYER V2 ;
      RECT 1645 177165 1795 177315 ;
    LAYER V2 ;
      RECT 1645 183045 1795 183195 ;
    LAYER V2 ;
      RECT 1645 188925 1795 189075 ;
    LAYER V2 ;
      RECT 1645 194805 1795 194955 ;
    LAYER V2 ;
      RECT 1645 200685 1795 200835 ;
    LAYER V2 ;
      RECT 1645 206565 1795 206715 ;
    LAYER V2 ;
      RECT 1645 212445 1795 212595 ;
    LAYER V2 ;
      RECT 1645 218325 1795 218475 ;
    LAYER V2 ;
      RECT 1645 224205 1795 224355 ;
    LAYER V2 ;
      RECT 1645 230085 1795 230235 ;
    LAYER V2 ;
      RECT 1645 235965 1795 236115 ;
    LAYER V2 ;
      RECT 1645 241845 1795 241995 ;
    LAYER V2 ;
      RECT 1645 247725 1795 247875 ;
    LAYER V2 ;
      RECT 1645 253605 1795 253755 ;
    LAYER V2 ;
      RECT 1645 259485 1795 259635 ;
    LAYER V2 ;
      RECT 1645 265365 1795 265515 ;
    LAYER V2 ;
      RECT 1645 271245 1795 271395 ;
    LAYER V2 ;
      RECT 1645 277125 1795 277275 ;
    LAYER V2 ;
      RECT 1645 283005 1795 283155 ;
    LAYER V2 ;
      RECT 1645 288885 1795 289035 ;
    LAYER V2 ;
      RECT 1645 294765 1795 294915 ;
    LAYER V2 ;
      RECT 1645 300645 1795 300795 ;
    LAYER V2 ;
      RECT 1645 306525 1795 306675 ;
    LAYER V2 ;
      RECT 1645 312405 1795 312555 ;
    LAYER V2 ;
      RECT 1645 318285 1795 318435 ;
    LAYER V2 ;
      RECT 1645 324165 1795 324315 ;
    LAYER V2 ;
      RECT 1645 330045 1795 330195 ;
    LAYER V2 ;
      RECT 1645 335925 1795 336075 ;
    LAYER V2 ;
      RECT 1645 341805 1795 341955 ;
    LAYER V2 ;
      RECT 1645 347685 1795 347835 ;
    LAYER V2 ;
      RECT 1645 353565 1795 353715 ;
    LAYER V2 ;
      RECT 1645 359445 1795 359595 ;
    LAYER V2 ;
      RECT 1645 365325 1795 365475 ;
    LAYER V2 ;
      RECT 1645 371205 1795 371355 ;
    LAYER V2 ;
      RECT 1645 377085 1795 377235 ;
    LAYER V2 ;
      RECT 1645 382965 1795 383115 ;
    LAYER V2 ;
      RECT 1645 388845 1795 388995 ;
    LAYER V2 ;
      RECT 1645 394725 1795 394875 ;
    LAYER V2 ;
      RECT 1645 400605 1795 400755 ;
    LAYER V2 ;
      RECT 1645 406485 1795 406635 ;
    LAYER V2 ;
      RECT 1645 412365 1795 412515 ;
    LAYER V2 ;
      RECT 1645 418245 1795 418395 ;
    LAYER V2 ;
      RECT 1645 424125 1795 424275 ;
    LAYER V2 ;
      RECT 1645 430005 1795 430155 ;
    LAYER V2 ;
      RECT 1645 435885 1795 436035 ;
    LAYER V2 ;
      RECT 1645 441765 1795 441915 ;
    LAYER V2 ;
      RECT 1645 447645 1795 447795 ;
    LAYER V2 ;
      RECT 1645 453525 1795 453675 ;
    LAYER V2 ;
      RECT 1645 459405 1795 459555 ;
    LAYER V2 ;
      RECT 1645 465285 1795 465435 ;
    LAYER V2 ;
      RECT 1645 471165 1795 471315 ;
    LAYER V2 ;
      RECT 1645 477045 1795 477195 ;
    LAYER V2 ;
      RECT 1645 482925 1795 483075 ;
    LAYER V2 ;
      RECT 1645 488805 1795 488955 ;
    LAYER V2 ;
      RECT 1645 494685 1795 494835 ;
    LAYER V2 ;
      RECT 1645 500565 1795 500715 ;
    LAYER V2 ;
      RECT 1645 506445 1795 506595 ;
    LAYER V2 ;
      RECT 1645 512325 1795 512475 ;
    LAYER V2 ;
      RECT 1645 518205 1795 518355 ;
    LAYER V2 ;
      RECT 1645 524085 1795 524235 ;
    LAYER V2 ;
      RECT 1645 529965 1795 530115 ;
    LAYER V2 ;
      RECT 1645 535845 1795 535995 ;
    LAYER V2 ;
      RECT 1645 541725 1795 541875 ;
    LAYER V2 ;
      RECT 1645 547605 1795 547755 ;
    LAYER V2 ;
      RECT 1645 553485 1795 553635 ;
    LAYER V2 ;
      RECT 1645 559365 1795 559515 ;
    LAYER V2 ;
      RECT 1645 565245 1795 565395 ;
    LAYER V2 ;
      RECT 1645 571125 1795 571275 ;
    LAYER V2 ;
      RECT 1645 577005 1795 577155 ;
    LAYER V2 ;
      RECT 1645 582885 1795 583035 ;
    LAYER V2 ;
      RECT 1645 588765 1795 588915 ;
    LAYER V2 ;
      RECT 1645 594645 1795 594795 ;
    LAYER V2 ;
      RECT 1645 600525 1795 600675 ;
    LAYER V2 ;
      RECT 1645 606405 1795 606555 ;
    LAYER V2 ;
      RECT 1645 612285 1795 612435 ;
    LAYER V2 ;
      RECT 1645 618165 1795 618315 ;
    LAYER V2 ;
      RECT 1645 624045 1795 624195 ;
    LAYER V2 ;
      RECT 1645 629925 1795 630075 ;
    LAYER V2 ;
      RECT 1645 635805 1795 635955 ;
    LAYER V2 ;
      RECT 1645 641685 1795 641835 ;
    LAYER V2 ;
      RECT 1645 647565 1795 647715 ;
    LAYER V2 ;
      RECT 1645 653445 1795 653595 ;
    LAYER V2 ;
      RECT 1645 659325 1795 659475 ;
    LAYER V2 ;
      RECT 1645 665205 1795 665355 ;
    LAYER V2 ;
      RECT 1645 671085 1795 671235 ;
    LAYER V2 ;
      RECT 1645 676965 1795 677115 ;
    LAYER V2 ;
      RECT 1645 682845 1795 682995 ;
    LAYER V2 ;
      RECT 1645 688725 1795 688875 ;
    LAYER V2 ;
      RECT 1645 694605 1795 694755 ;
    LAYER V2 ;
      RECT 1645 700485 1795 700635 ;
    LAYER V2 ;
      RECT 1645 706365 1795 706515 ;
    LAYER V2 ;
      RECT 1645 712245 1795 712395 ;
    LAYER V2 ;
      RECT 1645 718125 1795 718275 ;
    LAYER V2 ;
      RECT 1645 724005 1795 724155 ;
    LAYER V2 ;
      RECT 1645 729885 1795 730035 ;
    LAYER V2 ;
      RECT 1645 735765 1795 735915 ;
    LAYER V2 ;
      RECT 1645 741645 1795 741795 ;
    LAYER V2 ;
      RECT 1645 747525 1795 747675 ;
    LAYER V2 ;
      RECT 1645 753405 1795 753555 ;
    LAYER V2 ;
      RECT 1645 759285 1795 759435 ;
    LAYER V2 ;
      RECT 1645 765165 1795 765315 ;
    LAYER V2 ;
      RECT 1645 771045 1795 771195 ;
    LAYER V2 ;
      RECT 1645 776925 1795 777075 ;
    LAYER V2 ;
      RECT 1645 782805 1795 782955 ;
    LAYER V2 ;
      RECT 1645 788685 1795 788835 ;
    LAYER V2 ;
      RECT 1645 794565 1795 794715 ;
    LAYER V2 ;
      RECT 1645 800445 1795 800595 ;
    LAYER V2 ;
      RECT 1645 806325 1795 806475 ;
    LAYER V2 ;
      RECT 1645 812205 1795 812355 ;
    LAYER V2 ;
      RECT 1645 818085 1795 818235 ;
    LAYER V2 ;
      RECT 1645 823965 1795 824115 ;
    LAYER V2 ;
      RECT 1645 829845 1795 829995 ;
    LAYER V2 ;
      RECT 1645 835725 1795 835875 ;
    LAYER V2 ;
      RECT 1645 841605 1795 841755 ;
    LAYER V2 ;
      RECT 1645 847485 1795 847635 ;
    LAYER V2 ;
      RECT 1645 853365 1795 853515 ;
    LAYER V2 ;
      RECT 1645 859245 1795 859395 ;
    LAYER V2 ;
      RECT 1645 865125 1795 865275 ;
    LAYER V2 ;
      RECT 1645 871005 1795 871155 ;
  END
END NMOS_S_12565100_X1_Y148
