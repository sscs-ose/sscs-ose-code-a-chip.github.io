# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.41000 BY  11.69000 ;
  OBS
    LAYER li1 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.330000  0.140000 11.220000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.280000  0.470000  0.420000 11.360000 ;
      RECT  0.560000  0.330000  0.700000 11.220000 ;
      RECT  0.840000  0.470000  0.980000 11.360000 ;
      RECT  1.120000  0.330000  1.260000 11.220000 ;
      RECT  1.400000  0.470000  1.540000 11.360000 ;
      RECT  1.680000  0.330000  1.820000 11.220000 ;
      RECT  1.960000  0.470000  2.100000 11.360000 ;
      RECT  2.240000  0.330000  2.380000 11.220000 ;
      RECT  2.520000  0.470000  2.660000 11.360000 ;
      RECT  2.800000  0.330000  2.940000 11.220000 ;
      RECT  3.080000  0.470000  3.220000 11.360000 ;
      RECT  3.360000  0.330000  3.500000 11.220000 ;
      RECT  3.640000  0.470000  3.780000 11.360000 ;
      RECT  3.920000  0.330000  4.060000 11.220000 ;
      RECT  4.200000  0.470000  4.340000 11.360000 ;
      RECT  4.480000  0.330000  4.620000 11.220000 ;
      RECT  4.760000  0.470000  4.900000 11.360000 ;
      RECT  5.040000  0.330000  5.180000 11.220000 ;
      RECT  5.320000  0.470000  5.460000 11.360000 ;
      RECT  5.600000  0.330000  5.740000 11.220000 ;
      RECT  5.880000  0.470000  6.020000 11.360000 ;
      RECT  6.160000  0.330000  6.300000 11.220000 ;
      RECT  6.440000  0.470000  6.580000 11.360000 ;
      RECT  6.720000  0.330000  6.860000 11.220000 ;
      RECT  7.000000  0.470000  7.140000 11.360000 ;
      RECT  7.280000  0.330000  7.420000 11.220000 ;
      RECT  7.560000  0.470000  7.700000 11.360000 ;
      RECT  7.840000  0.330000  7.980000 11.220000 ;
      RECT  8.120000  0.470000  8.260000 11.360000 ;
      RECT  8.400000  0.330000  8.540000 11.220000 ;
      RECT  8.680000  0.470000  8.820000 11.360000 ;
      RECT  8.960000  0.330000  9.100000 11.220000 ;
      RECT  9.240000  0.470000  9.380000 11.360000 ;
      RECT  9.520000  0.330000  9.660000 11.220000 ;
      RECT  9.800000  0.470000  9.940000 11.360000 ;
      RECT 10.080000  0.330000 10.220000 11.220000 ;
      RECT 10.360000  0.470000 10.500000 11.360000 ;
      RECT 10.640000  0.330000 10.780000 11.220000 ;
      RECT 10.920000  0.470000 11.060000 11.360000 ;
      RECT 11.200000  0.330000 11.410000 11.220000 ;
    LAYER mcon ;
      RECT  0.190000  0.080000  0.360000  0.250000 ;
      RECT  0.190000 11.440000  0.360000 11.610000 ;
      RECT  0.550000  0.080000  0.720000  0.250000 ;
      RECT  0.550000 11.440000  0.720000 11.610000 ;
      RECT  0.910000  0.080000  1.080000  0.250000 ;
      RECT  0.910000 11.440000  1.080000 11.610000 ;
      RECT  1.270000  0.080000  1.440000  0.250000 ;
      RECT  1.270000 11.440000  1.440000 11.610000 ;
      RECT  1.630000  0.080000  1.800000  0.250000 ;
      RECT  1.630000 11.440000  1.800000 11.610000 ;
      RECT  1.990000  0.080000  2.160000  0.250000 ;
      RECT  1.990000 11.440000  2.160000 11.610000 ;
      RECT  2.350000  0.080000  2.520000  0.250000 ;
      RECT  2.350000 11.440000  2.520000 11.610000 ;
      RECT  2.710000  0.080000  2.880000  0.250000 ;
      RECT  2.710000 11.440000  2.880000 11.610000 ;
      RECT  3.070000  0.080000  3.240000  0.250000 ;
      RECT  3.070000 11.440000  3.240000 11.610000 ;
      RECT  3.430000  0.080000  3.600000  0.250000 ;
      RECT  3.430000 11.440000  3.600000 11.610000 ;
      RECT  3.790000  0.080000  3.960000  0.250000 ;
      RECT  3.790000 11.440000  3.960000 11.610000 ;
      RECT  4.150000  0.080000  4.320000  0.250000 ;
      RECT  4.150000 11.440000  4.320000 11.610000 ;
      RECT  4.510000  0.080000  4.680000  0.250000 ;
      RECT  4.510000 11.440000  4.680000 11.610000 ;
      RECT  4.870000  0.080000  5.040000  0.250000 ;
      RECT  4.870000 11.440000  5.040000 11.610000 ;
      RECT  5.230000  0.080000  5.400000  0.250000 ;
      RECT  5.230000 11.440000  5.400000 11.610000 ;
      RECT  5.590000  0.080000  5.760000  0.250000 ;
      RECT  5.590000 11.440000  5.760000 11.610000 ;
      RECT  5.950000  0.080000  6.120000  0.250000 ;
      RECT  5.950000 11.440000  6.120000 11.610000 ;
      RECT  6.310000  0.080000  6.480000  0.250000 ;
      RECT  6.310000 11.440000  6.480000 11.610000 ;
      RECT  6.670000  0.080000  6.840000  0.250000 ;
      RECT  6.670000 11.440000  6.840000 11.610000 ;
      RECT  7.030000  0.080000  7.200000  0.250000 ;
      RECT  7.030000 11.440000  7.200000 11.610000 ;
      RECT  7.390000  0.080000  7.560000  0.250000 ;
      RECT  7.390000 11.440000  7.560000 11.610000 ;
      RECT  7.750000  0.080000  7.920000  0.250000 ;
      RECT  7.750000 11.440000  7.920000 11.610000 ;
      RECT  8.110000  0.080000  8.280000  0.250000 ;
      RECT  8.110000 11.440000  8.280000 11.610000 ;
      RECT  8.470000  0.080000  8.640000  0.250000 ;
      RECT  8.470000 11.440000  8.640000 11.610000 ;
      RECT  8.830000  0.080000  9.000000  0.250000 ;
      RECT  8.830000 11.440000  9.000000 11.610000 ;
      RECT  9.190000  0.080000  9.360000  0.250000 ;
      RECT  9.190000 11.440000  9.360000 11.610000 ;
      RECT  9.550000  0.080000  9.720000  0.250000 ;
      RECT  9.550000 11.440000  9.720000 11.610000 ;
      RECT  9.910000  0.080000 10.080000  0.250000 ;
      RECT  9.910000 11.440000 10.080000 11.610000 ;
      RECT 10.270000  0.080000 10.440000  0.250000 ;
      RECT 10.270000 11.440000 10.440000 11.610000 ;
      RECT 10.630000  0.080000 10.800000  0.250000 ;
      RECT 10.630000 11.440000 10.800000 11.610000 ;
      RECT 10.990000  0.080000 11.160000  0.250000 ;
      RECT 10.990000 11.440000 11.160000 11.610000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.470000  0.140000 11.360000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.280000  0.330000  0.420000 11.220000 ;
      RECT  0.560000  0.470000  0.700000 11.360000 ;
      RECT  0.840000  0.330000  0.980000 11.220000 ;
      RECT  1.120000  0.470000  1.260000 11.360000 ;
      RECT  1.400000  0.330000  1.540000 11.220000 ;
      RECT  1.680000  0.470000  1.820000 11.360000 ;
      RECT  1.960000  0.330000  2.100000 11.220000 ;
      RECT  2.240000  0.470000  2.380000 11.360000 ;
      RECT  2.520000  0.330000  2.660000 11.220000 ;
      RECT  2.800000  0.470000  2.940000 11.360000 ;
      RECT  3.080000  0.330000  3.220000 11.220000 ;
      RECT  3.360000  0.470000  3.500000 11.360000 ;
      RECT  3.640000  0.330000  3.780000 11.220000 ;
      RECT  3.920000  0.470000  4.060000 11.360000 ;
      RECT  4.200000  0.330000  4.340000 11.220000 ;
      RECT  4.480000  0.470000  4.620000 11.360000 ;
      RECT  4.760000  0.330000  4.900000 11.220000 ;
      RECT  5.040000  0.470000  5.180000 11.360000 ;
      RECT  5.320000  0.330000  5.460000 11.220000 ;
      RECT  5.600000  0.470000  5.740000 11.360000 ;
      RECT  5.880000  0.330000  6.020000 11.220000 ;
      RECT  6.160000  0.470000  6.300000 11.360000 ;
      RECT  6.440000  0.330000  6.580000 11.220000 ;
      RECT  6.720000  0.470000  6.860000 11.360000 ;
      RECT  7.000000  0.330000  7.140000 11.220000 ;
      RECT  7.280000  0.470000  7.420000 11.360000 ;
      RECT  7.560000  0.330000  7.700000 11.220000 ;
      RECT  7.840000  0.470000  7.980000 11.360000 ;
      RECT  8.120000  0.330000  8.260000 11.220000 ;
      RECT  8.400000  0.470000  8.540000 11.360000 ;
      RECT  8.680000  0.330000  8.820000 11.220000 ;
      RECT  8.960000  0.470000  9.100000 11.360000 ;
      RECT  9.240000  0.330000  9.380000 11.220000 ;
      RECT  9.520000  0.470000  9.660000 11.360000 ;
      RECT  9.800000  0.330000  9.940000 11.220000 ;
      RECT 10.080000  0.470000 10.220000 11.360000 ;
      RECT 10.360000  0.330000 10.500000 11.220000 ;
      RECT 10.640000  0.470000 10.780000 11.360000 ;
      RECT 10.920000  0.330000 11.060000 11.220000 ;
      RECT 11.200000  0.470000 11.410000 11.360000 ;
    LAYER met2 ;
      RECT  0.000000  0.000000  0.700000  0.330000 ;
      RECT  0.000000  0.330000  0.140000 11.690000 ;
      RECT  0.280000  0.470000  0.420000 11.360000 ;
      RECT  0.280000 11.360000  0.980000 11.690000 ;
      RECT  0.560000  0.330000  0.700000 11.220000 ;
      RECT  0.840000  0.000000  0.980000 11.360000 ;
      RECT  1.120000  0.000000  1.820000  0.330000 ;
      RECT  1.120000  0.330000  1.260000 11.690000 ;
      RECT  1.400000  0.470000  1.540000 11.360000 ;
      RECT  1.400000 11.360000  2.100000 11.690000 ;
      RECT  1.680000  0.330000  1.820000 11.220000 ;
      RECT  1.960000  0.000000  2.100000 11.360000 ;
      RECT  2.240000  0.000000  2.940000  0.330000 ;
      RECT  2.240000  0.330000  2.380000 11.690000 ;
      RECT  2.520000  0.470000  2.660000 11.360000 ;
      RECT  2.520000 11.360000  3.220000 11.690000 ;
      RECT  2.800000  0.330000  2.940000 11.220000 ;
      RECT  3.080000  0.000000  3.220000 11.360000 ;
      RECT  3.360000  0.000000  4.060000  0.330000 ;
      RECT  3.360000  0.330000  3.500000 11.690000 ;
      RECT  3.640000  0.470000  3.780000 11.360000 ;
      RECT  3.640000 11.360000  4.340000 11.690000 ;
      RECT  3.920000  0.330000  4.060000 11.220000 ;
      RECT  4.200000  0.000000  4.340000 11.360000 ;
      RECT  4.480000  0.000000  5.180000  0.330000 ;
      RECT  4.480000  0.330000  4.620000 11.690000 ;
      RECT  4.760000  0.470000  4.900000 11.360000 ;
      RECT  4.760000 11.360000  5.460000 11.690000 ;
      RECT  5.040000  0.330000  5.180000 11.220000 ;
      RECT  5.320000  0.000000  5.460000 11.360000 ;
      RECT  5.600000  0.000000  6.300000  0.330000 ;
      RECT  5.600000  0.330000  5.740000 11.690000 ;
      RECT  5.880000  0.470000  6.020000 11.360000 ;
      RECT  5.880000 11.360000  6.580000 11.690000 ;
      RECT  6.160000  0.330000  6.300000 11.220000 ;
      RECT  6.440000  0.000000  6.580000 11.360000 ;
      RECT  6.720000  0.000000  7.420000  0.330000 ;
      RECT  6.720000  0.330000  6.860000 11.690000 ;
      RECT  7.000000  0.470000  7.140000 11.360000 ;
      RECT  7.000000 11.360000  7.700000 11.690000 ;
      RECT  7.280000  0.330000  7.420000 11.220000 ;
      RECT  7.560000  0.000000  7.700000 11.360000 ;
      RECT  7.840000  0.000000  8.540000  0.330000 ;
      RECT  7.840000  0.330000  7.980000 11.690000 ;
      RECT  8.120000  0.470000  8.260000 11.360000 ;
      RECT  8.120000 11.360000  8.820000 11.690000 ;
      RECT  8.400000  0.330000  8.540000 11.220000 ;
      RECT  8.680000  0.000000  8.820000 11.360000 ;
      RECT  8.960000  0.000000  9.660000  0.330000 ;
      RECT  8.960000  0.330000  9.100000 11.690000 ;
      RECT  9.240000  0.470000  9.380000 11.360000 ;
      RECT  9.240000 11.360000 11.410000 11.690000 ;
      RECT  9.520000  0.330000  9.660000 11.220000 ;
      RECT  9.800000  0.000000  9.940000 11.360000 ;
      RECT 10.080000  0.000000 11.410000  0.330000 ;
      RECT 10.080000  0.330000 10.220000 11.220000 ;
      RECT 10.360000  0.470000 10.500000 11.360000 ;
      RECT 10.640000  0.330000 10.780000 11.220000 ;
      RECT 10.920000  0.470000 11.060000 11.360000 ;
      RECT 11.200000  0.330000 11.410000 11.220000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.630000  0.300000 11.360000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.600000  0.330000  0.900000 11.060000 ;
      RECT  1.200000  0.630000  1.500000 11.360000 ;
      RECT  1.800000  0.330000  2.100000 11.060000 ;
      RECT  2.400000  0.630000  2.700000 11.360000 ;
      RECT  3.000000  0.330000  3.300000 11.060000 ;
      RECT  3.600000  0.630000  3.900000 11.360000 ;
      RECT  4.200000  0.330000  4.500000 11.060000 ;
      RECT  4.800000  0.630000  5.100000 11.360000 ;
      RECT  5.400000  0.330000  5.700000 11.060000 ;
      RECT  6.000000  0.630000  6.300000 11.360000 ;
      RECT  6.600000  0.330000  6.900000 11.060000 ;
      RECT  7.200000  0.630000  7.500000 11.360000 ;
      RECT  7.800000  0.330000  8.100000 11.060000 ;
      RECT  8.400000  0.630000  8.700000 11.360000 ;
      RECT  9.000000  0.330000  9.300000 11.060000 ;
      RECT  9.600000  0.630000  9.900000 11.360000 ;
      RECT 10.200000  0.330000 10.500000 11.060000 ;
      RECT 10.800000  0.630000 11.410000 11.360000 ;
    LAYER met4 ;
      RECT  0.000000  0.000000 11.410000  0.330000 ;
      RECT  0.000000  0.330000  0.300000 11.060000 ;
      RECT  0.000000 11.360000 11.410000 11.690000 ;
      RECT  0.600000  0.630000  0.900000 10.135000 ;
      RECT  0.600000 10.135000  2.100000 11.360000 ;
      RECT  1.200000  0.330000  2.700000  1.555000 ;
      RECT  1.200000  1.555000  1.500000  9.835000 ;
      RECT  1.800000  1.855000  2.100000 10.135000 ;
      RECT  2.400000  1.555000  2.700000 11.060000 ;
      RECT  3.000000  0.630000  3.300000 11.360000 ;
      RECT  3.600000  0.330000  3.900000 11.060000 ;
      RECT  4.200000  0.630000  4.500000 11.360000 ;
      RECT  4.800000  0.330000  5.100000 11.060000 ;
      RECT  5.400000  0.630000  5.700000 11.360000 ;
      RECT  6.000000  0.330000  6.300000 11.060000 ;
      RECT  6.600000  0.630000  6.900000 11.360000 ;
      RECT  7.200000  0.330000  7.500000 11.060000 ;
      RECT  7.800000  0.630000  8.100000 10.135000 ;
      RECT  7.800000 10.135000  9.300000 11.360000 ;
      RECT  8.400000  0.330000  9.900000  1.555000 ;
      RECT  8.400000  1.555000  8.700000  9.835000 ;
      RECT  9.000000  1.855000  9.300000 10.135000 ;
      RECT  9.600000  1.555000  9.900000 11.060000 ;
      RECT 10.200000  0.630000 10.500000 11.360000 ;
      RECT 10.800000  0.330000 11.410000 11.060000 ;
    LAYER met5 ;
      RECT 0.000000  0.000000 11.410000  1.675000 ;
      RECT 0.000000  3.275000  1.600000 10.015000 ;
      RECT 0.000000 10.015000 11.410000 11.690000 ;
      RECT 3.200000  1.675000  4.800000  8.415000 ;
      RECT 6.400000  3.275000  8.000000 10.015000 ;
      RECT 9.600000  1.675000 11.410000  8.415000 ;
    LAYER via ;
      RECT  0.120000  0.035000  0.380000  0.295000 ;
      RECT  0.340000 11.395000  0.600000 11.655000 ;
      RECT  0.440000  0.035000  0.700000  0.295000 ;
      RECT  0.660000 11.395000  0.920000 11.655000 ;
      RECT  1.180000  0.035000  1.440000  0.295000 ;
      RECT  1.460000 11.395000  1.720000 11.655000 ;
      RECT  1.500000  0.035000  1.760000  0.295000 ;
      RECT  1.780000 11.395000  2.040000 11.655000 ;
      RECT  2.300000  0.035000  2.560000  0.295000 ;
      RECT  2.580000 11.395000  2.840000 11.655000 ;
      RECT  2.620000  0.035000  2.880000  0.295000 ;
      RECT  2.900000 11.395000  3.160000 11.655000 ;
      RECT  3.420000  0.035000  3.680000  0.295000 ;
      RECT  3.700000 11.395000  3.960000 11.655000 ;
      RECT  3.740000  0.035000  4.000000  0.295000 ;
      RECT  4.020000 11.395000  4.280000 11.655000 ;
      RECT  4.540000  0.035000  4.800000  0.295000 ;
      RECT  4.820000 11.395000  5.080000 11.655000 ;
      RECT  4.860000  0.035000  5.120000  0.295000 ;
      RECT  5.140000 11.395000  5.400000 11.655000 ;
      RECT  5.660000  0.035000  5.920000  0.295000 ;
      RECT  5.940000 11.395000  6.200000 11.655000 ;
      RECT  5.980000  0.035000  6.240000  0.295000 ;
      RECT  6.260000 11.395000  6.520000 11.655000 ;
      RECT  6.780000  0.035000  7.040000  0.295000 ;
      RECT  7.060000 11.395000  7.320000 11.655000 ;
      RECT  7.100000  0.035000  7.360000  0.295000 ;
      RECT  7.380000 11.395000  7.640000 11.655000 ;
      RECT  7.900000  0.035000  8.160000  0.295000 ;
      RECT  8.180000 11.395000  8.440000 11.655000 ;
      RECT  8.220000  0.035000  8.480000  0.295000 ;
      RECT  8.500000 11.395000  8.760000 11.655000 ;
      RECT  9.020000  0.035000  9.280000  0.295000 ;
      RECT  9.300000 11.395000  9.560000 11.655000 ;
      RECT  9.340000  0.035000  9.600000  0.295000 ;
      RECT  9.620000 11.395000  9.880000 11.655000 ;
      RECT 10.140000  0.035000 10.400000  0.295000 ;
      RECT 10.420000 11.395000 10.680000 11.655000 ;
      RECT 10.460000  0.035000 10.720000  0.295000 ;
      RECT 10.740000 11.395000 11.000000 11.655000 ;
    LAYER via2 ;
      RECT  0.210000  0.025000  0.490000  0.305000 ;
      RECT  0.490000 11.385000  0.770000 11.665000 ;
      RECT  1.330000  0.025000  1.610000  0.305000 ;
      RECT  1.610000 11.385000  1.890000 11.665000 ;
      RECT  2.450000  0.025000  2.730000  0.305000 ;
      RECT  2.730000 11.385000  3.010000 11.665000 ;
      RECT  3.570000  0.025000  3.850000  0.305000 ;
      RECT  3.850000 11.385000  4.130000 11.665000 ;
      RECT  4.690000  0.025000  4.970000  0.305000 ;
      RECT  4.970000 11.385000  5.250000 11.665000 ;
      RECT  5.810000  0.025000  6.090000  0.305000 ;
      RECT  6.090000 11.385000  6.370000 11.665000 ;
      RECT  6.930000  0.025000  7.210000  0.305000 ;
      RECT  7.210000 11.385000  7.490000 11.665000 ;
      RECT  8.050000  0.025000  8.330000  0.305000 ;
      RECT  8.330000 11.385000  8.610000 11.665000 ;
      RECT  9.170000  0.025000  9.450000  0.305000 ;
      RECT  9.450000 11.385000  9.730000 11.665000 ;
      RECT 10.290000  0.025000 10.570000  0.305000 ;
      RECT 10.570000 11.385000 10.850000 11.665000 ;
    LAYER via3 ;
      RECT  0.140000  0.005000  0.460000  0.325000 ;
      RECT  0.140000 11.365000  0.460000 11.685000 ;
      RECT  0.540000  0.005000  0.860000  0.325000 ;
      RECT  0.540000 11.365000  0.860000 11.685000 ;
      RECT  0.940000  0.005000  1.260000  0.325000 ;
      RECT  0.940000 11.365000  1.260000 11.685000 ;
      RECT  1.340000  0.005000  1.660000  0.325000 ;
      RECT  1.340000 11.365000  1.660000 11.685000 ;
      RECT  1.740000  0.005000  2.060000  0.325000 ;
      RECT  1.740000 11.365000  2.060000 11.685000 ;
      RECT  2.140000  0.005000  2.460000  0.325000 ;
      RECT  2.140000 11.365000  2.460000 11.685000 ;
      RECT  2.540000  0.005000  2.860000  0.325000 ;
      RECT  2.540000 11.365000  2.860000 11.685000 ;
      RECT  2.940000  0.005000  3.260000  0.325000 ;
      RECT  2.940000 11.365000  3.260000 11.685000 ;
      RECT  3.340000  0.005000  3.660000  0.325000 ;
      RECT  3.340000 11.365000  3.660000 11.685000 ;
      RECT  3.740000  0.005000  4.060000  0.325000 ;
      RECT  3.740000 11.365000  4.060000 11.685000 ;
      RECT  4.140000  0.005000  4.460000  0.325000 ;
      RECT  4.140000 11.365000  4.460000 11.685000 ;
      RECT  4.540000  0.005000  4.860000  0.325000 ;
      RECT  4.540000 11.365000  4.860000 11.685000 ;
      RECT  4.940000  0.005000  5.260000  0.325000 ;
      RECT  4.940000 11.365000  5.260000 11.685000 ;
      RECT  5.340000  0.005000  5.660000  0.325000 ;
      RECT  5.340000 11.365000  5.660000 11.685000 ;
      RECT  5.740000  0.005000  6.060000  0.325000 ;
      RECT  5.740000 11.365000  6.060000 11.685000 ;
      RECT  6.140000  0.005000  6.460000  0.325000 ;
      RECT  6.140000 11.365000  6.460000 11.685000 ;
      RECT  6.540000  0.005000  6.860000  0.325000 ;
      RECT  6.540000 11.365000  6.860000 11.685000 ;
      RECT  6.940000  0.005000  7.260000  0.325000 ;
      RECT  6.940000 11.365000  7.260000 11.685000 ;
      RECT  7.340000  0.005000  7.660000  0.325000 ;
      RECT  7.340000 11.365000  7.660000 11.685000 ;
      RECT  7.740000  0.005000  8.060000  0.325000 ;
      RECT  7.740000 11.365000  8.060000 11.685000 ;
      RECT  8.140000  0.005000  8.460000  0.325000 ;
      RECT  8.140000 11.365000  8.460000 11.685000 ;
      RECT  8.540000  0.005000  8.860000  0.325000 ;
      RECT  8.540000 11.365000  8.860000 11.685000 ;
      RECT  8.940000  0.005000  9.260000  0.325000 ;
      RECT  8.940000 11.365000  9.260000 11.685000 ;
      RECT  9.340000  0.005000  9.660000  0.325000 ;
      RECT  9.340000 11.365000  9.660000 11.685000 ;
      RECT  9.740000  0.005000 10.060000  0.325000 ;
      RECT  9.740000 11.365000 10.060000 11.685000 ;
      RECT 10.140000  0.005000 10.460000  0.325000 ;
      RECT 10.140000 11.365000 10.460000 11.685000 ;
      RECT 10.540000  0.005000 10.860000  0.325000 ;
      RECT 10.540000 11.365000 10.860000 11.685000 ;
      RECT 10.940000  0.005000 11.260000  0.325000 ;
      RECT 10.940000 11.365000 11.260000 11.685000 ;
    LAYER via4 ;
      RECT 0.760000 10.135000 1.940000 11.315000 ;
      RECT 1.360000  0.375000 2.540000  1.555000 ;
      RECT 7.960000 10.135000 9.140000 11.315000 ;
      RECT 8.560000  0.375000 9.740000  1.555000 ;
  END
END sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield
END LIBRARY
