# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.900000 BY  5.900000 ;
  PIN C0
    PORT
      LAYER met4 ;
        RECT 0.000000 0.000000 5.900000 0.330000 ;
        RECT 0.000000 0.330000 0.330000 1.230000 ;
        RECT 0.000000 1.230000 5.130000 1.530000 ;
        RECT 0.000000 1.530000 0.330000 2.430000 ;
        RECT 0.000000 2.430000 5.130000 2.730000 ;
        RECT 0.000000 2.730000 0.330000 3.630000 ;
        RECT 0.000000 3.630000 5.130000 3.930000 ;
        RECT 0.000000 3.930000 0.330000 4.830000 ;
        RECT 0.000000 4.830000 5.130000 5.130000 ;
        RECT 0.000000 5.130000 0.330000 5.900000 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met4 ;
        RECT 0.630000 0.630000 5.900000 0.930000 ;
        RECT 0.630000 1.830000 5.900000 2.130000 ;
        RECT 0.630000 3.030000 5.900000 3.330000 ;
        RECT 0.630000 4.230000 5.900000 4.530000 ;
        RECT 0.630000 5.430000 5.900000 5.900000 ;
        RECT 5.430000 0.930000 5.900000 1.830000 ;
        RECT 5.430000 2.130000 5.900000 3.030000 ;
        RECT 5.430000 3.330000 5.900000 4.230000 ;
        RECT 5.430000 4.530000 5.900000 5.430000 ;
    END
  END C1
  PIN SUB
    PORT
      LAYER pwell ;
        RECT 2.615000 4.085000 2.720000 4.330000 ;
    END
  END SUB
  OBS
    LAYER li1 ;
      RECT 0.080000 0.080000 5.750000 0.250000 ;
      RECT 0.080000 0.250000 0.250000 5.580000 ;
      RECT 0.080000 5.580000 5.750000 5.750000 ;
      RECT 5.580000 0.250000 5.750000 5.580000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 5.820000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 5.820000 ;
      RECT 0.470000 0.470000 0.610000 5.510000 ;
      RECT 0.470000 5.510000 5.820000 5.820000 ;
      RECT 0.750000 0.330000 0.890000 5.370000 ;
      RECT 1.030000 0.470000 1.170000 5.510000 ;
      RECT 1.310000 0.330000 1.450000 5.370000 ;
      RECT 1.590000 0.470000 1.730000 5.510000 ;
      RECT 1.870000 0.330000 2.010000 5.370000 ;
      RECT 2.150000 0.470000 2.290000 5.510000 ;
      RECT 2.430000 0.330000 2.570000 5.370000 ;
      RECT 2.710000 0.470000 2.850000 5.510000 ;
      RECT 2.990000 0.330000 3.130000 5.370000 ;
      RECT 3.270000 0.470000 3.410000 5.510000 ;
      RECT 3.550000 0.330000 3.690000 5.370000 ;
      RECT 3.830000 0.470000 3.970000 5.510000 ;
      RECT 4.110000 0.330000 4.250000 5.370000 ;
      RECT 4.390000 0.470000 4.530000 5.510000 ;
      RECT 4.670000 0.330000 4.810000 5.370000 ;
      RECT 4.950000 0.470000 5.090000 5.510000 ;
      RECT 5.230000 0.330000 5.370000 5.370000 ;
      RECT 5.510000 0.470000 5.820000 5.510000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 5.370000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 0.750000 ;
      RECT 0.000000 0.750000 5.370000 0.890000 ;
      RECT 0.000000 0.890000 0.330000 1.310000 ;
      RECT 0.000000 1.310000 5.370000 1.450000 ;
      RECT 0.000000 1.450000 0.330000 1.870000 ;
      RECT 0.000000 1.870000 5.370000 2.010000 ;
      RECT 0.000000 2.010000 0.330000 2.430000 ;
      RECT 0.000000 2.430000 5.370000 2.570000 ;
      RECT 0.000000 2.570000 0.330000 2.990000 ;
      RECT 0.000000 2.990000 5.370000 3.130000 ;
      RECT 0.000000 3.130000 0.330000 3.550000 ;
      RECT 0.000000 3.550000 5.370000 3.690000 ;
      RECT 0.000000 3.690000 0.330000 4.110000 ;
      RECT 0.000000 4.110000 5.370000 4.250000 ;
      RECT 0.000000 4.250000 0.330000 4.670000 ;
      RECT 0.000000 4.670000 5.370000 4.810000 ;
      RECT 0.000000 4.810000 0.330000 5.230000 ;
      RECT 0.000000 5.230000 5.370000 5.370000 ;
      RECT 0.330000 5.510000 5.820000 5.820000 ;
      RECT 0.470000 0.470000 5.820000 0.610000 ;
      RECT 0.470000 1.030000 5.820000 1.170000 ;
      RECT 0.470000 1.590000 5.820000 1.730000 ;
      RECT 0.470000 2.150000 5.820000 2.290000 ;
      RECT 0.470000 2.710000 5.820000 2.850000 ;
      RECT 0.470000 3.270000 5.820000 3.410000 ;
      RECT 0.470000 3.830000 5.820000 3.970000 ;
      RECT 0.470000 4.390000 5.820000 4.530000 ;
      RECT 0.470000 4.950000 5.820000 5.090000 ;
      RECT 5.510000 0.330000 5.820000 0.470000 ;
      RECT 5.510000 0.610000 5.820000 1.030000 ;
      RECT 5.510000 1.170000 5.820000 1.590000 ;
      RECT 5.510000 1.730000 5.820000 2.150000 ;
      RECT 5.510000 2.290000 5.820000 2.710000 ;
      RECT 5.510000 2.850000 5.820000 3.270000 ;
      RECT 5.510000 3.410000 5.820000 3.830000 ;
      RECT 5.510000 3.970000 5.820000 4.390000 ;
      RECT 5.510000 4.530000 5.820000 4.950000 ;
      RECT 5.510000 5.090000 5.820000 5.510000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 5.130000 0.330000 ;
      RECT 0.000000 0.330000 0.330000 5.130000 ;
      RECT 0.330000 5.430000 5.900000 5.900000 ;
      RECT 0.630000 0.630000 0.930000 5.430000 ;
      RECT 1.230000 0.330000 1.530000 5.130000 ;
      RECT 1.830000 0.630000 2.130000 5.430000 ;
      RECT 2.430000 0.330000 2.730000 5.130000 ;
      RECT 3.030000 0.630000 3.330000 5.430000 ;
      RECT 3.630000 0.330000 3.930000 5.130000 ;
      RECT 4.230000 0.630000 4.530000 5.430000 ;
      RECT 4.830000 0.330000 5.130000 5.130000 ;
      RECT 5.430000 0.330000 5.900000 5.430000 ;
    LAYER via ;
      RECT 0.035000 0.680000 0.295000 0.940000 ;
      RECT 0.035000 1.080000 0.295000 1.340000 ;
      RECT 0.035000 1.480000 0.295000 1.740000 ;
      RECT 0.035000 1.880000 0.295000 2.140000 ;
      RECT 0.035000 2.280000 0.295000 2.540000 ;
      RECT 0.035000 2.680000 0.295000 2.940000 ;
      RECT 0.035000 3.080000 0.295000 3.340000 ;
      RECT 0.035000 3.480000 0.295000 3.740000 ;
      RECT 0.035000 3.880000 0.295000 4.140000 ;
      RECT 0.035000 4.280000 0.295000 4.540000 ;
      RECT 0.035000 4.680000 0.295000 4.940000 ;
      RECT 0.035000 5.080000 0.295000 5.340000 ;
      RECT 0.280000 0.035000 0.540000 0.295000 ;
      RECT 0.680000 0.035000 0.940000 0.295000 ;
      RECT 0.735000 5.535000 0.995000 5.795000 ;
      RECT 1.080000 0.035000 1.340000 0.295000 ;
      RECT 1.135000 5.535000 1.395000 5.795000 ;
      RECT 1.480000 0.035000 1.740000 0.295000 ;
      RECT 1.535000 5.535000 1.795000 5.795000 ;
      RECT 1.880000 0.035000 2.140000 0.295000 ;
      RECT 1.935000 5.535000 2.195000 5.795000 ;
      RECT 2.280000 0.035000 2.540000 0.295000 ;
      RECT 2.335000 5.535000 2.595000 5.795000 ;
      RECT 2.680000 0.035000 2.940000 0.295000 ;
      RECT 2.735000 5.535000 2.995000 5.795000 ;
      RECT 3.080000 0.035000 3.340000 0.295000 ;
      RECT 3.135000 5.535000 3.395000 5.795000 ;
      RECT 3.480000 0.035000 3.740000 0.295000 ;
      RECT 3.535000 5.535000 3.795000 5.795000 ;
      RECT 3.880000 0.035000 4.140000 0.295000 ;
      RECT 3.935000 5.535000 4.195000 5.795000 ;
      RECT 4.280000 0.035000 4.540000 0.295000 ;
      RECT 4.335000 5.535000 4.595000 5.795000 ;
      RECT 4.680000 0.035000 4.940000 0.295000 ;
      RECT 4.735000 5.535000 4.995000 5.795000 ;
      RECT 5.080000 0.035000 5.340000 0.295000 ;
      RECT 5.135000 5.535000 5.395000 5.795000 ;
      RECT 5.535000 0.735000 5.795000 0.995000 ;
      RECT 5.535000 1.135000 5.795000 1.395000 ;
      RECT 5.535000 1.535000 5.795000 1.795000 ;
      RECT 5.535000 1.935000 5.795000 2.195000 ;
      RECT 5.535000 2.335000 5.795000 2.595000 ;
      RECT 5.535000 2.735000 5.795000 2.995000 ;
      RECT 5.535000 3.135000 5.795000 3.395000 ;
      RECT 5.535000 3.535000 5.795000 3.795000 ;
      RECT 5.535000 3.935000 5.795000 4.195000 ;
      RECT 5.535000 4.335000 5.795000 4.595000 ;
      RECT 5.535000 4.735000 5.795000 4.995000 ;
      RECT 5.535000 5.135000 5.795000 5.395000 ;
    LAYER via2 ;
      RECT 0.025000 0.390000 0.305000 0.670000 ;
      RECT 0.025000 1.020000 0.305000 1.300000 ;
      RECT 0.025000 1.650000 0.305000 1.930000 ;
      RECT 0.025000 2.280000 0.305000 2.560000 ;
      RECT 0.025000 2.910000 0.305000 3.190000 ;
      RECT 0.025000 3.540000 0.305000 3.820000 ;
      RECT 0.025000 4.170000 0.305000 4.450000 ;
      RECT 0.025000 4.800000 0.305000 5.080000 ;
      RECT 0.390000 0.025000 0.670000 0.305000 ;
      RECT 0.485000 5.525000 0.765000 5.805000 ;
      RECT 1.020000 0.025000 1.300000 0.305000 ;
      RECT 1.115000 5.525000 1.395000 5.805000 ;
      RECT 1.650000 0.025000 1.930000 0.305000 ;
      RECT 1.745000 5.525000 2.025000 5.805000 ;
      RECT 2.280000 0.025000 2.560000 0.305000 ;
      RECT 2.375000 5.525000 2.655000 5.805000 ;
      RECT 2.910000 0.025000 3.190000 0.305000 ;
      RECT 3.005000 5.525000 3.285000 5.805000 ;
      RECT 3.540000 0.025000 3.820000 0.305000 ;
      RECT 3.635000 5.525000 3.915000 5.805000 ;
      RECT 4.170000 0.025000 4.450000 0.305000 ;
      RECT 4.265000 5.525000 4.545000 5.805000 ;
      RECT 4.800000 0.025000 5.080000 0.305000 ;
      RECT 4.895000 5.525000 5.175000 5.805000 ;
      RECT 5.525000 0.485000 5.805000 0.765000 ;
      RECT 5.525000 1.115000 5.805000 1.395000 ;
      RECT 5.525000 1.745000 5.805000 2.025000 ;
      RECT 5.525000 2.375000 5.805000 2.655000 ;
      RECT 5.525000 3.005000 5.805000 3.285000 ;
      RECT 5.525000 3.635000 5.805000 3.915000 ;
      RECT 5.525000 4.265000 5.805000 4.545000 ;
      RECT 5.525000 4.895000 5.805000 5.175000 ;
    LAYER via3 ;
      RECT 0.005000 0.370000 0.325000 0.690000 ;
      RECT 0.005000 1.000000 0.325000 1.320000 ;
      RECT 0.005000 1.630000 0.325000 1.950000 ;
      RECT 0.005000 2.260000 0.325000 2.580000 ;
      RECT 0.005000 2.890000 0.325000 3.210000 ;
      RECT 0.005000 3.520000 0.325000 3.840000 ;
      RECT 0.005000 4.150000 0.325000 4.470000 ;
      RECT 0.005000 4.780000 0.325000 5.100000 ;
      RECT 0.370000 0.005000 0.690000 0.325000 ;
      RECT 1.000000 0.005000 1.320000 0.325000 ;
      RECT 1.095000 5.505000 1.415000 5.825000 ;
      RECT 1.630000 0.005000 1.950000 0.325000 ;
      RECT 1.725000 5.505000 2.045000 5.825000 ;
      RECT 2.260000 0.005000 2.580000 0.325000 ;
      RECT 2.355000 5.505000 2.675000 5.825000 ;
      RECT 2.890000 0.005000 3.210000 0.325000 ;
      RECT 2.985000 5.505000 3.305000 5.825000 ;
      RECT 3.520000 0.005000 3.840000 0.325000 ;
      RECT 3.615000 5.505000 3.935000 5.825000 ;
      RECT 4.150000 0.005000 4.470000 0.325000 ;
      RECT 4.245000 5.505000 4.565000 5.825000 ;
      RECT 4.780000 0.005000 5.100000 0.325000 ;
      RECT 4.875000 5.505000 5.195000 5.825000 ;
      RECT 5.505000 1.095000 5.825000 1.415000 ;
      RECT 5.505000 1.725000 5.825000 2.045000 ;
      RECT 5.505000 2.355000 5.825000 2.675000 ;
      RECT 5.505000 2.985000 5.825000 3.305000 ;
      RECT 5.505000 3.615000 5.825000 3.935000 ;
      RECT 5.505000 4.245000 5.825000 4.565000 ;
      RECT 5.505000 4.875000 5.825000 5.195000 ;
      RECT 5.505000 5.505000 5.825000 5.825000 ;
  END
END sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap
END LIBRARY
