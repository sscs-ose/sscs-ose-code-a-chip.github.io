magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -307 -4582 307 4582
<< psubdiff >>
rect -271 4512 -175 4546
rect 175 4512 271 4546
rect -271 4450 -237 4512
rect 237 4450 271 4512
rect -271 -4512 -237 -4450
rect 237 -4512 271 -4450
rect -271 -4546 -175 -4512
rect 175 -4546 271 -4512
<< psubdiffcont >>
rect -175 4512 175 4546
rect -271 -4450 -237 4450
rect 237 -4450 271 4450
rect -175 -4546 175 -4512
<< xpolycontact >>
rect -141 3984 141 4416
rect -141 -4416 141 -3984
<< ppolyres >>
rect -141 -3984 141 3984
<< locali >>
rect -271 4512 -175 4546
rect 175 4512 271 4546
rect -271 4450 -237 4512
rect 237 4450 271 4512
rect -271 -4512 -237 -4450
rect 237 -4512 271 -4450
rect -271 -4546 -175 -4512
rect 175 -4546 271 -4512
<< viali >>
rect -125 4001 125 4398
rect -125 -4398 125 -4001
<< metal1 >>
rect -131 4398 131 4410
rect -131 4001 -125 4398
rect 125 4001 131 4398
rect -131 3989 131 4001
rect -131 -4001 131 -3989
rect -131 -4398 -125 -4001
rect 125 -4398 131 -4001
rect -131 -4410 131 -4398
<< labels >>
rlabel psubdiffcont 0 -4529 0 -4529 0 B
port 1 nsew
rlabel xpolycontact 0 4381 0 4381 0 R1
port 2 nsew
rlabel xpolycontact 0 -4381 0 -4381 0 R2
port 3 nsew
<< properties >>
string FIXED_BBOX -254 -4529 254 4529
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 40.0 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 319.8 val 9.348k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1 mult 1
<< end >>
