magic
tech sky130A
magscale 1 2
timestamp 1762084523
<< error_p >>
rect -29 -24007 29 -24001
rect -29 -24041 -17 -24007
rect -29 -24047 29 -24041
<< pwell >>
rect -211 -24179 211 24179
<< nmos >>
rect -15 -23969 15 24031
<< ndiff >>
rect -73 24019 -15 24031
rect -73 -23957 -61 24019
rect -27 -23957 -15 24019
rect -73 -23969 -15 -23957
rect 15 24019 73 24031
rect 15 -23957 27 24019
rect 61 -23957 73 24019
rect 15 -23969 73 -23957
<< ndiffc >>
rect -61 -23957 -27 24019
rect 27 -23957 61 24019
<< psubdiff >>
rect -175 24109 -79 24143
rect 79 24109 175 24143
rect -175 24047 -141 24109
rect 141 24047 175 24109
rect -175 -24109 -141 -24047
rect 141 -24109 175 -24047
rect -175 -24143 -79 -24109
rect 79 -24143 175 -24109
<< psubdiffcont >>
rect -79 24109 79 24143
rect -175 -24047 -141 24047
rect 141 -24047 175 24047
rect -79 -24143 79 -24109
<< poly >>
rect -15 24031 15 24057
rect -15 -23991 15 -23969
rect -33 -24007 33 -23991
rect -33 -24041 -17 -24007
rect 17 -24041 33 -24007
rect -33 -24057 33 -24041
<< polycont >>
rect -17 -24041 17 -24007
<< locali >>
rect -175 24109 -79 24143
rect 79 24109 175 24143
rect -175 24047 -141 24109
rect 141 24047 175 24109
rect -61 24019 -27 24035
rect -61 -23973 -27 -23957
rect 27 24019 61 24035
rect 27 -23973 61 -23957
rect -33 -24041 -17 -24007
rect 17 -24041 33 -24007
rect -175 -24109 -141 -24047
rect 141 -24109 175 -24047
rect -175 -24143 -79 -24109
rect 79 -24143 175 -24109
<< viali >>
rect -61 -23957 -27 24019
rect 27 -23957 61 24019
rect -17 -24041 17 -24007
<< metal1 >>
rect -67 24019 -21 24031
rect -67 -23957 -61 24019
rect -27 -23957 -21 24019
rect -67 -23969 -21 -23957
rect 21 24019 67 24031
rect 21 -23957 27 24019
rect 61 -23957 67 24019
rect 21 -23969 67 -23957
rect -29 -24007 29 -24001
rect -29 -24041 -17 -24007
rect 17 -24041 29 -24007
rect -29 -24047 29 -24041
<< labels >>
rlabel psubdiffcont 0 -24126 0 -24126 0 B
port 1 nsew
rlabel ndiffc -44 31 -44 31 0 D
port 2 nsew
rlabel ndiffc 44 31 44 31 0 S
port 3 nsew
rlabel polycont 0 -24024 0 -24024 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -24126 158 24126
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 240 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
