VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_0kbytes_1rw_32x128_32
   CLASS BLOCK ;
   SIZE 288.4 BY 300.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.26 0.0 78.64 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.1 0.0 84.48 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.94 0.0 90.32 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.78 0.0 96.16 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  101.62 0.0 102.0 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.46 0.0 107.84 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.3 0.0 113.68 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.14 0.0 119.52 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  124.98 0.0 125.36 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.82 0.0 131.2 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.66 0.0 137.04 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.5 0.0 142.88 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.34 0.0 148.72 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.18 0.0 154.56 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.02 0.0 160.4 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.86 0.0 166.24 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.7 0.0 172.08 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.54 0.0 177.92 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.38 0.0 183.76 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.22 0.0 189.6 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.06 0.0 195.44 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  200.9 0.0 201.28 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.74 0.0 207.12 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.58 0.0 212.96 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.42 0.0 218.8 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.26 0.0 224.64 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.1 0.0 230.48 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.94 0.0 236.32 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.78 0.0 242.16 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.62 0.0 248.0 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.46 0.0 253.84 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.3 0.0 259.68 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 117.985 0.38 118.365 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 126.385 0.38 126.765 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 132.35 0.38 132.73 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.85 0.38 141.23 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 146.49 0.38 146.87 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.99 0.38 155.37 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 159.985 0.38 160.365 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.385 0.38 168.765 ;
      END
   END addr0[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 23.37 0.38 23.75 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.565 0.0 140.945 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  145.1 0.0 145.48 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.25 0.0 146.63 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.1 0.0 150.48 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.25 0.0 151.63 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.1 0.0 155.48 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  156.25 0.0 156.63 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.71 0.0 161.09 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.63 0.0 163.01 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.72 0.0 164.1 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.55 0.0 166.93 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  169.895 0.0 170.275 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.63 0.0 173.01 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  175.1 0.0 175.48 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.23 0.0 178.61 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.1 0.0 180.48 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  181.25 0.0 181.63 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.1 0.0 185.48 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.25 0.0 186.63 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.1 0.0 190.48 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.25 0.0 191.63 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.75 0.0 196.13 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.63 0.0 198.01 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.72 0.0 199.1 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.59 0.0 201.97 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.935 0.0 205.315 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.63 0.0 208.01 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.1 0.0 210.48 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.27 0.0 213.65 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.1 0.0 215.48 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.25 0.0 216.63 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.1 0.0 220.48 0.38 ;
      END
   END dout0[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 300.62 ;
         LAYER met3 ;
         RECT  0.0 0.0 288.4 1.74 ;
         LAYER met3 ;
         RECT  0.0 298.88 288.4 300.62 ;
         LAYER met4 ;
         RECT  286.66 0.0 288.4 300.62 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 3.48 284.92 5.22 ;
         LAYER met4 ;
         RECT  283.18 3.48 284.92 297.14 ;
         LAYER met3 ;
         RECT  3.48 295.4 284.92 297.14 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 297.14 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 287.78 300.0 ;
   LAYER  met2 ;
      RECT  0.62 0.62 287.78 300.0 ;
   LAYER  met3 ;
      RECT  0.98 117.385 287.78 118.965 ;
      RECT  0.62 118.965 0.98 125.785 ;
      RECT  0.62 127.365 0.98 131.75 ;
      RECT  0.62 133.33 0.98 140.25 ;
      RECT  0.62 141.83 0.98 145.89 ;
      RECT  0.62 147.47 0.98 154.39 ;
      RECT  0.62 155.97 0.98 159.385 ;
      RECT  0.62 160.965 0.98 167.785 ;
      RECT  0.62 15.85 0.98 22.77 ;
      RECT  0.62 24.35 0.98 117.385 ;
      RECT  0.62 2.34 0.98 14.27 ;
      RECT  0.62 169.365 0.98 298.28 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 117.385 ;
      RECT  2.88 2.34 285.52 2.88 ;
      RECT  2.88 5.82 285.52 117.385 ;
      RECT  285.52 2.34 287.78 2.88 ;
      RECT  285.52 2.88 287.78 5.82 ;
      RECT  285.52 5.82 287.78 117.385 ;
      RECT  0.98 118.965 2.88 294.8 ;
      RECT  0.98 294.8 2.88 297.74 ;
      RECT  0.98 297.74 2.88 298.28 ;
      RECT  2.88 118.965 285.52 294.8 ;
      RECT  2.88 297.74 285.52 298.28 ;
      RECT  285.52 118.965 287.78 294.8 ;
      RECT  285.52 294.8 287.78 297.74 ;
      RECT  285.52 297.74 287.78 298.28 ;
   LAYER  met4 ;
      RECT  77.66 0.98 79.24 300.0 ;
      RECT  79.24 0.62 83.5 0.98 ;
      RECT  85.08 0.62 89.34 0.98 ;
      RECT  90.92 0.62 95.18 0.98 ;
      RECT  96.76 0.62 101.02 0.98 ;
      RECT  102.6 0.62 106.86 0.98 ;
      RECT  108.44 0.62 112.7 0.98 ;
      RECT  114.28 0.62 118.54 0.98 ;
      RECT  120.12 0.62 124.38 0.98 ;
      RECT  125.96 0.62 130.22 0.98 ;
      RECT  131.8 0.62 136.06 0.98 ;
      RECT  225.24 0.62 229.5 0.98 ;
      RECT  231.08 0.62 235.34 0.98 ;
      RECT  236.92 0.62 241.18 0.98 ;
      RECT  242.76 0.62 247.02 0.98 ;
      RECT  248.6 0.62 252.86 0.98 ;
      RECT  254.44 0.62 258.7 0.98 ;
      RECT  260.28 0.62 264.54 0.98 ;
      RECT  32.08 0.62 77.66 0.98 ;
      RECT  266.12 0.62 270.38 0.98 ;
      RECT  137.64 0.62 139.965 0.98 ;
      RECT  141.545 0.62 141.9 0.98 ;
      RECT  143.48 0.62 144.5 0.98 ;
      RECT  147.23 0.62 147.74 0.98 ;
      RECT  149.32 0.62 149.5 0.98 ;
      RECT  152.23 0.62 153.58 0.98 ;
      RECT  157.23 0.62 159.42 0.98 ;
      RECT  161.69 0.62 162.03 0.98 ;
      RECT  164.7 0.62 165.26 0.98 ;
      RECT  167.53 0.62 169.295 0.98 ;
      RECT  170.875 0.62 171.1 0.98 ;
      RECT  173.61 0.62 174.5 0.98 ;
      RECT  176.08 0.62 176.94 0.98 ;
      RECT  179.21 0.62 179.5 0.98 ;
      RECT  182.23 0.62 182.78 0.98 ;
      RECT  184.36 0.62 184.5 0.98 ;
      RECT  187.23 0.62 188.62 0.98 ;
      RECT  192.23 0.62 194.46 0.98 ;
      RECT  196.73 0.62 197.03 0.98 ;
      RECT  199.7 0.62 200.3 0.98 ;
      RECT  202.57 0.62 204.335 0.98 ;
      RECT  205.915 0.62 206.14 0.98 ;
      RECT  208.61 0.62 209.5 0.98 ;
      RECT  211.08 0.62 211.98 0.98 ;
      RECT  214.25 0.62 214.5 0.98 ;
      RECT  217.23 0.62 217.82 0.98 ;
      RECT  219.4 0.62 219.5 0.98 ;
      RECT  222.23 0.62 223.66 0.98 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  271.96 0.62 286.06 0.98 ;
      RECT  79.24 0.98 282.58 2.88 ;
      RECT  79.24 2.88 282.58 297.74 ;
      RECT  79.24 297.74 282.58 300.0 ;
      RECT  282.58 0.98 285.52 2.88 ;
      RECT  282.58 297.74 285.52 300.0 ;
      RECT  285.52 0.98 286.06 2.88 ;
      RECT  285.52 2.88 286.06 297.74 ;
      RECT  285.52 297.74 286.06 300.0 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 297.74 ;
      RECT  2.34 297.74 2.88 300.0 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 297.74 5.82 300.0 ;
      RECT  5.82 0.98 77.66 2.88 ;
      RECT  5.82 2.88 77.66 297.74 ;
      RECT  5.82 297.74 77.66 300.0 ;
   END
END    sky130_sram_0kbytes_1rw_32x128_32
END    LIBRARY