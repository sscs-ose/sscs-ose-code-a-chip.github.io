* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 3
.param
+ sky130_fd_pr__esd_nfet_01v8__toxe_mult = 1.0365
+ sky130_fd_pr__esd_nfet_01v8__rshn_mult = 1.0
+ sky130_fd_pr__esd_nfet_01v8__overlap_mult = 1.0142
+ sky130_fd_pr__esd_nfet_01v8__ajunction_mult = 1.1505e+0
+ sky130_fd_pr__esd_nfet_01v8__pjunction_mult = 1.1793e+0
+ sky130_fd_pr__esd_nfet_01v8__lint_diff = -1.21275e-8
+ sky130_fd_pr__esd_nfet_01v8__wint_diff = 2.252e-8
+ sky130_fd_pr__esd_nfet_01v8__dlc_diff = -10.107e-9
+ sky130_fd_pr__esd_nfet_01v8__dwc_diff = 2.252e-8
*
* sky130_fd_pr__esd_nfet_01v8, Bin 000, W = 20.35, L = 0.165
* ----------------------------------------
+ sky130_fd_pr__esd_nfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_0 = 1.7885e-10
+ sky130_fd_pr__esd_nfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__voff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_0 = 0.0055748
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_0 = -7.1805e-20
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_0 = 0.042026
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_0 = 0.0012233
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_0 = 14958.0
+ sky130_fd_pr__esd_nfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0 = 0.27275
+ sky130_fd_pr__esd_nfet_01v8__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__ags_diff_0 = 0.0
*
* sky130_fd_pr__esd_nfet_01v8, Bin 001, W = 40.31, L = 0.165
* ----------------------------------------
+ sky130_fd_pr__esd_nfet_01v8__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_1 = 1.3726e-10
+ sky130_fd_pr__esd_nfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__voff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_1 = -0.013821
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_1 = 2.5211e-19
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_1 = 0.036092
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_1 = 0.0022928
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_1 = 5065.5
+ sky130_fd_pr__esd_nfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1 = -0.30661
+ sky130_fd_pr__esd_nfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__b0_diff_1 = 0.0
*
* sky130_fd_pr__esd_nfet_01v8, Bin 002, W = 5.4, L = 0.18
* -------------------------------------
+ sky130_fd_pr__esd_nfet_01v8__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__ags_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_2 = 1.5043e-10
+ sky130_fd_pr__esd_nfet_01v8__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__voff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_2 = -0.005198
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_2 = -2.1082e-19
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_2 = 0.035849
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_2 = 0.00062049
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_2 = 13857.0
+ sky130_fd_pr__esd_nfet_01v8__kt1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2 = -0.46399
+ sky130_fd_pr__esd_nfet_01v8__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2 = 0.0
.include "sky130_fd_pr__esd_nfet_01v8.pm3.spice"
