MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 19.51 BY 45.28 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.73 30.92 4.01 35.44 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 4.16 12.02 4.44 29.98 ;
      LAYER M3 ;
        RECT 16.2 6.56 16.48 30.4 ;
      LAYER M3 ;
        RECT 4.16 19.555 4.44 19.925 ;
      LAYER M2 ;
        RECT 4.3 19.6 16.34 19.88 ;
      LAYER M3 ;
        RECT 16.2 19.555 16.48 19.925 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 13.62 35.54 13.9 41.74 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 13.19 35.96 13.47 42.16 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 3.73 11.6 4.01 29.56 ;
  LAYER M2 ;
        RECT 3.27 31.36 5.33 31.64 ;
  LAYER M3 ;
        RECT 12.76 32.18 13.04 38.38 ;
  LAYER M3 ;
        RECT 3.73 28.795 4.01 29.165 ;
  LAYER M2 ;
        RECT 3.721 28.84 4.019 29.12 ;
  LAYER M1 ;
        RECT 3.745 28.98 3.995 31.5 ;
  LAYER M2 ;
        RECT 3.71 31.36 4.03 31.64 ;
  LAYER M2 ;
        RECT 5.16 31.36 10.32 31.64 ;
  LAYER M3 ;
        RECT 10.18 31.379 10.46 31.621 ;
  LAYER M4 ;
        RECT 10.32 31.1 12.9 31.9 ;
  LAYER M3 ;
        RECT 12.76 31.5 13.04 32.34 ;
  LAYER M1 ;
        RECT 3.745 28.895 3.995 29.065 ;
  LAYER M2 ;
        RECT 3.7 28.84 4.04 29.12 ;
  LAYER M1 ;
        RECT 3.745 31.415 3.995 31.585 ;
  LAYER M2 ;
        RECT 3.7 31.36 4.04 31.64 ;
  LAYER M2 ;
        RECT 3.71 28.84 4.03 29.12 ;
  LAYER M3 ;
        RECT 3.73 28.82 4.01 29.14 ;
  LAYER M1 ;
        RECT 3.745 31.415 3.995 31.585 ;
  LAYER M2 ;
        RECT 3.7 31.36 4.04 31.64 ;
  LAYER M1 ;
        RECT 3.745 31.415 3.995 31.585 ;
  LAYER M2 ;
        RECT 3.7 31.36 4.04 31.64 ;
  LAYER M2 ;
        RECT 10.16 31.36 10.48 31.64 ;
  LAYER M3 ;
        RECT 10.18 31.34 10.46 31.66 ;
  LAYER M3 ;
        RECT 10.18 31.315 10.46 31.685 ;
  LAYER M4 ;
        RECT 10.155 31.1 10.485 31.9 ;
  LAYER M3 ;
        RECT 12.76 31.315 13.04 31.685 ;
  LAYER M4 ;
        RECT 12.735 31.1 13.065 31.9 ;
  LAYER M1 ;
        RECT 3.745 31.415 3.995 31.585 ;
  LAYER M2 ;
        RECT 3.7 31.36 4.04 31.64 ;
  LAYER M3 ;
        RECT 12.76 31.315 13.04 31.685 ;
  LAYER M4 ;
        RECT 12.735 31.1 13.065 31.9 ;
  LAYER M3 ;
        RECT 15.77 2.78 16.05 30.82 ;
  LAYER M3 ;
        RECT 14.48 31.34 14.76 37.54 ;
  LAYER M3 ;
        RECT 15.77 30.66 16.05 31.08 ;
  LAYER M2 ;
        RECT 14.62 30.94 15.91 31.22 ;
  LAYER M3 ;
        RECT 14.48 31.08 14.76 31.5 ;
  LAYER M2 ;
        RECT 14.46 30.94 14.78 31.22 ;
  LAYER M3 ;
        RECT 14.48 30.92 14.76 31.24 ;
  LAYER M2 ;
        RECT 15.75 30.94 16.07 31.22 ;
  LAYER M3 ;
        RECT 15.77 30.92 16.05 31.24 ;
  LAYER M2 ;
        RECT 14.46 30.94 14.78 31.22 ;
  LAYER M3 ;
        RECT 14.48 30.92 14.76 31.24 ;
  LAYER M2 ;
        RECT 15.75 30.94 16.07 31.22 ;
  LAYER M3 ;
        RECT 15.77 30.92 16.05 31.24 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 30.82 ;
  LAYER M3 ;
        RECT 14.05 31.76 14.33 37.96 ;
  LAYER M3 ;
        RECT 11.47 30.66 11.75 31.08 ;
  LAYER M2 ;
        RECT 11.61 30.94 13.76 31.22 ;
  LAYER M3 ;
        RECT 13.62 31.08 13.9 31.5 ;
  LAYER M4 ;
        RECT 13.76 31.1 14.19 31.9 ;
  LAYER M3 ;
        RECT 14.05 31.5 14.33 31.92 ;
  LAYER M2 ;
        RECT 11.45 30.94 11.77 31.22 ;
  LAYER M3 ;
        RECT 11.47 30.92 11.75 31.24 ;
  LAYER M2 ;
        RECT 13.6 30.94 13.92 31.22 ;
  LAYER M3 ;
        RECT 13.62 30.92 13.9 31.24 ;
  LAYER M3 ;
        RECT 13.62 31.315 13.9 31.685 ;
  LAYER M4 ;
        RECT 13.595 31.1 13.925 31.9 ;
  LAYER M3 ;
        RECT 14.05 31.315 14.33 31.685 ;
  LAYER M4 ;
        RECT 14.025 31.1 14.355 31.9 ;
  LAYER M2 ;
        RECT 11.45 30.94 11.77 31.22 ;
  LAYER M3 ;
        RECT 11.47 30.92 11.75 31.24 ;
  LAYER M2 ;
        RECT 13.6 30.94 13.92 31.22 ;
  LAYER M3 ;
        RECT 13.62 30.92 13.9 31.24 ;
  LAYER M3 ;
        RECT 13.62 31.315 13.9 31.685 ;
  LAYER M4 ;
        RECT 13.595 31.1 13.925 31.9 ;
  LAYER M3 ;
        RECT 14.05 31.315 14.33 31.685 ;
  LAYER M4 ;
        RECT 14.025 31.1 14.355 31.9 ;
  LAYER M3 ;
        RECT 4.59 8.24 4.87 30.4 ;
  LAYER M3 ;
        RECT 11.04 6.56 11.32 30.4 ;
  LAYER M3 ;
        RECT 4.59 18.715 4.87 19.085 ;
  LAYER M4 ;
        RECT 4.73 18.5 11.18 19.3 ;
  LAYER M3 ;
        RECT 11.04 18.715 11.32 19.085 ;
  LAYER M3 ;
        RECT 4.59 18.715 4.87 19.085 ;
  LAYER M4 ;
        RECT 4.565 18.5 4.895 19.3 ;
  LAYER M3 ;
        RECT 11.04 18.715 11.32 19.085 ;
  LAYER M4 ;
        RECT 11.015 18.5 11.345 19.3 ;
  LAYER M3 ;
        RECT 4.59 18.715 4.87 19.085 ;
  LAYER M4 ;
        RECT 4.565 18.5 4.895 19.3 ;
  LAYER M3 ;
        RECT 11.04 18.715 11.32 19.085 ;
  LAYER M4 ;
        RECT 11.015 18.5 11.345 19.3 ;
  LAYER M1 ;
        RECT 1.595 30.995 1.845 34.525 ;
  LAYER M1 ;
        RECT 1.595 34.775 1.845 35.785 ;
  LAYER M1 ;
        RECT 1.595 36.875 1.845 37.885 ;
  LAYER M1 ;
        RECT 0.735 30.995 0.985 34.525 ;
  LAYER M1 ;
        RECT 2.455 30.995 2.705 34.525 ;
  LAYER M1 ;
        RECT 3.315 30.995 3.565 34.525 ;
  LAYER M1 ;
        RECT 3.315 34.775 3.565 35.785 ;
  LAYER M1 ;
        RECT 3.315 36.875 3.565 37.885 ;
  LAYER M1 ;
        RECT 4.175 30.995 4.425 34.525 ;
  LAYER M1 ;
        RECT 5.035 30.995 5.285 34.525 ;
  LAYER M1 ;
        RECT 5.035 34.775 5.285 35.785 ;
  LAYER M1 ;
        RECT 5.035 36.875 5.285 37.885 ;
  LAYER M1 ;
        RECT 5.895 30.995 6.145 34.525 ;
  LAYER M1 ;
        RECT 6.755 30.995 7.005 34.525 ;
  LAYER M1 ;
        RECT 6.755 34.775 7.005 35.785 ;
  LAYER M1 ;
        RECT 6.755 36.875 7.005 37.885 ;
  LAYER M1 ;
        RECT 7.615 30.995 7.865 34.525 ;
  LAYER M2 ;
        RECT 1.55 30.94 7.05 31.22 ;
  LAYER M2 ;
        RECT 1.55 35.14 7.05 35.42 ;
  LAYER M2 ;
        RECT 0.69 31.78 7.91 32.06 ;
  LAYER M2 ;
        RECT 1.55 37.24 7.05 37.52 ;
  LAYER M3 ;
        RECT 3.73 30.92 4.01 35.44 ;
  LAYER M2 ;
        RECT 3.27 31.36 5.33 31.64 ;
  LAYER M3 ;
        RECT 4.59 31.76 4.87 37.54 ;
  LAYER M1 ;
        RECT 15.355 27.215 15.605 30.745 ;
  LAYER M1 ;
        RECT 15.355 25.955 15.605 26.965 ;
  LAYER M1 ;
        RECT 15.355 21.335 15.605 24.865 ;
  LAYER M1 ;
        RECT 15.355 20.075 15.605 21.085 ;
  LAYER M1 ;
        RECT 15.355 15.455 15.605 18.985 ;
  LAYER M1 ;
        RECT 15.355 14.195 15.605 15.205 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 8.315 15.605 9.325 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 15.355 2.435 15.605 3.445 ;
  LAYER M1 ;
        RECT 15.355 0.335 15.605 1.345 ;
  LAYER M1 ;
        RECT 14.495 27.215 14.745 30.745 ;
  LAYER M1 ;
        RECT 14.495 21.335 14.745 24.865 ;
  LAYER M1 ;
        RECT 14.495 15.455 14.745 18.985 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 16.215 27.215 16.465 30.745 ;
  LAYER M1 ;
        RECT 16.215 21.335 16.465 24.865 ;
  LAYER M1 ;
        RECT 16.215 15.455 16.465 18.985 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 17.075 27.215 17.325 30.745 ;
  LAYER M1 ;
        RECT 17.075 25.955 17.325 26.965 ;
  LAYER M1 ;
        RECT 17.075 21.335 17.325 24.865 ;
  LAYER M1 ;
        RECT 17.075 20.075 17.325 21.085 ;
  LAYER M1 ;
        RECT 17.075 15.455 17.325 18.985 ;
  LAYER M1 ;
        RECT 17.075 14.195 17.325 15.205 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 8.315 17.325 9.325 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 17.075 2.435 17.325 3.445 ;
  LAYER M1 ;
        RECT 17.075 0.335 17.325 1.345 ;
  LAYER M1 ;
        RECT 17.935 27.215 18.185 30.745 ;
  LAYER M1 ;
        RECT 17.935 21.335 18.185 24.865 ;
  LAYER M1 ;
        RECT 17.935 15.455 18.185 18.985 ;
  LAYER M1 ;
        RECT 17.935 9.575 18.185 13.105 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M2 ;
        RECT 14.88 30.52 16.08 30.8 ;
  LAYER M2 ;
        RECT 15.31 26.32 17.37 26.6 ;
  LAYER M2 ;
        RECT 16.17 30.1 17.37 30.38 ;
  LAYER M2 ;
        RECT 14.45 29.68 18.23 29.96 ;
  LAYER M2 ;
        RECT 15.74 24.64 17.37 24.92 ;
  LAYER M2 ;
        RECT 15.31 20.44 17.37 20.72 ;
  LAYER M2 ;
        RECT 15.31 24.22 16.51 24.5 ;
  LAYER M2 ;
        RECT 14.45 23.8 18.23 24.08 ;
  LAYER M2 ;
        RECT 14.88 18.76 16.08 19.04 ;
  LAYER M2 ;
        RECT 15.31 14.56 17.37 14.84 ;
  LAYER M2 ;
        RECT 16.17 18.34 17.37 18.62 ;
  LAYER M2 ;
        RECT 14.45 17.92 18.23 18.2 ;
  LAYER M2 ;
        RECT 15.74 12.88 17.37 13.16 ;
  LAYER M2 ;
        RECT 15.31 8.68 17.37 8.96 ;
  LAYER M2 ;
        RECT 15.31 12.46 16.51 12.74 ;
  LAYER M2 ;
        RECT 14.45 12.04 18.23 12.32 ;
  LAYER M2 ;
        RECT 14.88 7 16.08 7.28 ;
  LAYER M2 ;
        RECT 15.31 2.8 17.37 3.08 ;
  LAYER M2 ;
        RECT 16.17 6.58 17.37 6.86 ;
  LAYER M2 ;
        RECT 14.45 6.16 18.23 6.44 ;
  LAYER M2 ;
        RECT 15.31 0.7 17.37 0.98 ;
  LAYER M3 ;
        RECT 15.77 2.78 16.05 30.82 ;
  LAYER M3 ;
        RECT 16.2 6.56 16.48 30.4 ;
  LAYER M3 ;
        RECT 16.63 0.68 16.91 29.98 ;
  LAYER M1 ;
        RECT 11.915 27.215 12.165 30.745 ;
  LAYER M1 ;
        RECT 11.915 25.955 12.165 26.965 ;
  LAYER M1 ;
        RECT 11.915 21.335 12.165 24.865 ;
  LAYER M1 ;
        RECT 11.915 20.075 12.165 21.085 ;
  LAYER M1 ;
        RECT 11.915 15.455 12.165 18.985 ;
  LAYER M1 ;
        RECT 11.915 14.195 12.165 15.205 ;
  LAYER M1 ;
        RECT 11.915 9.575 12.165 13.105 ;
  LAYER M1 ;
        RECT 11.915 8.315 12.165 9.325 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.915 2.435 12.165 3.445 ;
  LAYER M1 ;
        RECT 11.915 0.335 12.165 1.345 ;
  LAYER M1 ;
        RECT 12.775 27.215 13.025 30.745 ;
  LAYER M1 ;
        RECT 12.775 21.335 13.025 24.865 ;
  LAYER M1 ;
        RECT 12.775 15.455 13.025 18.985 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 11.055 27.215 11.305 30.745 ;
  LAYER M1 ;
        RECT 11.055 21.335 11.305 24.865 ;
  LAYER M1 ;
        RECT 11.055 15.455 11.305 18.985 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.195 27.215 10.445 30.745 ;
  LAYER M1 ;
        RECT 10.195 25.955 10.445 26.965 ;
  LAYER M1 ;
        RECT 10.195 21.335 10.445 24.865 ;
  LAYER M1 ;
        RECT 10.195 20.075 10.445 21.085 ;
  LAYER M1 ;
        RECT 10.195 15.455 10.445 18.985 ;
  LAYER M1 ;
        RECT 10.195 14.195 10.445 15.205 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 8.315 10.445 9.325 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.195 2.435 10.445 3.445 ;
  LAYER M1 ;
        RECT 10.195 0.335 10.445 1.345 ;
  LAYER M1 ;
        RECT 9.335 27.215 9.585 30.745 ;
  LAYER M1 ;
        RECT 9.335 21.335 9.585 24.865 ;
  LAYER M1 ;
        RECT 9.335 15.455 9.585 18.985 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 11.44 30.52 12.64 30.8 ;
  LAYER M2 ;
        RECT 10.15 26.32 12.21 26.6 ;
  LAYER M2 ;
        RECT 10.15 30.1 11.35 30.38 ;
  LAYER M2 ;
        RECT 9.29 29.68 13.07 29.96 ;
  LAYER M2 ;
        RECT 10.15 24.64 11.78 24.92 ;
  LAYER M2 ;
        RECT 10.15 20.44 12.21 20.72 ;
  LAYER M2 ;
        RECT 11.01 24.22 12.21 24.5 ;
  LAYER M2 ;
        RECT 9.29 23.8 13.07 24.08 ;
  LAYER M2 ;
        RECT 11.44 18.76 12.64 19.04 ;
  LAYER M2 ;
        RECT 10.15 14.56 12.21 14.84 ;
  LAYER M2 ;
        RECT 10.15 18.34 11.35 18.62 ;
  LAYER M2 ;
        RECT 9.29 17.92 13.07 18.2 ;
  LAYER M2 ;
        RECT 10.15 12.88 11.78 13.16 ;
  LAYER M2 ;
        RECT 10.15 8.68 12.21 8.96 ;
  LAYER M2 ;
        RECT 11.01 12.46 12.21 12.74 ;
  LAYER M2 ;
        RECT 9.29 12.04 13.07 12.32 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 10.15 2.8 12.21 3.08 ;
  LAYER M2 ;
        RECT 10.15 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 9.29 6.16 13.07 6.44 ;
  LAYER M2 ;
        RECT 10.15 0.7 12.21 0.98 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 30.82 ;
  LAYER M3 ;
        RECT 11.04 6.56 11.32 30.4 ;
  LAYER M3 ;
        RECT 10.61 0.68 10.89 29.98 ;
  LAYER M1 ;
        RECT 6.755 26.795 7.005 30.325 ;
  LAYER M1 ;
        RECT 6.755 25.535 7.005 26.545 ;
  LAYER M1 ;
        RECT 6.755 20.915 7.005 24.445 ;
  LAYER M1 ;
        RECT 6.755 19.655 7.005 20.665 ;
  LAYER M1 ;
        RECT 6.755 15.035 7.005 18.565 ;
  LAYER M1 ;
        RECT 6.755 13.775 7.005 14.785 ;
  LAYER M1 ;
        RECT 6.755 9.155 7.005 12.685 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 8.905 ;
  LAYER M1 ;
        RECT 6.755 5.795 7.005 6.805 ;
  LAYER M1 ;
        RECT 7.615 26.795 7.865 30.325 ;
  LAYER M1 ;
        RECT 7.615 20.915 7.865 24.445 ;
  LAYER M1 ;
        RECT 7.615 15.035 7.865 18.565 ;
  LAYER M1 ;
        RECT 7.615 9.155 7.865 12.685 ;
  LAYER M1 ;
        RECT 5.895 26.795 6.145 30.325 ;
  LAYER M1 ;
        RECT 5.895 20.915 6.145 24.445 ;
  LAYER M1 ;
        RECT 5.895 15.035 6.145 18.565 ;
  LAYER M1 ;
        RECT 5.895 9.155 6.145 12.685 ;
  LAYER M1 ;
        RECT 5.035 26.795 5.285 30.325 ;
  LAYER M1 ;
        RECT 5.035 25.535 5.285 26.545 ;
  LAYER M1 ;
        RECT 5.035 20.915 5.285 24.445 ;
  LAYER M1 ;
        RECT 5.035 19.655 5.285 20.665 ;
  LAYER M1 ;
        RECT 5.035 15.035 5.285 18.565 ;
  LAYER M1 ;
        RECT 5.035 13.775 5.285 14.785 ;
  LAYER M1 ;
        RECT 5.035 9.155 5.285 12.685 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 8.905 ;
  LAYER M1 ;
        RECT 5.035 5.795 5.285 6.805 ;
  LAYER M1 ;
        RECT 4.175 26.795 4.425 30.325 ;
  LAYER M1 ;
        RECT 4.175 20.915 4.425 24.445 ;
  LAYER M1 ;
        RECT 4.175 15.035 4.425 18.565 ;
  LAYER M1 ;
        RECT 4.175 9.155 4.425 12.685 ;
  LAYER M1 ;
        RECT 3.315 26.795 3.565 30.325 ;
  LAYER M1 ;
        RECT 3.315 25.535 3.565 26.545 ;
  LAYER M1 ;
        RECT 3.315 20.915 3.565 24.445 ;
  LAYER M1 ;
        RECT 3.315 19.655 3.565 20.665 ;
  LAYER M1 ;
        RECT 3.315 15.035 3.565 18.565 ;
  LAYER M1 ;
        RECT 3.315 13.775 3.565 14.785 ;
  LAYER M1 ;
        RECT 3.315 9.155 3.565 12.685 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 8.905 ;
  LAYER M1 ;
        RECT 3.315 5.795 3.565 6.805 ;
  LAYER M1 ;
        RECT 2.455 26.795 2.705 30.325 ;
  LAYER M1 ;
        RECT 2.455 20.915 2.705 24.445 ;
  LAYER M1 ;
        RECT 2.455 15.035 2.705 18.565 ;
  LAYER M1 ;
        RECT 2.455 9.155 2.705 12.685 ;
  LAYER M1 ;
        RECT 1.595 26.795 1.845 30.325 ;
  LAYER M1 ;
        RECT 1.595 25.535 1.845 26.545 ;
  LAYER M1 ;
        RECT 1.595 20.915 1.845 24.445 ;
  LAYER M1 ;
        RECT 1.595 19.655 1.845 20.665 ;
  LAYER M1 ;
        RECT 1.595 15.035 1.845 18.565 ;
  LAYER M1 ;
        RECT 1.595 13.775 1.845 14.785 ;
  LAYER M1 ;
        RECT 1.595 9.155 1.845 12.685 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 8.905 ;
  LAYER M1 ;
        RECT 1.595 5.795 1.845 6.805 ;
  LAYER M1 ;
        RECT 0.735 26.795 0.985 30.325 ;
  LAYER M1 ;
        RECT 0.735 20.915 0.985 24.445 ;
  LAYER M1 ;
        RECT 0.735 15.035 0.985 18.565 ;
  LAYER M1 ;
        RECT 0.735 9.155 0.985 12.685 ;
  LAYER M2 ;
        RECT 1.55 30.1 7.05 30.38 ;
  LAYER M2 ;
        RECT 1.55 25.9 7.05 26.18 ;
  LAYER M2 ;
        RECT 3.27 29.68 5.33 29.96 ;
  LAYER M2 ;
        RECT 0.69 29.26 7.91 29.54 ;
  LAYER M2 ;
        RECT 3.27 24.22 5.33 24.5 ;
  LAYER M2 ;
        RECT 1.55 20.02 7.05 20.3 ;
  LAYER M2 ;
        RECT 1.55 23.8 7.05 24.08 ;
  LAYER M2 ;
        RECT 0.69 23.38 7.91 23.66 ;
  LAYER M2 ;
        RECT 1.55 18.34 7.05 18.62 ;
  LAYER M2 ;
        RECT 1.55 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 3.27 17.92 5.33 18.2 ;
  LAYER M2 ;
        RECT 0.69 17.5 7.91 17.78 ;
  LAYER M2 ;
        RECT 3.27 12.46 5.33 12.74 ;
  LAYER M2 ;
        RECT 1.55 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 1.55 12.04 7.05 12.32 ;
  LAYER M2 ;
        RECT 0.69 11.62 7.91 11.9 ;
  LAYER M2 ;
        RECT 1.55 6.16 7.05 6.44 ;
  LAYER M3 ;
        RECT 4.59 8.24 4.87 30.4 ;
  LAYER M3 ;
        RECT 4.16 12.02 4.44 29.98 ;
  LAYER M3 ;
        RECT 3.73 11.6 4.01 29.56 ;
  LAYER M1 ;
        RECT 16.215 31.415 16.465 34.945 ;
  LAYER M1 ;
        RECT 16.215 35.195 16.465 36.205 ;
  LAYER M1 ;
        RECT 16.215 37.295 16.465 40.825 ;
  LAYER M1 ;
        RECT 16.215 41.075 16.465 42.085 ;
  LAYER M1 ;
        RECT 16.215 43.175 16.465 44.185 ;
  LAYER M1 ;
        RECT 17.075 31.415 17.325 34.945 ;
  LAYER M1 ;
        RECT 17.075 37.295 17.325 40.825 ;
  LAYER M1 ;
        RECT 15.355 31.415 15.605 34.945 ;
  LAYER M1 ;
        RECT 15.355 37.295 15.605 40.825 ;
  LAYER M1 ;
        RECT 14.495 31.415 14.745 34.945 ;
  LAYER M1 ;
        RECT 14.495 35.195 14.745 36.205 ;
  LAYER M1 ;
        RECT 14.495 37.295 14.745 40.825 ;
  LAYER M1 ;
        RECT 14.495 41.075 14.745 42.085 ;
  LAYER M1 ;
        RECT 14.495 43.175 14.745 44.185 ;
  LAYER M1 ;
        RECT 13.635 31.415 13.885 34.945 ;
  LAYER M1 ;
        RECT 13.635 37.295 13.885 40.825 ;
  LAYER M1 ;
        RECT 12.775 31.415 13.025 34.945 ;
  LAYER M1 ;
        RECT 12.775 35.195 13.025 36.205 ;
  LAYER M1 ;
        RECT 12.775 37.295 13.025 40.825 ;
  LAYER M1 ;
        RECT 12.775 41.075 13.025 42.085 ;
  LAYER M1 ;
        RECT 12.775 43.175 13.025 44.185 ;
  LAYER M1 ;
        RECT 11.915 31.415 12.165 34.945 ;
  LAYER M1 ;
        RECT 11.915 37.295 12.165 40.825 ;
  LAYER M1 ;
        RECT 11.055 31.415 11.305 34.945 ;
  LAYER M1 ;
        RECT 11.055 35.195 11.305 36.205 ;
  LAYER M1 ;
        RECT 11.055 37.295 11.305 40.825 ;
  LAYER M1 ;
        RECT 11.055 41.075 11.305 42.085 ;
  LAYER M1 ;
        RECT 11.055 43.175 11.305 44.185 ;
  LAYER M1 ;
        RECT 10.195 31.415 10.445 34.945 ;
  LAYER M1 ;
        RECT 10.195 37.295 10.445 40.825 ;
  LAYER M2 ;
        RECT 11.01 31.36 16.51 31.64 ;
  LAYER M2 ;
        RECT 12.73 31.78 14.79 32.06 ;
  LAYER M2 ;
        RECT 11.01 35.56 16.51 35.84 ;
  LAYER M2 ;
        RECT 12.73 35.98 14.79 36.26 ;
  LAYER M2 ;
        RECT 10.15 32.2 17.37 32.48 ;
  LAYER M2 ;
        RECT 12.73 37.24 14.79 37.52 ;
  LAYER M2 ;
        RECT 11.01 37.66 16.51 37.94 ;
  LAYER M2 ;
        RECT 12.73 41.44 14.79 41.72 ;
  LAYER M2 ;
        RECT 11.01 41.86 16.51 42.14 ;
  LAYER M2 ;
        RECT 10.15 38.08 17.37 38.36 ;
  LAYER M2 ;
        RECT 11.01 43.54 16.51 43.82 ;
  LAYER M3 ;
        RECT 14.48 31.34 14.76 37.54 ;
  LAYER M3 ;
        RECT 14.05 31.76 14.33 37.96 ;
  LAYER M3 ;
        RECT 13.62 35.54 13.9 41.74 ;
  LAYER M3 ;
        RECT 13.19 35.96 13.47 42.16 ;
  LAYER M3 ;
        RECT 12.76 32.18 13.04 38.38 ;
  END 
END CURRENT_MIRROR_OTA
