# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25 ;
  ORIGIN -0.050000 -0.050000 ;
  SIZE  2.720000 BY  5.970000 ;
  PIN GATE
    ANTENNAGATEAREA  2.525000 ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.150000 1.915000 0.320000 ;
        RECT 0.905000 5.750000 1.915000 5.920000 ;
      LAYER mcon ;
        RECT 0.965000 0.150000 1.135000 0.320000 ;
        RECT 0.965000 5.750000 1.135000 5.920000 ;
        RECT 1.325000 0.150000 1.495000 0.320000 ;
        RECT 1.325000 5.750000 1.495000 5.920000 ;
        RECT 1.685000 0.150000 1.855000 0.320000 ;
        RECT 1.685000 5.750000 1.855000 5.920000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.905000 0.050000 1.915000 0.380000 ;
        RECT 0.905000 5.690000 1.915000 6.020000 ;
    END
  END GATE
  OBS
    LAYER li1 ;
      RECT 0.240000 0.610000 0.410000 5.460000 ;
      RECT 0.795000 0.490000 0.965000 5.580000 ;
      RECT 1.325000 0.490000 1.495000 5.580000 ;
      RECT 1.855000 0.490000 2.025000 5.580000 ;
      RECT 2.410000 0.610000 2.580000 5.460000 ;
    LAYER mcon ;
      RECT 0.240000 0.970000 0.410000 1.140000 ;
      RECT 0.240000 1.330000 0.410000 1.500000 ;
      RECT 0.240000 1.690000 0.410000 1.860000 ;
      RECT 0.240000 2.050000 0.410000 2.220000 ;
      RECT 0.240000 2.410000 0.410000 2.580000 ;
      RECT 0.240000 2.770000 0.410000 2.940000 ;
      RECT 0.240000 3.130000 0.410000 3.300000 ;
      RECT 0.240000 3.490000 0.410000 3.660000 ;
      RECT 0.240000 3.850000 0.410000 4.020000 ;
      RECT 0.240000 4.210000 0.410000 4.380000 ;
      RECT 0.240000 4.570000 0.410000 4.740000 ;
      RECT 0.240000 4.930000 0.410000 5.100000 ;
      RECT 0.240000 5.290000 0.410000 5.460000 ;
      RECT 0.795000 0.610000 0.965000 0.780000 ;
      RECT 0.795000 0.970000 0.965000 1.140000 ;
      RECT 0.795000 1.330000 0.965000 1.500000 ;
      RECT 0.795000 1.690000 0.965000 1.860000 ;
      RECT 0.795000 2.050000 0.965000 2.220000 ;
      RECT 0.795000 2.410000 0.965000 2.580000 ;
      RECT 0.795000 2.770000 0.965000 2.940000 ;
      RECT 0.795000 3.130000 0.965000 3.300000 ;
      RECT 0.795000 3.490000 0.965000 3.660000 ;
      RECT 0.795000 3.850000 0.965000 4.020000 ;
      RECT 0.795000 4.210000 0.965000 4.380000 ;
      RECT 0.795000 4.570000 0.965000 4.740000 ;
      RECT 0.795000 4.930000 0.965000 5.100000 ;
      RECT 0.795000 5.290000 0.965000 5.460000 ;
      RECT 1.325000 0.610000 1.495000 0.780000 ;
      RECT 1.325000 0.970000 1.495000 1.140000 ;
      RECT 1.325000 1.330000 1.495000 1.500000 ;
      RECT 1.325000 1.690000 1.495000 1.860000 ;
      RECT 1.325000 2.050000 1.495000 2.220000 ;
      RECT 1.325000 2.410000 1.495000 2.580000 ;
      RECT 1.325000 2.770000 1.495000 2.940000 ;
      RECT 1.325000 3.130000 1.495000 3.300000 ;
      RECT 1.325000 3.490000 1.495000 3.660000 ;
      RECT 1.325000 3.850000 1.495000 4.020000 ;
      RECT 1.325000 4.210000 1.495000 4.380000 ;
      RECT 1.325000 4.570000 1.495000 4.740000 ;
      RECT 1.325000 4.930000 1.495000 5.100000 ;
      RECT 1.325000 5.290000 1.495000 5.460000 ;
      RECT 1.855000 0.610000 2.025000 0.780000 ;
      RECT 1.855000 0.970000 2.025000 1.140000 ;
      RECT 1.855000 1.330000 2.025000 1.500000 ;
      RECT 1.855000 1.690000 2.025000 1.860000 ;
      RECT 1.855000 2.050000 2.025000 2.220000 ;
      RECT 1.855000 2.410000 2.025000 2.580000 ;
      RECT 1.855000 2.770000 2.025000 2.940000 ;
      RECT 1.855000 3.130000 2.025000 3.300000 ;
      RECT 1.855000 3.490000 2.025000 3.660000 ;
      RECT 1.855000 3.850000 2.025000 4.020000 ;
      RECT 1.855000 4.210000 2.025000 4.380000 ;
      RECT 1.855000 4.570000 2.025000 4.740000 ;
      RECT 1.855000 4.930000 2.025000 5.100000 ;
      RECT 1.855000 5.290000 2.025000 5.460000 ;
      RECT 2.410000 0.970000 2.580000 1.140000 ;
      RECT 2.410000 1.330000 2.580000 1.500000 ;
      RECT 2.410000 1.690000 2.580000 1.860000 ;
      RECT 2.410000 2.050000 2.580000 2.220000 ;
      RECT 2.410000 2.410000 2.580000 2.580000 ;
      RECT 2.410000 2.770000 2.580000 2.940000 ;
      RECT 2.410000 3.130000 2.580000 3.300000 ;
      RECT 2.410000 3.490000 2.580000 3.660000 ;
      RECT 2.410000 3.850000 2.580000 4.020000 ;
      RECT 2.410000 4.210000 2.580000 4.380000 ;
      RECT 2.410000 4.570000 2.580000 4.740000 ;
      RECT 2.410000 4.930000 2.580000 5.100000 ;
      RECT 2.410000 5.290000 2.580000 5.460000 ;
    LAYER met1 ;
      RECT 0.180000 0.550000 0.470000 5.520000 ;
      RECT 0.750000 0.550000 1.010000 5.520000 ;
      RECT 1.280000 0.550000 1.540000 5.520000 ;
      RECT 1.810000 0.550000 2.070000 5.520000 ;
      RECT 2.350000 0.550000 2.640000 5.520000 ;
    LAYER met2 ;
      RECT 0.050000 0.550000 2.770000 2.910000 ;
      RECT 0.050000 3.160000 2.770000 5.520000 ;
    LAYER via ;
      RECT 0.750000 0.580000 1.010000 0.840000 ;
      RECT 0.750000 0.900000 1.010000 1.160000 ;
      RECT 0.750000 1.220000 1.010000 1.480000 ;
      RECT 0.750000 1.540000 1.010000 1.800000 ;
      RECT 0.750000 1.860000 1.010000 2.120000 ;
      RECT 0.750000 2.180000 1.010000 2.440000 ;
      RECT 0.750000 2.500000 1.010000 2.760000 ;
      RECT 1.280000 3.310000 1.540000 3.570000 ;
      RECT 1.280000 3.630000 1.540000 3.890000 ;
      RECT 1.280000 3.950000 1.540000 4.210000 ;
      RECT 1.280000 4.270000 1.540000 4.530000 ;
      RECT 1.280000 4.590000 1.540000 4.850000 ;
      RECT 1.280000 4.910000 1.540000 5.170000 ;
      RECT 1.280000 5.230000 1.540000 5.490000 ;
      RECT 1.810000 0.580000 2.070000 0.840000 ;
      RECT 1.810000 0.900000 2.070000 1.160000 ;
      RECT 1.810000 1.220000 2.070000 1.480000 ;
      RECT 1.810000 1.540000 2.070000 1.800000 ;
      RECT 1.810000 1.860000 2.070000 2.120000 ;
      RECT 1.810000 2.180000 2.070000 2.440000 ;
      RECT 1.810000 2.500000 2.070000 2.760000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25
END LIBRARY
