* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__nfet_20v0__toxe_mult = 1.06
+ sky130_fd_pr__nfet_20v0__rshn_mult = 1.0
+ sky130_fd_pr__nfet_20v0__overlap_mult = 0.10
+ sky130_fd_pr__nfet_20v0__ajunction_mult = 1.6
+ sky130_fd_pr__nfet_20v0__pjunction_mult = 1.6
+ sky130_fd_pr__nfet_20v0__lint_diff = -1.7325e-8
+ sky130_fd_pr__nfet_20v0__wint_diff = 3.2175e-8
+ sky130_fd_pr__nfet_20v0__dlc_diff = -1.7325e-8
+ sky130_fd_pr__nfet_20v0__dwc_diff = 3.2175e-8
.param
+ sky130_fd_pr__nfet_20v0__rdrift_mult = 1.8205
+ sky130_fd_pr__nfet_20v0__hvvsat_mult = 1.3172
+ sky130_fd_pr__nfet_20v0__vth0_diff = 1.7977e-1
+ sky130_fd_pr__nfet_20v0__k2_diff = -2.5783e-2
.param
+ sky130_fd_pr__nfet_20v0_iso__rdrift_mult = 2.3846
+ sky130_fd_pr__nfet_20v0_iso__hvvsat_mult = 2.4860
+ sky130_fd_pr__nfet_20v0_iso__vth0_diff = 1.4387e-1
+ sky130_fd_pr__nfet_20v0_iso__k2_diff = -1.9447e-2
.include "sky130_fd_pr__nfet_20v0__subcircuit.pm3.spice"
.include "../nfet_20v0_iso/sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice"
.include "../nfet_20v0_zvt/sky130_fd_pr__nfet_20v0_zvt__fs_discrete.corner.spice"
