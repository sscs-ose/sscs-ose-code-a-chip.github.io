# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.000000 BY  12.50000 ;
  PIN BULK
    ANTENNADIFFAREA  2.929000 ;
    PORT
      LAYER met1 ;
        RECT 0.920000 3.765000 1.210000 8.735000 ;
        RECT 4.785000 3.765000 5.075000 8.735000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  6.262000 ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.000000 6.000000 7.500000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  3.030000 ;
    PORT
      LAYER met1 ;
        RECT 1.700000 3.190000 4.510000 3.480000 ;
        RECT 1.700000 9.020000 4.510000 9.310000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  6.034750 ;
    PORT
      LAYER met3 ;
        RECT 0.000000  0.000000 6.000000  2.500000 ;
        RECT 0.000000 10.000000 6.000000 12.500000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.980000 3.825000 1.150000 8.675000 ;
      RECT 1.535000 3.705000 1.705000 8.795000 ;
      RECT 1.760000 3.250000 4.470000 3.420000 ;
      RECT 1.760000 9.080000 4.470000 9.250000 ;
      RECT 1.955000 3.705000 2.485000 8.795000 ;
      RECT 2.725000 3.705000 3.255000 8.795000 ;
      RECT 3.495000 3.705000 4.025000 8.795000 ;
      RECT 4.275000 3.705000 4.445000 8.795000 ;
      RECT 4.845000 3.825000 5.015000 8.675000 ;
    LAYER mcon ;
      RECT 0.980000 4.185000 1.150000 4.355000 ;
      RECT 0.980000 4.545000 1.150000 4.715000 ;
      RECT 0.980000 4.905000 1.150000 5.075000 ;
      RECT 0.980000 5.265000 1.150000 5.435000 ;
      RECT 0.980000 5.625000 1.150000 5.795000 ;
      RECT 0.980000 5.985000 1.150000 6.155000 ;
      RECT 0.980000 6.345000 1.150000 6.515000 ;
      RECT 0.980000 6.705000 1.150000 6.875000 ;
      RECT 0.980000 7.065000 1.150000 7.235000 ;
      RECT 0.980000 7.425000 1.150000 7.595000 ;
      RECT 0.980000 7.785000 1.150000 7.955000 ;
      RECT 0.980000 8.145000 1.150000 8.315000 ;
      RECT 0.980000 8.505000 1.150000 8.675000 ;
      RECT 1.535000 3.825000 1.705000 3.995000 ;
      RECT 1.535000 4.185000 1.705000 4.355000 ;
      RECT 1.535000 4.545000 1.705000 4.715000 ;
      RECT 1.535000 4.905000 1.705000 5.075000 ;
      RECT 1.535000 5.265000 1.705000 5.435000 ;
      RECT 1.535000 5.625000 1.705000 5.795000 ;
      RECT 1.535000 5.985000 1.705000 6.155000 ;
      RECT 1.535000 6.345000 1.705000 6.515000 ;
      RECT 1.535000 6.705000 1.705000 6.875000 ;
      RECT 1.535000 7.065000 1.705000 7.235000 ;
      RECT 1.535000 7.425000 1.705000 7.595000 ;
      RECT 1.535000 7.785000 1.705000 7.955000 ;
      RECT 1.535000 8.145000 1.705000 8.315000 ;
      RECT 1.535000 8.505000 1.705000 8.675000 ;
      RECT 1.760000 3.250000 1.930000 3.420000 ;
      RECT 1.760000 9.080000 1.930000 9.250000 ;
      RECT 1.955000 3.825000 2.485000 8.675000 ;
      RECT 2.120000 3.250000 2.290000 3.420000 ;
      RECT 2.120000 9.080000 2.290000 9.250000 ;
      RECT 2.480000 3.250000 2.650000 3.420000 ;
      RECT 2.480000 9.080000 2.650000 9.250000 ;
      RECT 2.725000 3.825000 3.255000 8.675000 ;
      RECT 2.840000 3.250000 3.010000 3.420000 ;
      RECT 2.840000 9.080000 3.010000 9.250000 ;
      RECT 3.200000 3.250000 3.370000 3.420000 ;
      RECT 3.200000 9.080000 3.370000 9.250000 ;
      RECT 3.495000 3.825000 4.025000 8.675000 ;
      RECT 3.560000 3.250000 3.730000 3.420000 ;
      RECT 3.560000 9.080000 3.730000 9.250000 ;
      RECT 3.920000 3.250000 4.090000 3.420000 ;
      RECT 3.920000 9.080000 4.090000 9.250000 ;
      RECT 4.275000 3.825000 4.445000 3.995000 ;
      RECT 4.275000 4.185000 4.445000 4.355000 ;
      RECT 4.275000 4.545000 4.445000 4.715000 ;
      RECT 4.275000 4.905000 4.445000 5.075000 ;
      RECT 4.275000 5.265000 4.445000 5.435000 ;
      RECT 4.275000 5.625000 4.445000 5.795000 ;
      RECT 4.275000 5.985000 4.445000 6.155000 ;
      RECT 4.275000 6.345000 4.445000 6.515000 ;
      RECT 4.275000 6.705000 4.445000 6.875000 ;
      RECT 4.275000 7.065000 4.445000 7.235000 ;
      RECT 4.275000 7.425000 4.445000 7.595000 ;
      RECT 4.275000 7.785000 4.445000 7.955000 ;
      RECT 4.275000 8.145000 4.445000 8.315000 ;
      RECT 4.275000 8.505000 4.445000 8.675000 ;
      RECT 4.280000 3.250000 4.450000 3.420000 ;
      RECT 4.280000 9.080000 4.450000 9.250000 ;
      RECT 4.845000 4.185000 5.015000 4.355000 ;
      RECT 4.845000 4.545000 5.015000 4.715000 ;
      RECT 4.845000 4.905000 5.015000 5.075000 ;
      RECT 4.845000 5.265000 5.015000 5.435000 ;
      RECT 4.845000 5.625000 5.015000 5.795000 ;
      RECT 4.845000 5.985000 5.015000 6.155000 ;
      RECT 4.845000 6.345000 5.015000 6.515000 ;
      RECT 4.845000 6.705000 5.015000 6.875000 ;
      RECT 4.845000 7.065000 5.015000 7.235000 ;
      RECT 4.845000 7.425000 5.015000 7.595000 ;
      RECT 4.845000 7.785000 5.015000 7.955000 ;
      RECT 4.845000 8.145000 5.015000 8.315000 ;
      RECT 4.845000 8.505000 5.015000 8.675000 ;
    LAYER met1 ;
      RECT 1.490000 3.620000 1.750000 3.765000 ;
      RECT 1.490000 3.765000 1.765000 8.735000 ;
      RECT 1.490000 8.735000 1.750000 8.880000 ;
      RECT 1.905000 3.765000 2.535000 8.735000 ;
      RECT 2.675000 3.765000 3.305000 8.735000 ;
      RECT 2.700000 3.620000 3.280000 3.765000 ;
      RECT 2.700000 8.735000 3.280000 8.880000 ;
      RECT 3.445000 3.765000 4.075000 8.735000 ;
      RECT 4.215000 3.765000 4.505000 8.735000 ;
      RECT 4.230000 3.620000 4.490000 3.765000 ;
      RECT 4.230000 8.735000 4.490000 8.880000 ;
    LAYER met2 ;
      RECT 0.790000 0.360000 5.210000  4.370000 ;
      RECT 0.790000 4.370000 1.750000  5.220000 ;
      RECT 0.790000 5.220000 1.070000  7.280000 ;
      RECT 0.790000 7.280000 1.750000  8.130000 ;
      RECT 0.790000 8.130000 5.210000 12.140000 ;
      RECT 1.930000 4.650000 2.510000  5.360000 ;
      RECT 1.930000 5.360000 4.050000  7.140000 ;
      RECT 1.930000 7.140000 2.510000  7.850000 ;
      RECT 2.700000 4.370000 3.280000  5.220000 ;
      RECT 2.700000 7.280000 3.280000  8.130000 ;
      RECT 3.470000 4.650000 4.050000  5.360000 ;
      RECT 3.470000 7.140000 4.050000  7.850000 ;
      RECT 4.230000 4.370000 5.210000  5.220000 ;
      RECT 4.230000 7.280000 5.210000  8.130000 ;
      RECT 4.930000 5.220000 5.210000  7.280000 ;
    LAYER via ;
      RECT 1.490000 3.650000 1.750000 3.910000 ;
      RECT 1.490000 3.970000 1.750000 4.230000 ;
      RECT 1.490000 4.290000 1.750000 4.550000 ;
      RECT 1.490000 4.610000 1.750000 4.870000 ;
      RECT 1.490000 4.930000 1.750000 5.190000 ;
      RECT 1.490000 7.310000 1.750000 7.570000 ;
      RECT 1.490000 7.630000 1.750000 7.890000 ;
      RECT 1.490000 7.950000 1.750000 8.210000 ;
      RECT 1.490000 8.270000 1.750000 8.530000 ;
      RECT 1.490000 8.590000 1.750000 8.850000 ;
      RECT 1.930000 4.680000 2.510000 7.820000 ;
      RECT 2.700000 3.650000 3.280000 5.190000 ;
      RECT 2.700000 7.310000 3.280000 8.850000 ;
      RECT 3.470000 4.680000 4.050000 7.820000 ;
      RECT 4.230000 3.650000 4.490000 3.910000 ;
      RECT 4.230000 3.970000 4.490000 4.230000 ;
      RECT 4.230000 4.290000 4.490000 4.550000 ;
      RECT 4.230000 4.610000 4.490000 4.870000 ;
      RECT 4.230000 4.930000 4.490000 5.190000 ;
      RECT 4.230000 7.310000 4.490000 7.570000 ;
      RECT 4.230000 7.630000 4.490000 7.890000 ;
      RECT 4.230000 7.950000 4.490000 8.210000 ;
      RECT 4.230000 8.270000 4.490000 8.530000 ;
      RECT 4.230000 8.590000 4.490000 8.850000 ;
    LAYER via2 ;
      RECT 2.350000  0.610000 3.630000  1.890000 ;
      RECT 2.350000  5.610000 3.630000  6.890000 ;
      RECT 2.350000 10.610000 3.630000 11.890000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15
END LIBRARY
