* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 40
.param
+ sky130_fd_pr__pfet_01v8_lvt__toxe_mult = 1.0365
+ sky130_fd_pr__pfet_01v8_lvt__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8_lvt__overlap_mult = 0.1
+ sky130_fd_pr__pfet_01v8_lvt__ajunction_mult = 1.0625e+0
+ sky130_fd_pr__pfet_01v8_lvt__pjunction_mult = 1.0675e+0
+ sky130_fd_pr__pfet_01v8_lvt__lint_diff = -1.21275e-8
+ sky130_fd_pr__pfet_01v8_lvt__wint_diff = 2.252e-8
+ sky130_fd_pr__pfet_01v8_lvt__dlc_diff = -5.0625e-8
+ sky130_fd_pr__pfet_01v8_lvt__dwc_diff = 2.252e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 000, W = 1.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_0 = -7.9865e-5
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_0 = 0.26574
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0 = -0.12644
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_0 = 0.013397
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_0 = -0.031262
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 001, W = 1.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_1 = -0.026236
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_1 = -0.00012786
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_1 = 0.16579
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1 = -0.078037
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_1 = 0.081181
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 002, W = 1.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_2 = 0.081703
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_2 = -0.020702
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_2 = -0.00022389
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_2 = 0.183
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2 = -0.077468
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 003, W = 1.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_3 = 0.045553
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_3 = -0.031278
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_3 = -0.00011891
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_3 = 0.25821
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3 = -0.098522
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 004, W = 1.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4 = -0.21233
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_4 = -4.0845e-7
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_4 = -0.055821
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_4 = -0.00010561
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4 = 22877.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_4 = 2.0229e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 005, W = 1.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5 = -0.14333
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_5 = -3.3163e-7
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_5 = -0.03971
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_5 = -4.1155e-6
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5 = -16718.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_5 = 2.0889e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 006, W = 3.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_6 = 0.31235
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6 = -0.12188
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_6 = 0.0033223
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_6 = -0.028586
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_6 = -0.00010427
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_6 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 007, W = 3.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_7 = 0.28274
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7 = -0.11161
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_7 = 0.050471
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_7 = -0.041535
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_7 = 2.937e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 008, W = 3.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_8 = 0.24672
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8 = -0.10446
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_8 = 0.048259
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_8 = -0.028313
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_8 = -9.7474e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 009, W = 3.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_9 = 0.23037
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9 = -0.11028
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_9 = 0.06987
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_9 = -0.02342
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_9 = -0.0001049
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 010, W = 3.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_10 = -4.5499e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10 = -0.09476
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_10 = -0.024151
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_10 = 0.14637
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_10 = 0.10102
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 011, W = 3.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_11 = -7.0217e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11 = 23349.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11 = -0.13201
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_11 = -0.022
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_11 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 012, W = 3.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_12 = -0.020745
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_12 = 0.067887
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_12 = -0.00020593
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12 = -2327.4
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12 = -0.1054
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_12 = -1.5721e-6
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_12 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 013, W = 5.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_13 = -0.029978
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_13 = 0.15367
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_13 = 0.1035
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_13 = 3.1431e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13 = -0.11225
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 014, W = 5.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_14 = -0.027419
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_14 = 0.14457
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_14 = 0.09664
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_14 = 9.0274e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14 = -0.10521
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 015, W = 5.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_15 = -0.032015
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_15 = 0.19313
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_15 = 0.0963
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_15 = 0.00015852
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15 = -0.13808
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 016, W = 5.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_16 = -0.031826
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_16 = 0.10669
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_16 = 0.11957
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_16 = 5.5834e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16 = -0.11322
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 017, W = 5.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_17 = -0.024784
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_17 = 0.11407
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_17 = 0.11413
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_17 = 2.3472e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17 = -0.10164
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 018, W = 5.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_18 = -0.023553
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_18 = -0.00012549
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18 = 42777.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18 = -0.14765
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 019, W = 5.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_19 = -2.1376e-6
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_19 = -0.025587
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_19 = 0.026955
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_19 = 7.7099e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19 = -4093.1
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19 = -0.14239
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 020, W = 7.0, L = 1.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_20 = -0.03401
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_20 = 0.22865
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_20 = 0.01776
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_20 = 9.2552e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20 = -0.12381
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 021, W = 7.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_21 = 8.4983e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21 = -0.12337
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_21 = -0.042648
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_21 = 0.31403
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_21 = 0.044806
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 022, W = 7.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_22 = 0.25061
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_22 = 0.051013
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_22 = 0.00011455
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22 = -0.12704
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_22 = -0.049808
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_22 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 023, W = 7.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_23 = -0.027279
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_23 = 0.07464
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_23 = 0.12836
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_23 = 0.00012004
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23 = -0.11276
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_23 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 024, W = 7.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_24 = -0.027321
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_24 = 0.095877
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_24 = 0.11944
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_24 = 0.00014347
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24 = -0.12483
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 025, W = 7.0, L = 0.35
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_25 = -0.02542
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_25 = 6.1758e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25 = 15561.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25 = -0.15314
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 026, W = 7.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_26 = -0.028935
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_26 = 0.040782
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_26 = 1.7596e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26 = 30959.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26 = -0.11716
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_26 = -1.3309e-6
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 027, W = 0.42, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_27 = -3.5263e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_27 = 4.9834e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_27 = -0.053258
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_27 = 0.00037297
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27 = -0.18802
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 028, W = 0.42, L = 20.0
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_28 = -1.3381e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_28 = 2.0394e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_28 = -0.0209
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_28 = -0.00013203
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28 = -0.039406
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 029, W = 0.42, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_29 = -1.645e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_29 = 2.3047e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_29 = -0.03151
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_29 = -7.8723e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29 = -0.083464
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 030, W = 0.42, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_30 = -1.5578e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_30 = 2.0496e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_30 = -0.03191
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_30 = 8.7575e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30 = -0.1002
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_30 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 031, W = 0.42, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_31 = -1.0904e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_31 = 2.0176e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_31 = -0.030874
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_31 = -2.7331e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31 = -0.076934
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 032, W = 0.42, L = 0.35
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_32 = -0.00022831
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32 = 22176.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32 = -0.028993
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_32 = -0.021402
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 033, W = 0.42, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_33 = -3.7451e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33 = -16660.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33 = -0.1555
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_33 = -3.2745e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_33 = 2.075e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_33 = -0.045013
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_33 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 034, W = 0.55, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_34 = -0.03876
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_34 = -5.9923e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34 = -0.09247
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_34 = -2.1647e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_34 = 4.5689e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_34 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 035, W = 0.55, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_35 = -0.014723
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_35 = -2.2899e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35 = -0.099678
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_35 = -2.0612e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_35 = 2.0168e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 036, W = 0.55, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_36 = -0.018294
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_36 = -3.6145e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36 = -0.10614
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_36 = -3.745e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_36 = 1.9928e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 037, W = 0.55, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_37 = 2.0388e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_37 = -0.012579
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_37 = 1.3378e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37 = -0.083362
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_37 = -1.7748e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 038, W = 0.55, L = 0.35
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_38 = -0.037031
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_38 = -0.0001037
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38 = 46735.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38 = -0.18084
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 039, W = 0.55, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_39 = -4.3799e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_39 = 4.8359e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_39 = -0.054464
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_39 = 0.00041255
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39 = -11942.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39 = -0.23487
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_39 = 0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"
