module approxMult_signed8x8 (A, B, OUT);
  input  [7:0] A;
  input  [7:0] B;
  output [15:0] OUT;
  wire n10, n11, n12, n13, n14, n15, n2, n3, n4, n5, n6, n7, n8, v0_0, v100_0, v101_0, v102_0, v103_0, v104_0, v105_0, v106_0, v107_0, v108_0, v109_0, v10_0, v110_0, v111_0, v112_0, v113_0, v114_0, v115_0, v116_0, v117_0, v118_0, v119_0, v11_0, v120_0, v121_0, v122_0, v123_0, v124_0, v125_0, v126_0, v127_0, v128_0, v129_0, v12_0, v130_0, v131_0, v132_0, v133_0, v134_0, v135_0, v136_0, v137_0, v138_0, v139_0, v13_0, v140_0, v141_0, v142_0, v143_0, v144_0, v145_0, v146_0, v147_0, v148_0, v149_0, v14_0, v150_0, v151_0, v152_0, v153_0, v154_0, v155_0, v156_0, v157_0, v158_0, v159_0, v15_0, v160_0, v161_0, v162_0, v163_0, v164_0, v165_0, v166_0, v167_0, v168_0, v169_0, v16_0, v170_0, v171_0, v172_0, v173_0, v174_0, v175_0, v176_0, v177_0, v178_0, v179_0, v17_0, v180_0, v181_0, v182_0, v183_0, v184_0, v185_0, v186_0, v187_0, v188_0, v18_0, v19_0, v1_0, v20_0, v21_0, v22_0, v23_0, v24_0, v25_0, v26_0, v27_0, v28_0, v29_0, v2_0, v30_0, v31_0, v32_0, v33_0, v34_0, v35_0, v36_0, v37_0, v38_0, v39_0, v3_0, v40_0, v41_0, v42_0, v43_0, v44_0, v45_0, v46_0, v47_0, v48_0, v49_0, v4_0, v50_0, v51_0, v52_0, v53_0, v54_0, v55_0, v56_0, v57_0, v58_0, v59_0, v5_0, v60_0, v61_0, v62_0, v63_0, v64_0, v65_0, v66_0, v67_0, v68_0, v69_0, v6_0, v70_0, v71_0, v72_0, v73_0, v74_0, v75_0, v76_0, v77_0, v78_0, v79_0, v7_0, v80_0, v81_0, v82_0, v83_0, v84_0, v85_0, v86_0, v87_0, v88_0, v89_0, v8_0, v90_0, v91_0, v92_0, v93_0, v94_0, v95_0, v96_0, v97_0, v98_0, v99_0, v9_0;

  // Map n0..n7 to A[0..7], n8..n15 to B[0..7]
  assign n0 = A[0];
  assign n1 = A[1];
  assign n2 = A[2];
  assign n3 = A[3];
  assign n4 = A[4];
  assign n5 = A[5];
  assign n6 = A[6];
  assign n7 = A[7];
  assign n8 = B[0];
  assign n9 = B[1];
  assign n10 = B[2];
  assign n11 = B[3];
  assign n12 = B[4];
  assign n13 = B[5];
  assign n14 = B[6];
  assign n15 = B[7];

  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0001_ (
    .I(n2),
    .ZN(v0_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0002_ (
    .A1(n12),
    .A2(n5),
    .ZN(v1_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0003_ (
    .I(n4),
    .ZN(v2_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0004_ (
    .I(n15),
    .ZN(v3_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0005_ (
    .A1(n5),
    .A2(n11),
    .ZN(v4_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0006_ (
    .A1(v2_0),
    .A2(v1_0),
    .Z(v5_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0007_ (
    .I(n7),
    .ZN(v6_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0008_ (
    .I(n3),
    .ZN(v7_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0009_ (
    .A1(v3_0),
    .A2(v7_0),
    .Z(v8_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0010_ (
    .I(v8_0),
    .ZN(v9_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0011_ (
    .I(n11),
    .ZN(v10_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0012_ (
    .A1(v0_0),
    .A2(v3_0),
    .ZN(v11_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0013_ (
    .A1(n11),
    .A2(n6),
    .ZN(v12_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0014_ (
    .A1(v1_0),
    .A2(v12_0),
    .ZN(v13_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0015_ (
    .I(v13_0),
    .ZN(v14_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0016_ (
    .A1(n4),
    .A2(n13),
    .ZN(v15_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0017_ (
    .A1(v14_0),
    .A2(v15_0),
    .Z(v16_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0018_ (
    .A1(v14_0),
    .A2(v15_0),
    .ZN(v17_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0019_ (
    .I(v6_0),
    .ZN(v18_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0020_ (
    .I(v5_0),
    .ZN(v19_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0021_ (
    .A1(n11),
    .A2(v19_0),
    .Z(v20_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0022_ (
    .A1(v6_0),
    .A2(n10),
    .Z(v21_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0023_ (
    .A1(v10_0),
    .A2(v21_0),
    .Z(v22_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0024_ (
    .A1(n3),
    .A2(v3_0),
    .ZN(v23_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0025_ (
    .I(v23_0),
    .ZN(v24_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0026_ (
    .A1(v22_0),
    .A2(v24_0),
    .Z(v25_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0027_ (
    .A1(v22_0),
    .A2(v24_0),
    .ZN(v26_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0028_ (
    .A1(v25_0),
    .A2(v26_0),
    .Z(v27_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0029_ (
    .A1(v27_0),
    .A2(v9_0),
    .Z(v28_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0030_ (
    .A1(v22_0),
    .A2(v10_0),
    .Z(v29_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0031_ (
    .I(v29_0),
    .ZN(v30_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0032_ (
    .A1(v19_0),
    .A2(n14),
    .ZN(v31_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0033_ (
    .I(v31_0),
    .ZN(v32_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0034_ (
    .A1(n4),
    .A2(n14),
    .ZN(v33_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0035_ (
    .A1(v8_0),
    .A2(n15),
    .ZN(v34_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0036_ (
    .A1(v33_0),
    .A2(v34_0),
    .Z(v35_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0037_ (
    .A1(n12),
    .A2(n6),
    .ZN(v36_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0038_ (
    .A1(v4_0),
    .A2(v36_0),
    .Z(v37_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0039_ (
    .A1(v16_0),
    .A2(v37_0),
    .ZN(v38_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0040_ (
    .A1(v35_0),
    .A2(v38_0),
    .Z(v39_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0041_ (
    .I(v39_0),
    .ZN(v40_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0042_ (
    .A1(n11),
    .A2(n7),
    .ZN(v41_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0043_ (
    .A1(v36_0),
    .A2(v41_0),
    .Z(v42_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0044_ (
    .I(v42_0),
    .ZN(v43_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0045_ (
    .A1(n5),
    .A2(n13),
    .ZN(v44_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0046_ (
    .A1(v43_0),
    .A2(v44_0),
    .Z(v45_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0047_ (
    .A1(v43_0),
    .A2(v44_0),
    .ZN(v46_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0048_ (
    .A1(v45_0),
    .A2(v46_0),
    .Z(v47_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0049_ (
    .I(v47_0),
    .ZN(v48_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0050_ (
    .A1(v6_0),
    .A2(v48_0),
    .Z(v49_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0051_ (
    .I(v49_0),
    .ZN(v50_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0052_ (
    .A1(v40_0),
    .A2(v50_0),
    .Z(v51_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0053_ (
    .A1(v17_0),
    .A2(v11_0),
    .ZN(v52_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0054_ (
    .A1(v20_0),
    .A2(v52_0),
    .ZN(v53_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0055_ (
    .A1(v51_0),
    .A2(v53_0),
    .Z(v54_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0056_ (
    .A1(v32_0),
    .A2(v54_0),
    .Z(v55_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0057_ (
    .A1(v30_0),
    .A2(v55_0),
    .Z(v56_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0058_ (
    .I(v28_0),
    .ZN(v57_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0059_ (
    .A1(v57_0),
    .A2(v25_0),
    .ZN(v58_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0060_ (
    .I(v58_0),
    .ZN(v59_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0061_ (
    .A1(v56_0),
    .A2(v59_0),
    .Z(v60_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0062_ (
    .A1(v38_0),
    .A2(v35_0),
    .ZN(v61_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0063_ (
    .I(v61_0),
    .ZN(v62_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0064_ (
    .A1(v50_0),
    .A2(v40_0),
    .Z(v63_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0065_ (
    .I(v63_0),
    .ZN(v64_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0066_ (
    .A1(n5),
    .A2(n14),
    .ZN(v65_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0067_ (
    .A1(v2_0),
    .A2(n15),
    .ZN(v66_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0068_ (
    .A1(v65_0),
    .A2(v66_0),
    .Z(v67_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0069_ (
    .A1(v36_0),
    .A2(v42_0),
    .Z(v68_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0070_ (
    .A1(v45_0),
    .A2(v68_0),
    .ZN(v69_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0071_ (
    .A1(v67_0),
    .A2(v69_0),
    .Z(v70_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0072_ (
    .I(v70_0),
    .ZN(v71_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0073_ (
    .A1(v34_0),
    .A2(v33_0),
    .Z(v72_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0074_ (
    .A1(v71_0),
    .A2(v72_0),
    .Z(v73_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0075_ (
    .A1(v71_0),
    .A2(v72_0),
    .ZN(v74_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0076_ (
    .A1(v73_0),
    .A2(v74_0),
    .Z(v75_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0077_ (
    .A1(v18_0),
    .A2(v47_0),
    .ZN(v76_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0078_ (
    .I(v76_0),
    .ZN(v77_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0079_ (
    .I(v41_0),
    .ZN(v78_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0080_ (
    .A1(v78_0),
    .A2(n12),
    .ZN(v79_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0081_ (
    .A1(n12),
    .A2(n7),
    .ZN(v80_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0082_ (
    .A1(v41_0),
    .A2(v80_0),
    .ZN(v81_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0083_ (
    .A1(v79_0),
    .A2(v81_0),
    .ZN(v82_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0084_ (
    .A1(n13),
    .A2(n6),
    .ZN(v83_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0085_ (
    .A1(v82_0),
    .A2(v83_0),
    .Z(v84_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0086_ (
    .A1(v82_0),
    .A2(v83_0),
    .ZN(v85_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0087_ (
    .A1(v84_0),
    .A2(v85_0),
    .Z(v86_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0088_ (
    .I(v86_0),
    .ZN(v87_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0089_ (
    .A1(v87_0),
    .A2(v6_0),
    .Z(v88_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0090_ (
    .A1(v77_0),
    .A2(v88_0),
    .Z(v89_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0091_ (
    .A1(v77_0),
    .A2(v87_0),
    .ZN(v90_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0092_ (
    .A1(v89_0),
    .A2(v90_0),
    .Z(v91_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0093_ (
    .A1(v75_0),
    .A2(v91_0),
    .Z(v92_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0094_ (
    .A1(v64_0),
    .A2(v92_0),
    .Z(v93_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0095_ (
    .A1(v62_0),
    .A2(v93_0),
    .Z(v94_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0096_ (
    .A1(v54_0),
    .A2(v32_0),
    .ZN(v95_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0097_ (
    .A1(v53_0),
    .A2(v51_0),
    .ZN(v96_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0098_ (
    .A1(v95_0),
    .A2(v96_0),
    .ZN(v97_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0099_ (
    .A1(v94_0),
    .A2(v97_0),
    .Z(v98_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0100_ (
    .A1(v94_0),
    .A2(v97_0),
    .ZN(v99_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0101_ (
    .A1(v98_0),
    .A2(v99_0),
    .Z(v100_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0102_ (
    .A1(v59_0),
    .A2(v56_0),
    .ZN(v101_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0103_ (
    .A1(v55_0),
    .A2(v30_0),
    .ZN(v102_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0104_ (
    .A1(v101_0),
    .A2(v102_0),
    .ZN(v103_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0105_ (
    .A1(v100_0),
    .A2(v103_0),
    .Z(v104_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0106_ (
    .A1(v93_0),
    .A2(v62_0),
    .ZN(v105_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0107_ (
    .A1(v92_0),
    .A2(v64_0),
    .ZN(v106_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0108_ (
    .A1(v105_0),
    .A2(v106_0),
    .ZN(v107_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0109_ (
    .A1(v69_0),
    .A2(v71_0),
    .ZN(v108_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0110_ (
    .A1(v73_0),
    .A2(v108_0),
    .ZN(v109_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0111_ (
    .A1(v91_0),
    .A2(v75_0),
    .ZN(v110_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0112_ (
    .A1(v110_0),
    .A2(v90_0),
    .ZN(v111_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0113_ (
    .A1(n6),
    .A2(n14),
    .ZN(v112_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0114_ (
    .I(n5),
    .ZN(v113_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0115_ (
    .A1(v113_0),
    .A2(n15),
    .ZN(v114_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0116_ (
    .A1(v112_0),
    .A2(v114_0),
    .Z(v115_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0117_ (
    .A1(v84_0),
    .A2(v79_0),
    .ZN(v116_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0118_ (
    .A1(v115_0),
    .A2(v116_0),
    .Z(v117_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0119_ (
    .I(v117_0),
    .ZN(v118_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0120_ (
    .A1(v66_0),
    .A2(v65_0),
    .Z(v119_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0121_ (
    .A1(v118_0),
    .A2(v119_0),
    .Z(v120_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0122_ (
    .A1(v118_0),
    .A2(v119_0),
    .ZN(v121_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0123_ (
    .A1(v120_0),
    .A2(v121_0),
    .Z(v122_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0124_ (
    .A1(v18_0),
    .A2(v86_0),
    .ZN(v123_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0125_ (
    .I(v123_0),
    .ZN(v124_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0126_ (
    .A1(n13),
    .A2(n7),
    .ZN(v125_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0127_ (
    .A1(v125_0),
    .A2(v82_0),
    .Z(v126_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0128_ (
    .I(v126_0),
    .ZN(v127_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0129_ (
    .A1(v127_0),
    .A2(v6_0),
    .Z(v128_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0130_ (
    .A1(v124_0),
    .A2(v128_0),
    .Z(v129_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0131_ (
    .A1(v124_0),
    .A2(v127_0),
    .ZN(v130_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0132_ (
    .A1(v129_0),
    .A2(v130_0),
    .Z(v131_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0133_ (
    .A1(v122_0),
    .A2(v131_0),
    .Z(v132_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0134_ (
    .A1(v111_0),
    .A2(v132_0),
    .Z(v133_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0135_ (
    .A1(v109_0),
    .A2(v133_0),
    .Z(v134_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0136_ (
    .A1(v107_0),
    .A2(v134_0),
    .Z(v135_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0137_ (
    .A1(v104_0),
    .A2(v99_0),
    .Z(v136_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0138_ (
    .I(v136_0),
    .ZN(v137_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0139_ (
    .A1(v137_0),
    .A2(v98_0),
    .Z(v138_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0140_ (
    .A1(v135_0),
    .A2(v138_0),
    .Z(v139_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0141_ (
    .A1(v116_0),
    .A2(v115_0),
    .ZN(v140_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0142_ (
    .A1(v120_0),
    .A2(v140_0),
    .ZN(v141_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0143_ (
    .A1(v131_0),
    .A2(v122_0),
    .ZN(v142_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0144_ (
    .A1(v142_0),
    .A2(v130_0),
    .ZN(v143_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0145_ (
    .A1(v82_0),
    .A2(v125_0),
    .Z(v144_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0146_ (
    .A1(v144_0),
    .A2(v79_0),
    .ZN(v145_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0147_ (
    .I(v145_0),
    .ZN(v146_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0148_ (
    .A1(n14),
    .A2(v18_0),
    .ZN(v147_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0149_ (
    .I(v147_0),
    .ZN(v148_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0150_ (
    .A1(v3_0),
    .A2(n6),
    .Z(v149_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0151_ (
    .A1(v148_0),
    .A2(v149_0),
    .Z(v150_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0152_ (
    .A1(v146_0),
    .A2(v150_0),
    .Z(v151_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0153_ (
    .A1(v146_0),
    .A2(v150_0),
    .ZN(v152_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0154_ (
    .A1(v151_0),
    .A2(v152_0),
    .Z(v153_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0155_ (
    .I(v153_0),
    .ZN(v154_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0156_ (
    .A1(v115_0),
    .A2(v112_0),
    .Z(v155_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0157_ (
    .A1(v154_0),
    .A2(v155_0),
    .Z(v156_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0158_ (
    .A1(v154_0),
    .A2(v155_0),
    .ZN(v157_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0159_ (
    .A1(v156_0),
    .A2(v157_0),
    .Z(v158_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0160_ (
    .A1(v18_0),
    .A2(v158_0),
    .Z(v159_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0161_ (
    .A1(v143_0),
    .A2(v159_0),
    .Z(v160_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0162_ (
    .A1(v141_0),
    .A2(v160_0),
    .Z(v161_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0163_ (
    .A1(v133_0),
    .A2(v109_0),
    .ZN(v162_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0164_ (
    .A1(v132_0),
    .A2(v111_0),
    .ZN(v163_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0165_ (
    .A1(v162_0),
    .A2(v163_0),
    .ZN(v164_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0166_ (
    .A1(v161_0),
    .A2(v164_0),
    .Z(v165_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0167_ (
    .A1(v161_0),
    .A2(v164_0),
    .ZN(v166_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__and2_1 _0168_ (
    .A1(v165_0),
    .A2(v166_0),
    .Z(v167_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0169_ (
    .A1(v138_0),
    .A2(v135_0),
    .ZN(v168_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0170_ (
    .A1(v134_0),
    .A2(v107_0),
    .ZN(v169_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0171_ (
    .A1(v168_0),
    .A2(v169_0),
    .ZN(v170_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0172_ (
    .A1(v167_0),
    .A2(v170_0),
    .Z(v171_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0173_ (
    .A1(v156_0),
    .A2(v151_0),
    .ZN(v172_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0174_ (
    .A1(v149_0),
    .A2(v148_0),
    .ZN(v173_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__or2_1 _0175_ (
    .A1(v3_0),
    .A2(n7),
    .Z(v174_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0176_ (
    .A1(v173_0),
    .A2(v174_0),
    .ZN(v175_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0177_ (
    .A1(v175_0),
    .A2(v145_0),
    .Z(v176_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0178_ (
    .A1(v176_0),
    .A2(v18_0),
    .Z(v177_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0179_ (
    .A1(v158_0),
    .A2(v18_0),
    .ZN(v178_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__inv_1 _0180_ (
    .I(v178_0),
    .ZN(v179_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0181_ (
    .A1(v177_0),
    .A2(v179_0),
    .Z(v180_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0182_ (
    .A1(v172_0),
    .A2(v180_0),
    .Z(v181_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0183_ (
    .A1(v160_0),
    .A2(v141_0),
    .ZN(v182_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0184_ (
    .A1(v159_0),
    .A2(v143_0),
    .ZN(v183_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0185_ (
    .A1(v182_0),
    .A2(v183_0),
    .ZN(v184_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0186_ (
    .A1(v181_0),
    .A2(v184_0),
    .Z(v185_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0187_ (
    .A1(v170_0),
    .A2(v165_0),
    .ZN(v186_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__nand2_1 _0188_ (
    .A1(v186_0),
    .A2(v166_0),
    .ZN(v187_0)
  );
  gf180mcu_fd_sc_mcu9t5v0__xor2_1 _0189_ (
    .A1(v185_0),
    .A2(v187_0),
    .Z(v188_0)
  );

  assign OUT[0] = v42_0;
  assign OUT[1] = n8;
  assign OUT[2] = v112_0;
  assign OUT[3] = v157_0;
  assign OUT[4] = v141_0;
  assign OUT[5] = v115_0;
  assign OUT[6] = v85_0;
  assign OUT[7] = n10;
  assign OUT[8] = v116_0;
  assign OUT[9] = v28_0;
  assign OUT[10] = v60_0;
  assign OUT[11] = v104_0;
  assign OUT[12] = v139_0;
  assign OUT[13] = v171_0;
  assign OUT[14] = v188_0;
  assign OUT[15] = v188_0;
endmodule
