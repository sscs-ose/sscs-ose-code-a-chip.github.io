** MIYAHARA flat netlist
M2 NET1 VIN+ NET3 M2N7002 M=1
M4 GND CLK NET1 M2N7002 M=1
M5 NET1 VIN- NET2 M2N7002 M=1
M1 NET1 VB NET2 M2N7002 M=1
M3 NET1 VCH NET3 M2N7002 M=1
M6 GND NET2 NET4 M2N7002 M=1
M7 GND NET5 NET4 M2N7002 M=1
M8 GND NET4 NET5 M2N7002 M=1
M9 GND NET3 NET5 M2N7002 M=1
M10 GND NET2 NET6 M2N7002 M=1
M11 GND NET3 NET7 M2N7002 M=1
M12 NET5 NET4 NET7 DMP2035U M=1
M13 NET6 NET2 VDD DMP2035U M=1
M14 NET4 NET5 NET6 DMP2035U M=1
M15 NET7 NET3 VDD DMP2035U M=1
M16 NET2 CLK VDD DMP2035U M=1
M17 NET3 CLK VDD DMP2035U M=1
.end
