# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  1.470000 BY  4.120000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.840000 ;
    PORT
      LAYER met2 ;
        RECT 0.605000 2.440000 0.865000 3.080000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.900000 ;
    PORT
      LAYER met1 ;
        RECT 0.410000 3.365000 1.060000 3.655000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.590000 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.445000 1.280000 -0.145000 ;
        RECT 0.190000 -0.145000 0.420000  3.105000 ;
        RECT 1.050000 -0.145000 1.280000  3.105000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.235000 0.390000 3.105000 ;
      RECT 0.400000 3.335000 1.070000 3.675000 ;
      RECT 0.650000 0.255000 0.820000 3.105000 ;
      RECT 1.080000 0.255000 1.250000 3.105000 ;
    LAYER mcon ;
      RECT 0.220000 0.335000 0.390000 0.505000 ;
      RECT 0.220000 0.695000 0.390000 0.865000 ;
      RECT 0.220000 1.055000 0.390000 1.225000 ;
      RECT 0.220000 1.415000 0.390000 1.585000 ;
      RECT 0.220000 1.775000 0.390000 1.945000 ;
      RECT 0.220000 2.135000 0.390000 2.305000 ;
      RECT 0.220000 2.495000 0.390000 2.665000 ;
      RECT 0.220000 2.855000 0.390000 3.025000 ;
      RECT 0.470000 3.425000 0.640000 3.595000 ;
      RECT 0.650000 0.335000 0.820000 0.505000 ;
      RECT 0.650000 0.695000 0.820000 0.865000 ;
      RECT 0.650000 1.055000 0.820000 1.225000 ;
      RECT 0.650000 1.415000 0.820000 1.585000 ;
      RECT 0.650000 1.775000 0.820000 1.945000 ;
      RECT 0.650000 2.135000 0.820000 2.305000 ;
      RECT 0.650000 2.495000 0.820000 2.665000 ;
      RECT 0.650000 2.855000 0.820000 3.025000 ;
      RECT 0.830000 3.425000 1.000000 3.595000 ;
      RECT 1.080000 0.335000 1.250000 0.505000 ;
      RECT 1.080000 0.695000 1.250000 0.865000 ;
      RECT 1.080000 1.055000 1.250000 1.225000 ;
      RECT 1.080000 1.415000 1.250000 1.585000 ;
      RECT 1.080000 1.775000 1.250000 1.945000 ;
      RECT 1.080000 2.135000 1.250000 2.305000 ;
      RECT 1.080000 2.495000 1.250000 2.665000 ;
      RECT 1.080000 2.855000 1.250000 3.025000 ;
    LAYER met1 ;
      RECT 0.605000 0.255000 0.865000 3.105000 ;
    LAYER via ;
      RECT 0.605000 2.470000 0.865000 2.730000 ;
      RECT 0.605000 2.790000 0.865000 3.050000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15
END LIBRARY
