* SKY130 Spice File.
* Number of bins: 1
* 9 parameters
.param
+ sky130_fd_bs_flash__special_sonosfet_star__tox_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__overlap_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__lint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__wint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__dlc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__dwc_diff = 0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 000, W = 0.45, L = 0.22
* ------------------------------------
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0 = -1.3147e-1
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0 = 7.1682e-3
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0 = -4.1163e-1
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0 = 0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 001, W = 1.00, L = 0.50
* ------------------------------------
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_1 = 2.6332e-1
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_1 = -3.4880e-1
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_1 = -1.7269e-3
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_1 = 0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 002, W = 0.35, L = 0.15
* ------------------------------------
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_2 = -2.6498e-1
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_2 = -5.2454e-3
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_2 = -6.6727e-1
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_2 = 0.0
