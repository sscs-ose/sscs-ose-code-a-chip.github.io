* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p15 BULK DRAIN GATE SOURCE
X0 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u
X1 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u
X2 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u
X3 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u
.ends
