** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/tb_cm_ota_working_v2_extracted.sch
**.subckt tb_cm_ota_working_v2_extracted
V1 vdd GND 1.8
C1 out GND 4p m=1
V3 inn GND DC 1
V4 inp GND DC 1 AC 1
X1 vdd out inp inn itail GND cm_ota w1_2=1.13 w3_4=4.23 w5_6=11.67 w7_8=43.77 w9_10=2.26 beta=1 nf1_2=1 nf3_4=1 nf5_6=1 nf7_8=1
+ nf9_10=1
I3 GND itail 22u

V123 avdd_1v8_ext GND 1.8
C123 out_ext GND 4p m=1
V323 inn_ext GND DC 1 AC 1
V423 inp_ext GND 1
X123 iref_ext out_ext inn_ext inp_ext GND avdd_1v8_ext cm_ota_extracted
I123 GND iref_ext 35.2u



**** begin user architecture code

** opencircuitdesign pdks isntsall
.lib /opt/pdk/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.temp 27
.option savecurrents
.save all
.control
	op
	print I(V1)       ; Print the current through voltage source V1
	print I(V123)
	ac dec 10 1 1e15
	set filetype=ascii
	wrdata ac_output.txt frequency vdb(out) cph(out)
	wrdata ac_phase_output.txt frequency cph(out)
	wrdata ac_output_ext.txt frequency vdb(out_ext) cph(out_ext)
	wrdata ac_phase_output_ext.txt frequency cph(out_ext)
	plot vdb(out) vs frequency
	plot (180*cph(out)/pi) vs frequency
	let phase_vector = 180*cph(out)/pi
	let gain_vector = vdb(out)
	let phase_vector_ext = 180*cph(out_ext)/pi
	let gain_vector_ext = vdb(out_ext)
	meas ac unity_gain_freq_val when vdb(out)=0
	meas ac dc_gain_val find vdb(out) at=10Hz
	meas ac unity_gain_freq_val_ext when vdb(out_ext)=0
	meas ac dc_gain_val find vdb(out_ext) at=10Hz
	let dc_gain = dc_gain_val
	meas ac p1_val when phase_vector=-45 cross=1
	meas ac p2_val when phase_vector=-135 cross=1
	meas ac p1_val_ext when phase_vector_ext=-45 cross=1
	meas ac p2_val_ext when phase_vector_ext=-135 cross=1
	meas ac three_db when gain_vector=dc_gain_val -3 cross=1
	let p2 = p2_val
	let p1 = p1_val
	let dc_gain = dc_gain_val
	let unity_gain_freq = unity_gain_freq_val
	op
	print I(V1)       ; Print the current through voltage source V1
	print I(V123)
	write tb_cm_ota_working_v2_extracted_ac.raw

	let gm1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8[gm]
	let gm2 = @m.x1.xm2.msky130_fd_pr__nfet_01v8[gm]
	let gm3 = @m.x1.xm3.msky130_fd_pr__pfet_01v8[gm]
	let gm4 = @m.x1.xm4.msky130_fd_pr__pfet_01v8[gm]
	let gm5 = @m.x1.xm5.msky130_fd_pr__nfet_01v8[gm]
	let gm6 = @m.x1.xm6.msky130_fd_pr__nfet_01v8[gm]
	let gm7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8[gm]
	let gm8 = @m.x1.xm8.msky130_fd_pr__pfet_01v8[gm]

	let id1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8[id]
	let id2 = @m.x1.xm2.msky130_fd_pr__nfet_01v8[id]
	let id3 = @m.x1.xm3.msky130_fd_pr__pfet_01v8[id]
	let id4 = @m.x1.xm4.msky130_fd_pr__pfet_01v8[id]
	let id5 = @m.x1.xm5.msky130_fd_pr__nfet_01v8[id]
	let id6 = @m.x1.xm6.msky130_fd_pr__nfet_01v8[id]
	let id7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8[id]
	let id8 = @m.x1.xm8.msky130_fd_pr__pfet_01v8[id]

	let current_scale = id5/id1

	let kgm1 = gm1/id1
	let kgm2 = gm2/id2
	let kgm3 = gm3/id3
	let kgm4 = gm4/id4
	let kgm5 = gm5/id5
	let kgm6 = gm6/id6
	let kgm7 = gm7/id7
	let kgm8 = gm8/id8

	print kgm1
	print kgm2
	print kgm3
	print kgm4
	print kgm5
	print kgm6
	print kgm7
	print kgm8

	print id1
	print id2
	print id3
	print id4
	print id5
	print id6
	print id7
	print id8

	print current_scale
	print dc_gain_val
	print p1_val
	print p2_val
.endc


**** end user architecture code
**.ends

* expanding   symbol:  cm_ota.sym # of pins=6
** sym_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sym
** sch_path: /home/adair/Documents/CAD/xschem_library_adair/schematics/cm_ota.sch
.subckt cm_ota vdd out inp inn itail vss  w1_2=1 w3_4=1 w5_6=1 w7_8=1 w9_10=1 beta=2 nf1_2=2 nf3_4=2 nf5_6=2 nf7_8=2 nf9_10=2
*.iopin inn
*.iopin inp
*.iopin out
*.iopin vss
*.iopin vdd
*.iopin itail
XM1 ds1_3 inn source source sky130_fd_pr__nfet_01v8 L=0.500 W=w1_2 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM3 ds1_3 ds1_3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.500 W=w3_4 nf=nf3_4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 ds2_4 inp source source sky130_fd_pr__nfet_01v8 L=0.500 W=w1_2 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM4 ds2_4 ds2_4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.500 W=w3_4 nf=nf3_4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM7 ds5_7 ds1_3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.500 W=w7_8 nf=nf7_8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 ds5_7 ds5_7 vss vss sky130_fd_pr__nfet_01v8 L=0.500 W=w5_6 nf=nf5_6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 out ds5_7 vss vss sky130_fd_pr__nfet_01v8 L=0.500 W=w5_6 nf=nf5_6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xM8 out ds2_4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.500 W=w7_8 nf=nf7_8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 source itail vss vss sky130_fd_pr__nfet_01v8 L=0.500 W=w9_10 nf=nf9_10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 itail itail vss vss sky130_fd_pr__nfet_01v8 L=0.500 W=w9_10 nf=nf1_2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.subckt cm_ota_extracted ID VOUT VINN VINP VSS VDD
X0 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X1 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X2 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X3 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X4 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X5 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X6 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X7 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X8 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X9 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X10 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X11 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X12 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X13 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X14 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X15 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X16 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X17 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X18 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X19 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X20 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X21 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X22 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X23 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X24 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X25 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X26 VSS m2_8142_2604# m2_8142_2604# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X27 m2_8142_2604# m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X28 VDD m1_5762_1400# m1_5762_1400# VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X29 VDD m1_5762_1400# m1_5762_1400# VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X30 m1_5762_1400# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X31 m1_5762_1400# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X32 VDD m1_5762_1400# m1_5762_1400# VDD sky130_fd_pr__pfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X33 m1_5762_1400# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X34 VDD m1_5762_1400# m1_5762_1400# VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X35 VDD m1_5762_1400# m1_5762_1400# VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X36 m1_5762_1400# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X37 m1_5762_1400# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X38 VDD li_4705_1411# li_4705_1411# VDD sky130_fd_pr__pfet_01v8 ad=14 pd=168 as=0.588 ps=7 w=0.42 l=0.50
X39 VDD li_4705_1411# li_4705_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X40 li_4705_1411# li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X41 li_4705_1411# li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X42 VDD li_4705_1411# li_4705_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X43 li_4705_1411# li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X44 VDD li_4705_1411# li_4705_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X45 VDD li_4705_1411# li_4705_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X46 li_4705_1411# li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X47 li_4705_1411# li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X48 li_5393_1327# ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X49 VSS ID li_5393_1327# VSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X50 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X51 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X52 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X53 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X54 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X55 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X56 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X57 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X58 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X59 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X60 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X61 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X62 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X63 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X64 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X65 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X66 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X67 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X68 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X69 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X70 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X71 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X72 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X73 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X74 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X75 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X76 VSS m2_8142_2604# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X77 VOUT m2_8142_2604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X78 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X79 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X80 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X81 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X82 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X83 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X84 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X85 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X86 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X87 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X88 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X89 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X90 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X91 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X92 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X93 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X94 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X95 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X96 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X97 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X98 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X99 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X100 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X101 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X102 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X103 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X104 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X105 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X106 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X107 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X108 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X109 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X110 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X111 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X112 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X113 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X114 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X115 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X116 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X117 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X118 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X119 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X120 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X121 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X122 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X123 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X124 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X125 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X126 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X127 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X128 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X129 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X130 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X131 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X132 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X133 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X134 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X135 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X136 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X137 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X138 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X139 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X140 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X141 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X142 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X143 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X144 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X145 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X146 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X147 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X148 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X149 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X150 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X151 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X152 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X153 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X154 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X155 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X156 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X157 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X158 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X159 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X160 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X161 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X162 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X163 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X164 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X165 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X166 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X167 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X168 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X169 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X170 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X171 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X172 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X173 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X174 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X175 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X176 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X177 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X178 VDD li_4705_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X179 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X180 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X181 VOUT li_4705_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.50
X182 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=6.12 ps=72.8 w=0.42 l=0.50
X183 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X184 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X185 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X186 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X187 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X188 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X189 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X190 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X191 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X192 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X193 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X194 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X195 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X196 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X197 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X198 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X199 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X200 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X201 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X202 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X203 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X204 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X205 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X206 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X207 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X208 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X209 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X210 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X211 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X212 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X213 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X214 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X215 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X216 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X217 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X218 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X219 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X220 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X221 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X222 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X223 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X224 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X225 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X226 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X227 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X228 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X229 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X230 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X231 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X232 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X233 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X234 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X235 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X236 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X237 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X238 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X239 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X240 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X241 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X242 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X243 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X244 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X245 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X246 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X247 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X248 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X249 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X250 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X251 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X252 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X253 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X254 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X255 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X256 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X257 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X258 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X259 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X260 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X261 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X262 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X263 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X264 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X265 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X266 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X267 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X268 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X269 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X270 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X271 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X272 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X273 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X274 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X275 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X276 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X277 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X278 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X279 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X280 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X281 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X282 VDD m1_5762_1400# m2_8142_2604# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X283 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X284 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X285 m2_8142_2604# m1_5762_1400# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X286 m1_5762_1400# VINP li_5393_1327# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X287 li_5393_1327# VINP m1_5762_1400# VSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
X288 li_4705_1411# VINN li_5393_1327# VSS sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.563 ps=6.88 w=0.42 l=0.50
X289 li_5393_1327# VINN li_4705_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.50
X290 ID ID VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.50
X291 VSS ID ID VSS sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.50
C0 VINP VDD 0.043f
C1 li_4705_1411# VINN 0.151f
C2 m1_5762_1400# ID 0.0259f
C3 li_4705_1411# m1_5762_1400# 0.0211f
C4 li_5393_1327# VDD 0.221f
C5 m2_8142_2604# VDD 42.5f
C6 VINP ID 0.0019f
C7 VOUT m2_8142_2604# 1.44f
C8 VINP VINN 0.041f
C9 li_5393_1327# ID 0.168f
C10 li_5393_1327# li_4705_1411# 0.711f
C11 VINP m1_5762_1400# 0.151f
C12 li_5393_1327# VINN 0.103f
C13 m2_8142_2604# ID 0.0122f
C14 li_4705_1411# m2_8142_2604# 0.813f
C15 li_5393_1327# m1_5762_1400# 0.734f
C16 m1_5762_1400# m2_8142_2604# 8.09f
C17 VOUT VDD 40.2f
C18 VINP li_5393_1327# 0.104f
C19 VDD ID 0.12f
C20 li_4705_1411# VDD 38.4f
C21 VINN VDD 0.042f
C22 m1_5762_1400# VDD 38.7f
C23 VOUT ID 0.00132f
C24 li_4705_1411# VOUT 7.89f
C25 li_5393_1327# m2_8142_2604# 1.02e-19
C26 m1_5762_1400# VOUT 3.68e-20
C27 li_4705_1411# ID 0.0578f
C28 VINN ID 0.0026f
C29 ID VSS 3.4f
C30 VINN VSS 0.805f
C31 VINP VSS 0.798f
C32 li_4705_1411# VSS 4.61f
C33 VOUT VSS 11.9f
C34 li_5393_1327# VSS 1.76f
C35 VDD VSS 98.6f
C36 m1_5762_1400# VSS 4.44f
C37 m2_8142_2604# VSS 31.1f
.ends

.GLOBAL GND
.end
