* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
*   mismatch {
*   }
* }
* 4-terminal Vertical Parallel Plate Capacitor /w LI-M4 fingers and M5 Shield
* 4-terminal Vertical Parallel Plate Capacitor /w LI-M4 fingers and Poly/M5 Shield
* Layout: sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x
.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x c0 c1 b m5
+ 
.param  mult = 1 presim_flag = 0.0
+ 
+ ctot_a = {141.23e-15*sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor+1.5*0.00244/sqrt(mult/0.21936)*141.23e-15*sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor*sky130_fd_pr__model__cap_vpp_only_p__slope}
+ cm5_c0 = {((2.074e-15)*c0m5m4_vpp0p4shield+(2.916e-15*presim_flag))}
+ cm5_c1 = {((3.67e-15)*c1m5m4_vpp0p4shield)}
+ cpl2s = {((15.22e-15)*cpl2s_vpp0p4shield+(2.84e-15*presim_flag))}
+ rat_m4 = 0.1120
+ rat_m3 = 0.1120
+ rat_m2 = 0.2836
+ rat_m1 = 0.2801
+ rat_li = 0.1863
+ rat_li2p = 0.026
+ cap_m4 = {rat_m4*ctot_a}
+ cap_m3 = {rat_m3*ctot_a}
+ cap_m2 = {rat_m2*ctot_a}
+ cap_m1 = {rat_m1*ctot_a}
+ cap_li = {rat_li*ctot_a}
+ cap_li2p = {rat_li2p*ctot_a}
+ ll1 = 5.070
+ lm1 = 5.215
+ lm2 = 5.095
+ lm3 = 5.050
+ lm4 = 4.910
+ wl1 = 0.170
+ wm1 = 0.140
+ wm2 = 0.140
+ wm3 = 0.300
+ wm4 = 0.300
+ nfl1 = 62.0
+ nfm1 = 72.0
+ nfm2 = 72.0
+ nfm3 = 34.0
+ nfm4 = 34.0
+ nvia3_c0 = 103.0
+ nvia3_c1 = 49.0
+ nvia2_c0 = 104.0
+ nvia2_c1 = 49.0
+ nvia_c0 = 124.0
+ nvia_c1 = 62.0
+ ncon_c0 = 116.0
+ ncon_c1 = 28.0
+ nlicon = 126.0
ccmvpp11p5x11p7_polym50p4shield m5 a0  c = {cm5_c0}
cm5_1 m5 a1 c = {cm5_c1}
rsm4 a0 a2 r = {rm4*lm4/wm4*(1/3)*(1/nfm4)}
cm4 a2 a1 c = {cap_m4}
rvia3_0 a0 b0 r = {rcvia3/nvia3_c0}
rvia3_1 a1 b1 r = {rcvia3/nvia3_c1}
rsm3 b0 b2 r = {rm3*lm3/wm3*(1/3)*(1/nfm3)}
cm3 b2 b1 c = {cap_m3}
rvia2_0 b0 c0 r = {rcvia2/nvia2_c0}
rvia2_1 b1 c1 r = {rcvia2/nvia2_c1}
rsm2 c0 c2 r = {rm2*lm2/wm2*(1/3)*(1/nfm2)}
cm2 c2 c1 c = {cap_m2}
rvia_0 c0 d0 r = {rcvia/nvia_c0}
rvia_1 c1 d1 r = {rcvia/nvia_c1}
rsm1 d0 d2 r = {rm1*lm1/wm1*(1/3)*(1/nfm1)}
cm1 d2 d1 c = {cap_m1}
rcon1 d0 e0 r = {rcl1/ncon_c0}
rcon2 d1 e1 r = {rcl1/ncon_c1}
rli1 e0 e2 r = {rl1*ll1/wl1*(1/3)*(1/nfl1)}
cli e2 e1 c = {cap_li}
rlicon e0 f0 r = {rcp1/nlicon}
rpoly f0 f2 r = {rp1}
cl12p e1 f2 c = {cap_li2p}
cpl2b f0 b c = {cpl2s}
.ends sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x
