VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO myconfig
   CLASS BLOCK ;
   SIZE 454.62 BY 328.82 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.28 0.0 82.66 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.4 0.0 88.78 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 0.0 94.22 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.28 0.0 99.66 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.4 0.0 105.78 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 0.0 111.22 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.96 0.0 117.34 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 0.0 122.78 1.06 ;
      END
   END din0[7]
   PIN din1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  320.96 327.76 321.34 328.82 ;
      END
   END din1[0]
   PIN din1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.08 327.76 327.46 328.82 ;
      END
   END din1[1]
   PIN din1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  333.2 327.76 333.58 328.82 ;
      END
   END din1[2]
   PIN din1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  338.64 327.76 339.02 328.82 ;
      END
   END din1[3]
   PIN din1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.76 327.76 345.14 328.82 ;
      END
   END din1[4]
   PIN din1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 327.76 351.26 328.82 ;
      END
   END din1[5]
   PIN din1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  356.32 327.76 356.7 328.82 ;
      END
   END din1[6]
   PIN din1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  362.44 327.76 362.82 328.82 ;
      END
   END din1[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  64.6 0.0 64.98 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.04 0.0 70.42 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.48 0.0 75.86 1.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 134.64 1.06 135.02 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 144.84 1.06 145.22 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 1.06 149.98 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.76 1.06 158.14 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 164.56 1.06 164.94 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 172.04 1.06 172.42 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  383.52 327.76 383.9 328.82 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 327.76 377.78 328.82 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 327.76 372.34 328.82 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 97.92 454.62 98.3 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 89.76 454.62 90.14 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 84.32 454.62 84.7 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 75.48 454.62 75.86 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 70.04 454.62 70.42 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 61.88 454.62 62.26 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 42.16 1.06 42.54 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 285.6 454.62 285.98 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 50.32 1.06 50.7 ;
      END
   END web0
   PIN web1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 277.44 454.62 277.82 ;
      END
   END web1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 44.2 1.06 44.58 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  453.56 284.92 454.62 285.3 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  126.48 0.0 126.86 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  152.32 0.0 152.7 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 0.0 177.18 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.12 0.0 227.5 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 252.66 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 0.0 277.14 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.92 0.0 302.3 1.06 ;
      END
   END dout0[7]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 327.76 127.54 328.82 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  152.32 327.76 152.7 328.82 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 327.76 177.18 328.82 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 327.76 202.34 328.82 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.12 327.76 227.5 328.82 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 327.76 252.66 328.82 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 327.76 277.14 328.82 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.92 327.76 302.3 328.82 ;
      END
   END dout1[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.4 323.68 451.22 325.42 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 325.42 ;
         LAYER met3 ;
         RECT  3.4 3.4 451.22 5.14 ;
         LAYER met4 ;
         RECT  449.48 3.4 451.22 325.42 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 327.08 454.62 328.82 ;
         LAYER met3 ;
         RECT  0.0 0.0 454.62 1.74 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 328.82 ;
         LAYER met4 ;
         RECT  452.88 0.0 454.62 328.82 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 454.0 328.2 ;
   LAYER  met2 ;
      RECT  0.62 0.62 454.0 328.2 ;
   LAYER  met3 ;
      RECT  1.66 134.04 454.0 135.62 ;
      RECT  0.62 135.62 1.66 144.24 ;
      RECT  0.62 145.82 1.66 149.0 ;
      RECT  0.62 150.58 1.66 157.16 ;
      RECT  0.62 158.74 1.66 163.96 ;
      RECT  0.62 165.54 1.66 171.44 ;
      RECT  1.66 97.32 452.96 98.9 ;
      RECT  1.66 98.9 452.96 134.04 ;
      RECT  452.96 98.9 454.0 134.04 ;
      RECT  452.96 90.74 454.0 97.32 ;
      RECT  452.96 85.3 454.0 89.16 ;
      RECT  452.96 76.46 454.0 83.72 ;
      RECT  452.96 71.02 454.0 74.88 ;
      RECT  452.96 62.86 454.0 69.44 ;
      RECT  1.66 135.62 452.96 285.0 ;
      RECT  1.66 285.0 452.96 286.58 ;
      RECT  0.62 51.3 1.66 134.04 ;
      RECT  452.96 135.62 454.0 276.84 ;
      RECT  0.62 43.14 1.66 43.6 ;
      RECT  0.62 45.18 1.66 49.72 ;
      RECT  452.96 278.42 454.0 284.32 ;
      RECT  1.66 286.58 2.8 323.08 ;
      RECT  1.66 323.08 2.8 326.02 ;
      RECT  2.8 286.58 451.82 323.08 ;
      RECT  451.82 286.58 452.96 323.08 ;
      RECT  451.82 323.08 452.96 326.02 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 97.32 ;
      RECT  2.8 5.74 451.82 97.32 ;
      RECT  451.82 2.8 452.96 5.74 ;
      RECT  451.82 5.74 452.96 97.32 ;
      RECT  0.62 173.02 1.66 326.48 ;
      RECT  452.96 286.58 454.0 326.48 ;
      RECT  1.66 326.02 2.8 326.48 ;
      RECT  2.8 326.02 451.82 326.48 ;
      RECT  451.82 326.02 452.96 326.48 ;
      RECT  452.96 2.34 454.0 61.28 ;
      RECT  0.62 2.34 1.66 41.56 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 451.82 2.8 ;
      RECT  451.82 2.34 452.96 2.8 ;
   LAYER  met4 ;
      RECT  81.68 1.66 83.26 328.2 ;
      RECT  83.26 0.62 87.8 1.66 ;
      RECT  89.38 0.62 93.24 1.66 ;
      RECT  94.82 0.62 98.68 1.66 ;
      RECT  100.26 0.62 104.8 1.66 ;
      RECT  106.38 0.62 110.24 1.66 ;
      RECT  111.82 0.62 116.36 1.66 ;
      RECT  117.94 0.62 121.8 1.66 ;
      RECT  83.26 1.66 320.36 327.16 ;
      RECT  320.36 1.66 321.94 327.16 ;
      RECT  321.94 327.16 326.48 328.2 ;
      RECT  328.06 327.16 332.6 328.2 ;
      RECT  334.18 327.16 338.04 328.2 ;
      RECT  339.62 327.16 344.16 328.2 ;
      RECT  345.74 327.16 350.28 328.2 ;
      RECT  351.86 327.16 355.72 328.2 ;
      RECT  357.3 327.16 361.84 328.2 ;
      RECT  65.58 0.62 69.44 1.66 ;
      RECT  71.02 0.62 74.88 1.66 ;
      RECT  76.46 0.62 81.68 1.66 ;
      RECT  378.38 327.16 382.92 328.2 ;
      RECT  363.42 327.16 371.36 328.2 ;
      RECT  372.94 327.16 376.8 328.2 ;
      RECT  123.38 0.62 125.88 1.66 ;
      RECT  127.46 0.62 151.72 1.66 ;
      RECT  153.3 0.62 176.2 1.66 ;
      RECT  177.78 0.62 201.36 1.66 ;
      RECT  202.94 0.62 226.52 1.66 ;
      RECT  228.1 0.62 251.68 1.66 ;
      RECT  253.26 0.62 276.16 1.66 ;
      RECT  277.74 0.62 301.32 1.66 ;
      RECT  83.26 327.16 126.56 328.2 ;
      RECT  128.14 327.16 151.72 328.2 ;
      RECT  153.3 327.16 176.2 328.2 ;
      RECT  177.78 327.16 201.36 328.2 ;
      RECT  202.94 327.16 226.52 328.2 ;
      RECT  228.1 327.16 251.68 328.2 ;
      RECT  253.26 327.16 276.16 328.2 ;
      RECT  277.74 327.16 301.32 328.2 ;
      RECT  302.9 327.16 320.36 328.2 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 326.02 5.74 328.2 ;
      RECT  5.74 1.66 81.68 2.8 ;
      RECT  5.74 2.8 81.68 326.02 ;
      RECT  5.74 326.02 81.68 328.2 ;
      RECT  321.94 1.66 448.88 2.8 ;
      RECT  321.94 2.8 448.88 326.02 ;
      RECT  321.94 326.02 448.88 327.16 ;
      RECT  448.88 1.66 451.82 2.8 ;
      RECT  448.88 326.02 451.82 327.16 ;
      RECT  2.34 0.62 64.0 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 326.02 ;
      RECT  2.34 326.02 2.8 328.2 ;
      RECT  384.5 327.16 452.28 328.2 ;
      RECT  302.9 0.62 452.28 1.66 ;
      RECT  451.82 1.66 452.28 2.8 ;
      RECT  451.82 2.8 452.28 326.02 ;
      RECT  451.82 326.02 452.28 327.16 ;
   END
END    myconfig
END    LIBRARY
