# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50 ;
  ORIGIN -0.070000  0.000000 ;
  SIZE  6.670000 BY  8.980000 ;
  PIN DRAIN
    ANTENNADIFFAREA  3.970400 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 2.890000 6.740000 6.090000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  14.179999 ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.000000 4.810000 0.685000 ;
        RECT 2.000000 8.295000 4.810000 8.980000 ;
      LAYER mcon ;
        RECT 2.060000 0.095000 4.750000 0.625000 ;
        RECT 2.060000 8.355000 4.750000 8.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.000000 0.000000 4.810000 0.685000 ;
        RECT 2.000000 8.295000 4.810000 8.980000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  5.955600 ;
    PORT
      LAYER met2 ;
        RECT 0.070000 1.010000 6.740000 2.610000 ;
        RECT 0.070000 6.370000 6.740000 7.970000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    ANTENNADIFFAREA  7.090000 ;
    ANTENNAGATEAREA  3.545000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 1.010000 0.500000 7.970000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.310000 1.010000 6.605000 7.970000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.205000 0.925000 1.150000 8.055000 ;
      RECT 0.950000 0.485000 1.280000 0.815000 ;
      RECT 0.950000 0.815000 1.150000 0.925000 ;
      RECT 0.950000 8.055000 1.150000 8.165000 ;
      RECT 0.950000 8.165000 1.280000 8.495000 ;
      RECT 1.760000 0.925000 1.930000 8.055000 ;
      RECT 2.540000 0.925000 2.710000 8.055000 ;
      RECT 3.320000 0.925000 3.490000 8.055000 ;
      RECT 4.100000 0.925000 4.270000 8.055000 ;
      RECT 4.880000 0.925000 5.050000 8.055000 ;
      RECT 5.530000 0.485000 5.860000 0.815000 ;
      RECT 5.530000 8.165000 5.860000 8.495000 ;
      RECT 5.660000 0.815000 5.860000 0.925000 ;
      RECT 5.660000 0.925000 6.605000 8.055000 ;
      RECT 5.660000 8.055000 5.860000 8.165000 ;
    LAYER mcon ;
      RECT 0.300000 1.165000 0.470000 1.335000 ;
      RECT 0.300000 1.525000 0.470000 1.695000 ;
      RECT 0.300000 1.885000 0.470000 2.055000 ;
      RECT 0.300000 2.245000 0.470000 2.415000 ;
      RECT 0.300000 2.605000 0.470000 2.775000 ;
      RECT 0.300000 2.965000 0.470000 3.135000 ;
      RECT 0.300000 3.325000 0.470000 3.495000 ;
      RECT 0.300000 3.685000 0.470000 3.855000 ;
      RECT 0.300000 4.045000 0.470000 4.215000 ;
      RECT 0.300000 4.405000 0.470000 4.575000 ;
      RECT 0.300000 4.765000 0.470000 4.935000 ;
      RECT 0.300000 5.125000 0.470000 5.295000 ;
      RECT 0.300000 5.485000 0.470000 5.655000 ;
      RECT 0.300000 5.845000 0.470000 6.015000 ;
      RECT 0.300000 6.205000 0.470000 6.375000 ;
      RECT 0.300000 6.565000 0.470000 6.735000 ;
      RECT 0.300000 6.925000 0.470000 7.095000 ;
      RECT 0.300000 7.285000 0.470000 7.455000 ;
      RECT 0.300000 7.645000 0.470000 7.815000 ;
      RECT 1.760000 1.165000 1.930000 1.335000 ;
      RECT 1.760000 1.525000 1.930000 1.695000 ;
      RECT 1.760000 1.885000 1.930000 2.055000 ;
      RECT 1.760000 2.245000 1.930000 2.415000 ;
      RECT 1.760000 2.605000 1.930000 2.775000 ;
      RECT 1.760000 2.965000 1.930000 3.135000 ;
      RECT 1.760000 3.325000 1.930000 3.495000 ;
      RECT 1.760000 3.685000 1.930000 3.855000 ;
      RECT 1.760000 4.045000 1.930000 4.215000 ;
      RECT 1.760000 4.405000 1.930000 4.575000 ;
      RECT 1.760000 4.765000 1.930000 4.935000 ;
      RECT 1.760000 5.125000 1.930000 5.295000 ;
      RECT 1.760000 5.485000 1.930000 5.655000 ;
      RECT 1.760000 5.845000 1.930000 6.015000 ;
      RECT 1.760000 6.205000 1.930000 6.375000 ;
      RECT 1.760000 6.565000 1.930000 6.735000 ;
      RECT 1.760000 6.925000 1.930000 7.095000 ;
      RECT 1.760000 7.285000 1.930000 7.455000 ;
      RECT 1.760000 7.645000 1.930000 7.815000 ;
      RECT 2.540000 1.165000 2.710000 1.335000 ;
      RECT 2.540000 1.525000 2.710000 1.695000 ;
      RECT 2.540000 1.885000 2.710000 2.055000 ;
      RECT 2.540000 2.245000 2.710000 2.415000 ;
      RECT 2.540000 2.605000 2.710000 2.775000 ;
      RECT 2.540000 2.965000 2.710000 3.135000 ;
      RECT 2.540000 3.325000 2.710000 3.495000 ;
      RECT 2.540000 3.685000 2.710000 3.855000 ;
      RECT 2.540000 4.045000 2.710000 4.215000 ;
      RECT 2.540000 4.405000 2.710000 4.575000 ;
      RECT 2.540000 4.765000 2.710000 4.935000 ;
      RECT 2.540000 5.125000 2.710000 5.295000 ;
      RECT 2.540000 5.485000 2.710000 5.655000 ;
      RECT 2.540000 5.845000 2.710000 6.015000 ;
      RECT 2.540000 6.205000 2.710000 6.375000 ;
      RECT 2.540000 6.565000 2.710000 6.735000 ;
      RECT 2.540000 6.925000 2.710000 7.095000 ;
      RECT 2.540000 7.285000 2.710000 7.455000 ;
      RECT 2.540000 7.645000 2.710000 7.815000 ;
      RECT 3.320000 1.165000 3.490000 1.335000 ;
      RECT 3.320000 1.525000 3.490000 1.695000 ;
      RECT 3.320000 1.885000 3.490000 2.055000 ;
      RECT 3.320000 2.245000 3.490000 2.415000 ;
      RECT 3.320000 2.605000 3.490000 2.775000 ;
      RECT 3.320000 2.965000 3.490000 3.135000 ;
      RECT 3.320000 3.325000 3.490000 3.495000 ;
      RECT 3.320000 3.685000 3.490000 3.855000 ;
      RECT 3.320000 4.045000 3.490000 4.215000 ;
      RECT 3.320000 4.405000 3.490000 4.575000 ;
      RECT 3.320000 4.765000 3.490000 4.935000 ;
      RECT 3.320000 5.125000 3.490000 5.295000 ;
      RECT 3.320000 5.485000 3.490000 5.655000 ;
      RECT 3.320000 5.845000 3.490000 6.015000 ;
      RECT 3.320000 6.205000 3.490000 6.375000 ;
      RECT 3.320000 6.565000 3.490000 6.735000 ;
      RECT 3.320000 6.925000 3.490000 7.095000 ;
      RECT 3.320000 7.285000 3.490000 7.455000 ;
      RECT 3.320000 7.645000 3.490000 7.815000 ;
      RECT 4.100000 1.165000 4.270000 1.335000 ;
      RECT 4.100000 1.525000 4.270000 1.695000 ;
      RECT 4.100000 1.885000 4.270000 2.055000 ;
      RECT 4.100000 2.245000 4.270000 2.415000 ;
      RECT 4.100000 2.605000 4.270000 2.775000 ;
      RECT 4.100000 2.965000 4.270000 3.135000 ;
      RECT 4.100000 3.325000 4.270000 3.495000 ;
      RECT 4.100000 3.685000 4.270000 3.855000 ;
      RECT 4.100000 4.045000 4.270000 4.215000 ;
      RECT 4.100000 4.405000 4.270000 4.575000 ;
      RECT 4.100000 4.765000 4.270000 4.935000 ;
      RECT 4.100000 5.125000 4.270000 5.295000 ;
      RECT 4.100000 5.485000 4.270000 5.655000 ;
      RECT 4.100000 5.845000 4.270000 6.015000 ;
      RECT 4.100000 6.205000 4.270000 6.375000 ;
      RECT 4.100000 6.565000 4.270000 6.735000 ;
      RECT 4.100000 6.925000 4.270000 7.095000 ;
      RECT 4.100000 7.285000 4.270000 7.455000 ;
      RECT 4.100000 7.645000 4.270000 7.815000 ;
      RECT 4.880000 1.165000 5.050000 1.335000 ;
      RECT 4.880000 1.525000 5.050000 1.695000 ;
      RECT 4.880000 1.885000 5.050000 2.055000 ;
      RECT 4.880000 2.245000 5.050000 2.415000 ;
      RECT 4.880000 2.605000 5.050000 2.775000 ;
      RECT 4.880000 2.965000 5.050000 3.135000 ;
      RECT 4.880000 3.325000 5.050000 3.495000 ;
      RECT 4.880000 3.685000 5.050000 3.855000 ;
      RECT 4.880000 4.045000 5.050000 4.215000 ;
      RECT 4.880000 4.405000 5.050000 4.575000 ;
      RECT 4.880000 4.765000 5.050000 4.935000 ;
      RECT 4.880000 5.125000 5.050000 5.295000 ;
      RECT 4.880000 5.485000 5.050000 5.655000 ;
      RECT 4.880000 5.845000 5.050000 6.015000 ;
      RECT 4.880000 6.205000 5.050000 6.375000 ;
      RECT 4.880000 6.565000 5.050000 6.735000 ;
      RECT 4.880000 6.925000 5.050000 7.095000 ;
      RECT 4.880000 7.285000 5.050000 7.455000 ;
      RECT 4.880000 7.645000 5.050000 7.815000 ;
      RECT 6.340000 1.165000 6.510000 1.335000 ;
      RECT 6.340000 1.525000 6.510000 1.695000 ;
      RECT 6.340000 1.885000 6.510000 2.055000 ;
      RECT 6.340000 2.245000 6.510000 2.415000 ;
      RECT 6.340000 2.605000 6.510000 2.775000 ;
      RECT 6.340000 2.965000 6.510000 3.135000 ;
      RECT 6.340000 3.325000 6.510000 3.495000 ;
      RECT 6.340000 3.685000 6.510000 3.855000 ;
      RECT 6.340000 4.045000 6.510000 4.215000 ;
      RECT 6.340000 4.405000 6.510000 4.575000 ;
      RECT 6.340000 4.765000 6.510000 4.935000 ;
      RECT 6.340000 5.125000 6.510000 5.295000 ;
      RECT 6.340000 5.485000 6.510000 5.655000 ;
      RECT 6.340000 5.845000 6.510000 6.015000 ;
      RECT 6.340000 6.205000 6.510000 6.375000 ;
      RECT 6.340000 6.565000 6.510000 6.735000 ;
      RECT 6.340000 6.925000 6.510000 7.095000 ;
      RECT 6.340000 7.285000 6.510000 7.455000 ;
      RECT 6.340000 7.645000 6.510000 7.815000 ;
    LAYER met1 ;
      RECT 1.715000 1.010000 1.975000 7.970000 ;
      RECT 2.495000 1.010000 2.755000 7.970000 ;
      RECT 3.275000 1.010000 3.535000 7.970000 ;
      RECT 4.055000 1.010000 4.315000 7.970000 ;
      RECT 4.835000 1.010000 5.095000 7.970000 ;
    LAYER via ;
      RECT 1.715000 1.040000 1.975000 1.300000 ;
      RECT 1.715000 1.360000 1.975000 1.620000 ;
      RECT 1.715000 1.680000 1.975000 1.940000 ;
      RECT 1.715000 2.000000 1.975000 2.260000 ;
      RECT 1.715000 2.320000 1.975000 2.580000 ;
      RECT 1.715000 6.400000 1.975000 6.660000 ;
      RECT 1.715000 6.720000 1.975000 6.980000 ;
      RECT 1.715000 7.040000 1.975000 7.300000 ;
      RECT 1.715000 7.360000 1.975000 7.620000 ;
      RECT 1.715000 7.680000 1.975000 7.940000 ;
      RECT 2.495000 2.920000 2.755000 3.180000 ;
      RECT 2.495000 3.240000 2.755000 3.500000 ;
      RECT 2.495000 3.560000 2.755000 3.820000 ;
      RECT 2.495000 3.880000 2.755000 4.140000 ;
      RECT 2.495000 4.200000 2.755000 4.460000 ;
      RECT 2.495000 4.520000 2.755000 4.780000 ;
      RECT 2.495000 4.840000 2.755000 5.100000 ;
      RECT 2.495000 5.160000 2.755000 5.420000 ;
      RECT 2.495000 5.480000 2.755000 5.740000 ;
      RECT 2.495000 5.800000 2.755000 6.060000 ;
      RECT 3.275000 1.040000 3.535000 1.300000 ;
      RECT 3.275000 1.360000 3.535000 1.620000 ;
      RECT 3.275000 1.680000 3.535000 1.940000 ;
      RECT 3.275000 2.000000 3.535000 2.260000 ;
      RECT 3.275000 2.320000 3.535000 2.580000 ;
      RECT 3.275000 6.400000 3.535000 6.660000 ;
      RECT 3.275000 6.720000 3.535000 6.980000 ;
      RECT 3.275000 7.040000 3.535000 7.300000 ;
      RECT 3.275000 7.360000 3.535000 7.620000 ;
      RECT 3.275000 7.680000 3.535000 7.940000 ;
      RECT 4.055000 2.920000 4.315000 3.180000 ;
      RECT 4.055000 3.240000 4.315000 3.500000 ;
      RECT 4.055000 3.560000 4.315000 3.820000 ;
      RECT 4.055000 3.880000 4.315000 4.140000 ;
      RECT 4.055000 4.200000 4.315000 4.460000 ;
      RECT 4.055000 4.520000 4.315000 4.780000 ;
      RECT 4.055000 4.840000 4.315000 5.100000 ;
      RECT 4.055000 5.160000 4.315000 5.420000 ;
      RECT 4.055000 5.480000 4.315000 5.740000 ;
      RECT 4.055000 5.800000 4.315000 6.060000 ;
      RECT 4.835000 1.040000 5.095000 1.300000 ;
      RECT 4.835000 1.360000 5.095000 1.620000 ;
      RECT 4.835000 1.680000 5.095000 1.940000 ;
      RECT 4.835000 2.000000 5.095000 2.260000 ;
      RECT 4.835000 2.320000 5.095000 2.580000 ;
      RECT 4.835000 6.400000 5.095000 6.660000 ;
      RECT 4.835000 6.720000 5.095000 6.980000 ;
      RECT 4.835000 7.040000 5.095000 7.300000 ;
      RECT 4.835000 7.360000 5.095000 7.620000 ;
      RECT 4.835000 7.680000 5.095000 7.940000 ;
  END
END sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50
END LIBRARY
