# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.34000 BY  11.69000 ;
  PIN C0
    ANTENNAGATEAREA  80.00000 ;
    PORT
      LAYER met4 ;
        RECT  0.300000 0.075000  0.630000 11.615000 ;
        RECT  1.595000 0.800000  1.895000  5.600000 ;
        RECT  1.595000 5.600000  9.745000  5.930000 ;
        RECT  1.595000 5.930000  1.895000 10.730000 ;
        RECT  2.795000 0.800000  3.095000  5.600000 ;
        RECT  2.795000 5.930000  3.095000 10.730000 ;
        RECT  3.995000 0.800000  4.295000  5.600000 ;
        RECT  3.995000 5.930000  4.295000 10.730000 ;
        RECT  5.310000 0.800000  5.835000  5.600000 ;
        RECT  5.310000 5.930000  5.835000 10.730000 ;
        RECT  7.045000 0.800000  7.345000  5.600000 ;
        RECT  7.045000 5.930000  7.345000 10.730000 ;
        RECT  8.245000 0.800000  8.545000  5.600000 ;
        RECT  8.245000 5.930000  8.545000 10.730000 ;
        RECT  9.445000 0.800000  9.745000  5.600000 ;
        RECT  9.445000 5.930000  9.745000 10.730000 ;
        RECT 10.710000 0.075000 11.040000 11.615000 ;
    END
  END C0
  PIN C1
    ANTENNADIFFAREA  29.799999 ;
    PORT
      LAYER met4 ;
        RECT  0.965000  0.170000 10.375000  0.500000 ;
        RECT  0.965000  0.500000  1.295000 11.030000 ;
        RECT  0.965000 11.030000 10.375000 11.330000 ;
        RECT  0.965000 11.330000 10.045000 11.360000 ;
        RECT  2.195000  0.500000  2.495000  5.300000 ;
        RECT  2.195000  6.230000  2.495000 11.030000 ;
        RECT  3.395000  0.500000  3.695000  5.300000 ;
        RECT  3.395000  6.230000  3.695000 11.030000 ;
        RECT  4.595000  0.500000  5.010000  5.300000 ;
        RECT  4.595000  6.230000  5.010000 11.030000 ;
        RECT  6.135000  0.500000  6.745000  5.300000 ;
        RECT  6.135000  6.230000  6.745000 11.030000 ;
        RECT  7.645000  0.500000  7.945000  5.300000 ;
        RECT  7.645000  6.230000  7.945000 11.030000 ;
        RECT  8.845000  0.500000  9.145000  5.300000 ;
        RECT  8.845000  6.230000  9.145000 11.030000 ;
        RECT 10.045000  0.500000 10.375000 11.030000 ;
    END
  END C1
  PIN MET5
    PORT
      LAYER met5 ;
        RECT 0.000000 0.000000 11.340000 11.690000 ;
    END
  END MET5
  OBS
    LAYER li1 ;
      RECT  0.465000  0.825000 10.875000  1.625000 ;
      RECT  0.465000  1.625000  1.175000  9.935000 ;
      RECT  0.465000  9.935000 10.875000 10.735000 ;
      RECT  1.355000  0.290000  9.980000  0.335000 ;
      RECT  1.355000  0.335000  9.985000  0.505000 ;
      RECT  1.355000  0.505000  9.980000  0.550000 ;
      RECT  1.355000 11.140000  9.980000 11.185000 ;
      RECT  1.355000 11.185000  9.985000 11.355000 ;
      RECT  1.355000 11.355000  9.980000 11.400000 ;
      RECT  1.450000  1.795000  1.620000  5.465000 ;
      RECT  1.450000  5.465000  5.260000  6.095000 ;
      RECT  1.450000  6.095000  1.620000  9.765000 ;
      RECT  1.800000  1.625000  1.970000  5.295000 ;
      RECT  1.800000  6.265000  1.970000  9.935000 ;
      RECT  2.150000  1.795000  2.320000  5.465000 ;
      RECT  2.150000  6.095000  2.320000  9.765000 ;
      RECT  2.500000  1.625000  2.670000  5.295000 ;
      RECT  2.500000  6.265000  2.670000  9.935000 ;
      RECT  2.850000  1.795000  3.020000  5.465000 ;
      RECT  2.850000  6.095000  3.020000  9.765000 ;
      RECT  3.200000  1.625000  3.370000  5.295000 ;
      RECT  3.200000  6.265000  3.370000  9.935000 ;
      RECT  3.550000  1.795000  3.720000  5.465000 ;
      RECT  3.550000  6.095000  3.720000  9.765000 ;
      RECT  3.900000  1.625000  4.070000  5.295000 ;
      RECT  3.900000  6.265000  4.070000  9.935000 ;
      RECT  4.250000  1.795000  4.420000  5.465000 ;
      RECT  4.250000  6.095000  4.420000  9.765000 ;
      RECT  4.600000  1.625000  4.770000  5.295000 ;
      RECT  4.600000  6.265000  4.770000  9.935000 ;
      RECT  4.950000  1.795000  5.120000  5.465000 ;
      RECT  4.950000  6.095000  5.120000  9.765000 ;
      RECT  5.300000  1.625000  6.040000  5.285000 ;
      RECT  5.300000  6.275000  5.900000  6.280000 ;
      RECT  5.300000  6.280000  6.040000  9.935000 ;
      RECT  5.440000  5.285000  5.900000  6.275000 ;
      RECT  6.080000  5.465000  9.890000  6.095000 ;
      RECT  6.220000  1.795000  6.390000  5.465000 ;
      RECT  6.220000  6.095000  6.390000  9.765000 ;
      RECT  6.570000  1.625000  6.740000  5.295000 ;
      RECT  6.570000  6.265000  6.740000  9.935000 ;
      RECT  6.920000  1.795000  7.090000  5.465000 ;
      RECT  6.920000  6.095000  7.090000  9.765000 ;
      RECT  7.270000  1.625000  7.440000  5.295000 ;
      RECT  7.270000  6.265000  7.440000  9.935000 ;
      RECT  7.620000  1.795000  7.790000  5.465000 ;
      RECT  7.620000  6.095000  7.790000  9.765000 ;
      RECT  7.970000  1.625000  8.140000  5.295000 ;
      RECT  7.970000  6.265000  8.140000  9.935000 ;
      RECT  8.320000  1.795000  8.490000  5.465000 ;
      RECT  8.320000  6.095000  8.490000  9.765000 ;
      RECT  8.670000  1.625000  8.840000  5.295000 ;
      RECT  8.670000  6.265000  8.840000  9.935000 ;
      RECT  9.020000  1.795000  9.190000  5.465000 ;
      RECT  9.020000  6.095000  9.190000  9.765000 ;
      RECT  9.370000  1.625000  9.540000  5.295000 ;
      RECT  9.370000  6.265000  9.540000  9.935000 ;
      RECT  9.720000  1.795000  9.890000  5.465000 ;
      RECT  9.720000  6.095000  9.890000  9.765000 ;
      RECT 10.165000  1.625000 10.875000  9.935000 ;
    LAYER mcon ;
      RECT  0.645000  1.015000  1.175000 10.545000 ;
      RECT  1.415000  0.335000  1.585000  0.505000 ;
      RECT  1.415000 11.185000  1.585000 11.355000 ;
      RECT  1.595000  1.405000  1.765000  1.575000 ;
      RECT  1.595000  9.985000  1.765000 10.155000 ;
      RECT  1.720000  5.515000  5.130000  6.045000 ;
      RECT  1.775000  0.335000  1.945000  0.505000 ;
      RECT  1.775000 11.185000  1.945000 11.355000 ;
      RECT  1.955000  1.405000  2.125000  1.575000 ;
      RECT  1.955000  9.985000  2.125000 10.155000 ;
      RECT  2.135000  0.335000  2.305000  0.505000 ;
      RECT  2.135000 11.185000  2.305000 11.355000 ;
      RECT  2.315000  1.405000  2.485000  1.575000 ;
      RECT  2.315000  9.985000  2.485000 10.155000 ;
      RECT  2.495000  0.335000  2.665000  0.505000 ;
      RECT  2.495000 11.185000  2.665000 11.355000 ;
      RECT  2.675000  1.405000  2.845000  1.575000 ;
      RECT  2.675000  9.985000  2.845000 10.155000 ;
      RECT  2.855000  0.335000  3.025000  0.505000 ;
      RECT  2.855000 11.185000  3.025000 11.355000 ;
      RECT  3.035000  1.405000  3.205000  1.575000 ;
      RECT  3.035000  9.985000  3.205000 10.155000 ;
      RECT  3.215000  0.335000  3.385000  0.505000 ;
      RECT  3.215000 11.185000  3.385000 11.355000 ;
      RECT  3.395000  1.405000  3.565000  1.575000 ;
      RECT  3.395000  9.985000  3.565000 10.155000 ;
      RECT  3.575000  0.335000  3.745000  0.505000 ;
      RECT  3.575000 11.185000  3.745000 11.355000 ;
      RECT  3.755000  1.405000  3.925000  1.575000 ;
      RECT  3.755000  9.985000  3.925000 10.155000 ;
      RECT  3.935000  0.335000  4.105000  0.505000 ;
      RECT  3.935000 11.185000  4.105000 11.355000 ;
      RECT  4.115000  1.405000  4.285000  1.575000 ;
      RECT  4.115000  9.985000  4.285000 10.155000 ;
      RECT  4.295000  0.335000  4.465000  0.505000 ;
      RECT  4.295000 11.185000  4.465000 11.355000 ;
      RECT  4.475000  1.405000  4.645000  1.575000 ;
      RECT  4.475000  9.985000  4.645000 10.155000 ;
      RECT  4.655000  0.335000  4.825000  0.505000 ;
      RECT  4.655000 11.185000  4.825000 11.355000 ;
      RECT  4.835000  1.405000  5.005000  1.575000 ;
      RECT  4.835000  9.985000  5.005000 10.155000 ;
      RECT  5.015000  0.335000  5.185000  0.505000 ;
      RECT  5.015000 11.185000  5.185000 11.355000 ;
      RECT  5.375000  0.335000  5.545000  0.505000 ;
      RECT  5.375000 11.185000  5.545000 11.355000 ;
      RECT  5.735000  0.335000  5.905000  0.505000 ;
      RECT  5.735000 11.185000  5.905000 11.355000 ;
      RECT  6.095000  0.335000  6.265000  0.505000 ;
      RECT  6.095000 11.185000  6.265000 11.355000 ;
      RECT  6.210000  5.515000  9.620000  6.045000 ;
      RECT  6.335000  1.405000  6.505000  1.575000 ;
      RECT  6.335000  9.985000  6.505000 10.155000 ;
      RECT  6.455000  0.335000  6.625000  0.505000 ;
      RECT  6.455000 11.185000  6.625000 11.355000 ;
      RECT  6.695000  1.405000  6.865000  1.575000 ;
      RECT  6.695000  9.985000  6.865000 10.155000 ;
      RECT  6.815000  0.335000  6.985000  0.505000 ;
      RECT  6.815000 11.185000  6.985000 11.355000 ;
      RECT  7.055000  1.405000  7.225000  1.575000 ;
      RECT  7.055000  9.985000  7.225000 10.155000 ;
      RECT  7.175000  0.335000  7.345000  0.505000 ;
      RECT  7.175000 11.185000  7.345000 11.355000 ;
      RECT  7.415000  1.405000  7.585000  1.575000 ;
      RECT  7.415000  9.985000  7.585000 10.155000 ;
      RECT  7.535000  0.335000  7.705000  0.505000 ;
      RECT  7.535000 11.185000  7.705000 11.355000 ;
      RECT  7.775000  1.405000  7.945000  1.575000 ;
      RECT  7.775000  9.985000  7.945000 10.155000 ;
      RECT  7.895000  0.335000  8.065000  0.505000 ;
      RECT  7.895000 11.185000  8.065000 11.355000 ;
      RECT  8.135000  1.405000  8.305000  1.575000 ;
      RECT  8.135000  9.985000  8.305000 10.155000 ;
      RECT  8.255000  0.335000  8.425000  0.505000 ;
      RECT  8.255000 11.185000  8.425000 11.355000 ;
      RECT  8.495000  1.405000  8.665000  1.575000 ;
      RECT  8.495000  9.985000  8.665000 10.155000 ;
      RECT  8.615000  0.335000  8.785000  0.505000 ;
      RECT  8.615000 11.185000  8.785000 11.355000 ;
      RECT  8.855000  1.405000  9.025000  1.575000 ;
      RECT  8.855000  9.985000  9.025000 10.155000 ;
      RECT  8.975000  0.335000  9.145000  0.505000 ;
      RECT  8.975000 11.185000  9.145000 11.355000 ;
      RECT  9.215000  1.405000  9.385000  1.575000 ;
      RECT  9.215000  9.985000  9.385000 10.155000 ;
      RECT  9.335000  0.335000  9.505000  0.505000 ;
      RECT  9.335000 11.185000  9.505000 11.355000 ;
      RECT  9.575000  1.405000  9.745000  1.575000 ;
      RECT  9.575000  9.985000  9.745000 10.155000 ;
      RECT  9.695000  0.335000  9.865000  0.505000 ;
      RECT  9.695000 11.185000  9.865000 11.355000 ;
      RECT 10.165000  1.015000 10.695000 10.545000 ;
    LAYER met1 ;
      RECT  0.465000  0.000000 10.875000  0.150000 ;
      RECT  0.465000  0.150000  1.215000  1.355000 ;
      RECT  0.465000  1.355000  5.120000  1.625000 ;
      RECT  0.465000  1.625000  1.310000  2.075000 ;
      RECT  0.465000  2.075000  5.120000  2.215000 ;
      RECT  0.465000  2.215000  1.310000  2.635000 ;
      RECT  0.465000  2.635000  5.120000  2.775000 ;
      RECT  0.465000  2.775000  1.310000  3.195000 ;
      RECT  0.465000  3.195000  5.120000  3.335000 ;
      RECT  0.465000  3.335000  1.310000  3.755000 ;
      RECT  0.465000  3.755000  5.120000  3.895000 ;
      RECT  0.465000  3.895000  1.310000  4.315000 ;
      RECT  0.465000  4.315000  5.120000  4.455000 ;
      RECT  0.465000  4.455000  1.310000  4.875000 ;
      RECT  0.465000  4.875000  5.120000  5.015000 ;
      RECT  0.465000  5.015000  1.310000  6.545000 ;
      RECT  0.465000  6.545000  5.120000  6.685000 ;
      RECT  0.465000  6.685000  1.310000  7.105000 ;
      RECT  0.465000  7.105000  5.120000  7.245000 ;
      RECT  0.465000  7.245000  1.310000  7.665000 ;
      RECT  0.465000  7.665000  5.120000  7.805000 ;
      RECT  0.465000  7.805000  1.310000  8.225000 ;
      RECT  0.465000  8.225000  5.120000  8.365000 ;
      RECT  0.465000  8.365000  1.310000  8.785000 ;
      RECT  0.465000  8.785000  5.120000  8.925000 ;
      RECT  0.465000  8.925000  1.310000  9.345000 ;
      RECT  0.465000  9.345000  5.120000  9.485000 ;
      RECT  0.465000  9.485000  1.310000  9.935000 ;
      RECT  0.465000  9.935000  5.120000 10.205000 ;
      RECT  0.465000 10.205000  1.215000 11.540000 ;
      RECT  0.465000 11.540000 10.875000 11.690000 ;
      RECT  1.355000  0.290000  9.980000  1.205000 ;
      RECT  1.355000 10.355000  9.980000 11.400000 ;
      RECT  1.450000  1.795000  9.890000  1.935000 ;
      RECT  1.450000  2.355000  9.890000  2.495000 ;
      RECT  1.450000  2.915000  9.890000  3.055000 ;
      RECT  1.450000  3.475000  9.890000  3.615000 ;
      RECT  1.450000  4.035000  9.890000  4.175000 ;
      RECT  1.450000  4.595000  9.890000  4.735000 ;
      RECT  1.450000  5.155000  9.890000  5.295000 ;
      RECT  1.450000  5.465000  9.890000  6.095000 ;
      RECT  1.450000  6.265000  9.890000  6.405000 ;
      RECT  1.450000  6.825000  9.890000  6.965000 ;
      RECT  1.450000  7.385000  9.890000  7.525000 ;
      RECT  1.450000  7.945000  9.890000  8.085000 ;
      RECT  1.450000  8.505000  9.890000  8.645000 ;
      RECT  1.450000  9.065000  9.890000  9.205000 ;
      RECT  1.450000  9.625000  9.890000  9.765000 ;
      RECT  5.260000  1.205000  6.080000  1.795000 ;
      RECT  5.260000  1.935000  6.080000  2.355000 ;
      RECT  5.260000  2.495000  6.080000  2.915000 ;
      RECT  5.260000  3.055000  6.080000  3.475000 ;
      RECT  5.260000  3.615000  6.080000  4.035000 ;
      RECT  5.260000  4.175000  6.080000  4.595000 ;
      RECT  5.260000  4.735000  6.080000  5.155000 ;
      RECT  5.260000  5.295000  6.080000  5.465000 ;
      RECT  5.260000  6.095000  6.080000  6.265000 ;
      RECT  5.260000  6.405000  6.080000  6.825000 ;
      RECT  5.260000  6.965000  6.080000  7.385000 ;
      RECT  5.260000  7.525000  6.080000  7.945000 ;
      RECT  5.260000  8.085000  6.080000  8.505000 ;
      RECT  5.260000  8.645000  6.080000  9.065000 ;
      RECT  5.260000  9.205000  6.080000  9.625000 ;
      RECT  5.260000  9.765000  6.080000 10.355000 ;
      RECT  6.220000  1.355000 10.875000  1.625000 ;
      RECT  6.220000  2.075000 10.875000  2.215000 ;
      RECT  6.220000  2.635000 10.875000  2.775000 ;
      RECT  6.220000  3.195000 10.875000  3.335000 ;
      RECT  6.220000  3.755000 10.875000  3.895000 ;
      RECT  6.220000  4.315000 10.875000  4.455000 ;
      RECT  6.220000  4.875000 10.875000  5.015000 ;
      RECT  6.220000  6.545000 10.875000  6.685000 ;
      RECT  6.220000  7.105000 10.875000  7.245000 ;
      RECT  6.220000  7.665000 10.875000  7.805000 ;
      RECT  6.220000  8.225000 10.875000  8.365000 ;
      RECT  6.220000  8.785000 10.875000  8.925000 ;
      RECT  6.220000  9.345000 10.875000  9.485000 ;
      RECT  6.220000  9.935000 10.875000 10.205000 ;
      RECT 10.030000  1.625000 10.875000  2.075000 ;
      RECT 10.030000  2.215000 10.875000  2.635000 ;
      RECT 10.030000  2.775000 10.875000  3.195000 ;
      RECT 10.030000  3.335000 10.875000  3.755000 ;
      RECT 10.030000  3.895000 10.875000  4.315000 ;
      RECT 10.030000  4.455000 10.875000  4.875000 ;
      RECT 10.030000  5.015000 10.875000  6.545000 ;
      RECT 10.030000  6.685000 10.875000  7.105000 ;
      RECT 10.030000  7.245000 10.875000  7.665000 ;
      RECT 10.030000  7.805000 10.875000  8.225000 ;
      RECT 10.030000  8.365000 10.875000  8.785000 ;
      RECT 10.030000  8.925000 10.875000  9.345000 ;
      RECT 10.030000  9.485000 10.875000  9.935000 ;
      RECT 10.120000  0.150000 10.875000  1.355000 ;
      RECT 10.120000 10.205000 10.875000 11.540000 ;
    LAYER met2 ;
      RECT  0.325000  0.075000 11.015000  1.205000 ;
      RECT  0.325000  1.205000  0.845000 10.355000 ;
      RECT  0.325000 10.355000 11.015000 11.615000 ;
      RECT  0.990000  1.355000  5.120000  1.625000 ;
      RECT  0.990000  1.625000  1.310000  1.795000 ;
      RECT  0.990000  1.795000  5.120000  1.935000 ;
      RECT  0.990000  1.935000  1.310000  2.355000 ;
      RECT  0.990000  2.355000  5.120000  2.495000 ;
      RECT  0.990000  2.495000  1.310000  2.915000 ;
      RECT  0.990000  2.915000  5.120000  3.055000 ;
      RECT  0.990000  3.055000  1.310000  3.475000 ;
      RECT  0.990000  3.475000  5.120000  3.615000 ;
      RECT  0.990000  3.615000  1.310000  4.035000 ;
      RECT  0.990000  4.035000  5.120000  4.175000 ;
      RECT  0.990000  4.175000  1.310000  4.595000 ;
      RECT  0.990000  4.595000  5.120000  4.735000 ;
      RECT  0.990000  4.735000  1.310000  5.155000 ;
      RECT  0.990000  5.155000  5.120000  5.295000 ;
      RECT  0.990000  5.295000  1.310000  6.265000 ;
      RECT  0.990000  6.265000  5.120000  6.405000 ;
      RECT  0.990000  6.405000  1.310000  6.825000 ;
      RECT  0.990000  6.825000  5.120000  6.965000 ;
      RECT  0.990000  6.965000  1.310000  7.385000 ;
      RECT  0.990000  7.385000  5.120000  7.525000 ;
      RECT  0.990000  7.525000  1.310000  7.945000 ;
      RECT  0.990000  7.945000  5.120000  8.085000 ;
      RECT  0.990000  8.085000  1.310000  8.505000 ;
      RECT  0.990000  8.505000  5.120000  8.645000 ;
      RECT  0.990000  8.645000  1.310000  9.065000 ;
      RECT  0.990000  9.065000  5.120000  9.205000 ;
      RECT  0.990000  9.205000  1.310000  9.625000 ;
      RECT  0.990000  9.625000  5.120000  9.765000 ;
      RECT  0.990000  9.765000  1.310000  9.935000 ;
      RECT  0.990000  9.935000  5.120000 10.205000 ;
      RECT  1.450000  2.075000  9.890000  2.215000 ;
      RECT  1.450000  2.635000  9.890000  2.775000 ;
      RECT  1.450000  3.195000  9.890000  3.335000 ;
      RECT  1.450000  3.755000  9.890000  3.895000 ;
      RECT  1.450000  4.315000  9.890000  4.455000 ;
      RECT  1.450000  4.875000  9.890000  5.015000 ;
      RECT  1.450000  5.465000  9.890000  6.095000 ;
      RECT  1.450000  6.545000  9.890000  6.685000 ;
      RECT  1.450000  7.105000  9.890000  7.245000 ;
      RECT  1.450000  7.665000  9.890000  7.805000 ;
      RECT  1.450000  8.225000  9.890000  8.365000 ;
      RECT  1.450000  8.785000  9.890000  8.925000 ;
      RECT  1.450000  9.345000  9.890000  9.485000 ;
      RECT  5.260000  1.205000  6.080000  2.075000 ;
      RECT  5.260000  2.215000  6.080000  2.635000 ;
      RECT  5.260000  2.775000  6.080000  3.195000 ;
      RECT  5.260000  3.335000  6.080000  3.755000 ;
      RECT  5.260000  3.895000  6.080000  4.315000 ;
      RECT  5.260000  4.455000  6.080000  4.875000 ;
      RECT  5.260000  5.015000  6.080000  5.465000 ;
      RECT  5.260000  6.095000  6.080000  6.545000 ;
      RECT  5.260000  6.685000  6.080000  7.105000 ;
      RECT  5.260000  7.245000  6.080000  7.665000 ;
      RECT  5.260000  7.805000  6.080000  8.225000 ;
      RECT  5.260000  8.365000  6.080000  8.785000 ;
      RECT  5.260000  8.925000  6.080000  9.345000 ;
      RECT  5.260000  9.485000  6.080000 10.355000 ;
      RECT  6.220000  1.355000 10.350000  1.625000 ;
      RECT  6.220000  1.795000 10.350000  1.935000 ;
      RECT  6.220000  2.355000 10.350000  2.495000 ;
      RECT  6.220000  2.915000 10.350000  3.055000 ;
      RECT  6.220000  3.475000 10.350000  3.615000 ;
      RECT  6.220000  4.035000 10.350000  4.175000 ;
      RECT  6.220000  4.595000 10.350000  4.735000 ;
      RECT  6.220000  5.155000 10.350000  5.295000 ;
      RECT  6.220000  6.265000 10.350000  6.405000 ;
      RECT  6.220000  6.825000 10.350000  6.965000 ;
      RECT  6.220000  7.385000 10.350000  7.525000 ;
      RECT  6.220000  7.945000 10.350000  8.085000 ;
      RECT  6.220000  8.505000 10.350000  8.645000 ;
      RECT  6.220000  9.065000 10.350000  9.205000 ;
      RECT  6.220000  9.625000 10.350000  9.765000 ;
      RECT  6.220000  9.935000 10.350000 10.205000 ;
      RECT 10.030000  1.625000 10.350000  1.795000 ;
      RECT 10.030000  1.935000 10.350000  2.355000 ;
      RECT 10.030000  2.495000 10.350000  2.915000 ;
      RECT 10.030000  3.055000 10.350000  3.475000 ;
      RECT 10.030000  3.615000 10.350000  4.035000 ;
      RECT 10.030000  4.175000 10.350000  4.595000 ;
      RECT 10.030000  4.735000 10.350000  5.155000 ;
      RECT 10.030000  5.295000 10.350000  6.265000 ;
      RECT 10.030000  6.405000 10.350000  6.825000 ;
      RECT 10.030000  6.965000 10.350000  7.385000 ;
      RECT 10.030000  7.525000 10.350000  7.945000 ;
      RECT 10.030000  8.085000 10.350000  8.505000 ;
      RECT 10.030000  8.645000 10.350000  9.065000 ;
      RECT 10.030000  9.205000 10.350000  9.625000 ;
      RECT 10.030000  9.765000 10.350000  9.935000 ;
      RECT 10.490000  1.205000 11.015000 10.355000 ;
    LAYER met3 ;
      RECT  0.300000  0.075000  0.630000 11.615000 ;
      RECT  0.965000  0.170000 10.375000  0.500000 ;
      RECT  0.965000  0.500000  1.295000  1.400000 ;
      RECT  0.965000  1.400000  5.205000  1.700000 ;
      RECT  0.965000  1.700000  1.295000  2.600000 ;
      RECT  0.965000  2.600000  5.205000  2.900000 ;
      RECT  0.965000  2.900000  1.295000  3.800000 ;
      RECT  0.965000  3.800000  5.205000  4.100000 ;
      RECT  0.965000  4.100000  1.295000  5.000000 ;
      RECT  0.965000  5.000000  5.205000  5.300000 ;
      RECT  0.965000  5.300000  1.295000  6.230000 ;
      RECT  0.965000  6.230000  5.205000  6.530000 ;
      RECT  0.965000  6.530000  1.295000  7.430000 ;
      RECT  0.965000  7.430000  5.205000  7.730000 ;
      RECT  0.965000  7.730000  1.295000  8.630000 ;
      RECT  0.965000  8.630000  5.205000  8.930000 ;
      RECT  0.965000  8.930000  1.295000  9.830000 ;
      RECT  0.965000  9.830000  5.205000 10.130000 ;
      RECT  0.965000 10.130000  1.295000 11.030000 ;
      RECT  0.965000 11.030000 10.375000 11.360000 ;
      RECT  1.595000  0.800000  9.745000  1.100000 ;
      RECT  1.595000  2.000000  9.745000  2.300000 ;
      RECT  1.595000  3.200000  9.745000  3.500000 ;
      RECT  1.595000  4.400000  9.745000  4.700000 ;
      RECT  1.595000  5.600000  9.745000  5.930000 ;
      RECT  1.595000  6.830000  9.745000  7.130000 ;
      RECT  1.595000  8.030000  9.745000  8.330000 ;
      RECT  1.595000  9.230000  9.745000  9.530000 ;
      RECT  1.595000 10.430000  9.745000 10.730000 ;
      RECT  5.505000  1.100000  5.835000  2.000000 ;
      RECT  5.505000  2.300000  5.835000  3.200000 ;
      RECT  5.505000  3.500000  5.835000  4.400000 ;
      RECT  5.505000  4.700000  5.835000  5.600000 ;
      RECT  5.505000  5.930000  5.835000  6.830000 ;
      RECT  5.505000  7.130000  5.835000  8.030000 ;
      RECT  5.505000  8.330000  5.835000  9.230000 ;
      RECT  5.505000  9.530000  5.835000 10.430000 ;
      RECT  6.135000  1.400000 10.375000  1.700000 ;
      RECT  6.135000  2.600000 10.375000  2.900000 ;
      RECT  6.135000  3.800000 10.375000  4.100000 ;
      RECT  6.135000  5.000000 10.375000  5.300000 ;
      RECT  6.135000  6.230000 10.375000  6.530000 ;
      RECT  6.135000  7.430000 10.375000  7.730000 ;
      RECT  6.135000  8.630000 10.375000  8.930000 ;
      RECT  6.135000  9.830000 10.375000 10.130000 ;
      RECT 10.045000  0.500000 10.375000  1.400000 ;
      RECT 10.045000  1.700000 10.375000  2.600000 ;
      RECT 10.045000  2.900000 10.375000  3.800000 ;
      RECT 10.045000  4.100000 10.375000  5.000000 ;
      RECT 10.045000  5.300000 10.375000  6.230000 ;
      RECT 10.045000  6.530000 10.375000  7.430000 ;
      RECT 10.045000  7.730000 10.375000  8.630000 ;
      RECT 10.045000  8.930000 10.375000  9.830000 ;
      RECT 10.045000 10.130000 10.375000 11.030000 ;
      RECT 10.710000  0.075000 11.040000 11.615000 ;
    LAYER via ;
      RECT  1.020000  1.895000  1.280000  2.155000 ;
      RECT  1.020000  2.215000  1.280000  2.475000 ;
      RECT  1.020000  2.535000  1.280000  2.795000 ;
      RECT  1.020000  2.855000  1.280000  3.115000 ;
      RECT  1.020000  3.175000  1.280000  3.435000 ;
      RECT  1.020000  3.495000  1.280000  3.755000 ;
      RECT  1.020000  3.815000  1.280000  4.075000 ;
      RECT  1.020000  4.135000  1.280000  4.395000 ;
      RECT  1.020000  4.455000  1.280000  4.715000 ;
      RECT  1.020000  4.775000  1.280000  5.035000 ;
      RECT  1.020000  5.095000  1.280000  5.355000 ;
      RECT  1.020000  6.205000  1.280000  6.465000 ;
      RECT  1.020000  6.525000  1.280000  6.785000 ;
      RECT  1.020000  6.845000  1.280000  7.105000 ;
      RECT  1.020000  7.165000  1.280000  7.425000 ;
      RECT  1.020000  7.485000  1.280000  7.745000 ;
      RECT  1.020000  7.805000  1.280000  8.065000 ;
      RECT  1.020000  8.125000  1.280000  8.385000 ;
      RECT  1.020000  8.445000  1.280000  8.705000 ;
      RECT  1.020000  8.765000  1.280000  9.025000 ;
      RECT  1.020000  9.085000  1.280000  9.345000 ;
      RECT  1.020000  9.405000  1.280000  9.665000 ;
      RECT  1.385000  0.290000  1.645000  0.550000 ;
      RECT  1.385000 11.140000  1.645000 11.400000 ;
      RECT  1.535000  5.470000  1.795000  5.730000 ;
      RECT  1.535000  5.830000  1.795000  6.090000 ;
      RECT  1.630000  1.360000  1.890000  1.620000 ;
      RECT  1.630000  9.940000  1.890000 10.200000 ;
      RECT  1.705000  0.290000  1.965000  0.550000 ;
      RECT  1.705000 11.140000  1.965000 11.400000 ;
      RECT  1.855000  5.470000  2.115000  5.730000 ;
      RECT  1.855000  5.830000  2.115000  6.090000 ;
      RECT  1.950000  1.360000  2.210000  1.620000 ;
      RECT  1.950000  9.940000  2.210000 10.200000 ;
      RECT  2.025000  0.290000  2.285000  0.550000 ;
      RECT  2.025000 11.140000  2.285000 11.400000 ;
      RECT  2.175000  5.470000  2.435000  5.730000 ;
      RECT  2.175000  5.830000  2.435000  6.090000 ;
      RECT  2.270000  1.360000  2.530000  1.620000 ;
      RECT  2.270000  9.940000  2.530000 10.200000 ;
      RECT  2.345000  0.290000  2.605000  0.550000 ;
      RECT  2.345000 11.140000  2.605000 11.400000 ;
      RECT  2.495000  5.470000  2.755000  5.730000 ;
      RECT  2.495000  5.830000  2.755000  6.090000 ;
      RECT  2.590000  1.360000  2.850000  1.620000 ;
      RECT  2.590000  9.940000  2.850000 10.200000 ;
      RECT  2.665000  0.290000  2.925000  0.550000 ;
      RECT  2.665000 11.140000  2.925000 11.400000 ;
      RECT  2.815000  5.470000  3.075000  5.730000 ;
      RECT  2.815000  5.830000  3.075000  6.090000 ;
      RECT  2.910000  1.360000  3.170000  1.620000 ;
      RECT  2.910000  9.940000  3.170000 10.200000 ;
      RECT  2.985000  0.290000  3.245000  0.550000 ;
      RECT  2.985000 11.140000  3.245000 11.400000 ;
      RECT  3.135000  5.470000  3.395000  5.730000 ;
      RECT  3.135000  5.830000  3.395000  6.090000 ;
      RECT  3.230000  1.360000  3.490000  1.620000 ;
      RECT  3.230000  9.940000  3.490000 10.200000 ;
      RECT  3.305000  0.290000  3.565000  0.550000 ;
      RECT  3.305000 11.140000  3.565000 11.400000 ;
      RECT  3.455000  5.470000  3.715000  5.730000 ;
      RECT  3.455000  5.830000  3.715000  6.090000 ;
      RECT  3.550000  1.360000  3.810000  1.620000 ;
      RECT  3.550000  9.940000  3.810000 10.200000 ;
      RECT  3.625000  0.290000  3.885000  0.550000 ;
      RECT  3.625000 11.140000  3.885000 11.400000 ;
      RECT  3.775000  5.470000  4.035000  5.730000 ;
      RECT  3.775000  5.830000  4.035000  6.090000 ;
      RECT  3.870000  1.360000  4.130000  1.620000 ;
      RECT  3.870000  9.940000  4.130000 10.200000 ;
      RECT  3.945000  0.290000  4.205000  0.550000 ;
      RECT  3.945000 11.140000  4.205000 11.400000 ;
      RECT  4.095000  5.470000  4.355000  5.730000 ;
      RECT  4.095000  5.830000  4.355000  6.090000 ;
      RECT  4.190000  1.360000  4.450000  1.620000 ;
      RECT  4.190000  9.940000  4.450000 10.200000 ;
      RECT  4.265000  0.290000  4.525000  0.550000 ;
      RECT  4.265000 11.140000  4.525000 11.400000 ;
      RECT  4.415000  5.470000  4.675000  5.730000 ;
      RECT  4.415000  5.830000  4.675000  6.090000 ;
      RECT  4.510000  1.360000  4.770000  1.620000 ;
      RECT  4.510000  9.940000  4.770000 10.200000 ;
      RECT  4.585000  0.290000  4.845000  0.550000 ;
      RECT  4.585000 11.140000  4.845000 11.400000 ;
      RECT  4.735000  5.470000  4.995000  5.730000 ;
      RECT  4.735000  5.830000  4.995000  6.090000 ;
      RECT  4.830000  1.360000  5.090000  1.620000 ;
      RECT  4.830000  9.940000  5.090000 10.200000 ;
      RECT  4.905000  0.290000  5.165000  0.550000 ;
      RECT  4.905000 11.140000  5.165000 11.400000 ;
      RECT  5.055000  5.470000  5.315000  5.730000 ;
      RECT  5.055000  5.830000  5.315000  6.090000 ;
      RECT  5.225000  0.290000  5.485000  0.550000 ;
      RECT  5.225000 11.140000  5.485000 11.400000 ;
      RECT  5.290000  1.895000  5.550000  2.155000 ;
      RECT  5.290000  2.215000  5.550000  2.475000 ;
      RECT  5.290000  2.535000  5.550000  2.795000 ;
      RECT  5.290000  2.855000  5.550000  3.115000 ;
      RECT  5.290000  3.175000  5.550000  3.435000 ;
      RECT  5.290000  3.495000  5.550000  3.755000 ;
      RECT  5.290000  3.815000  5.550000  4.075000 ;
      RECT  5.290000  4.135000  5.550000  4.395000 ;
      RECT  5.290000  4.455000  5.550000  4.715000 ;
      RECT  5.290000  4.775000  5.550000  5.035000 ;
      RECT  5.290000  5.095000  5.550000  5.355000 ;
      RECT  5.290000  6.205000  5.550000  6.465000 ;
      RECT  5.290000  6.525000  5.550000  6.785000 ;
      RECT  5.290000  6.845000  5.550000  7.105000 ;
      RECT  5.290000  7.165000  5.550000  7.425000 ;
      RECT  5.290000  7.485000  5.550000  7.745000 ;
      RECT  5.290000  7.805000  5.550000  8.065000 ;
      RECT  5.290000  8.125000  5.550000  8.385000 ;
      RECT  5.290000  8.445000  5.550000  8.705000 ;
      RECT  5.290000  8.765000  5.550000  9.025000 ;
      RECT  5.290000  9.085000  5.550000  9.345000 ;
      RECT  5.290000  9.405000  5.550000  9.665000 ;
      RECT  5.545000  0.290000  5.805000  0.550000 ;
      RECT  5.545000 11.140000  5.805000 11.400000 ;
      RECT  5.790000  1.895000  6.050000  2.155000 ;
      RECT  5.790000  2.215000  6.050000  2.475000 ;
      RECT  5.790000  2.535000  6.050000  2.795000 ;
      RECT  5.790000  2.855000  6.050000  3.115000 ;
      RECT  5.790000  3.175000  6.050000  3.435000 ;
      RECT  5.790000  3.495000  6.050000  3.755000 ;
      RECT  5.790000  3.815000  6.050000  4.075000 ;
      RECT  5.790000  4.135000  6.050000  4.395000 ;
      RECT  5.790000  4.455000  6.050000  4.715000 ;
      RECT  5.790000  4.775000  6.050000  5.035000 ;
      RECT  5.790000  5.095000  6.050000  5.355000 ;
      RECT  5.790000  6.205000  6.050000  6.465000 ;
      RECT  5.790000  6.525000  6.050000  6.785000 ;
      RECT  5.790000  6.845000  6.050000  7.105000 ;
      RECT  5.790000  7.165000  6.050000  7.425000 ;
      RECT  5.790000  7.485000  6.050000  7.745000 ;
      RECT  5.790000  7.805000  6.050000  8.065000 ;
      RECT  5.790000  8.125000  6.050000  8.385000 ;
      RECT  5.790000  8.445000  6.050000  8.705000 ;
      RECT  5.790000  8.765000  6.050000  9.025000 ;
      RECT  5.790000  9.085000  6.050000  9.345000 ;
      RECT  5.790000  9.405000  6.050000  9.665000 ;
      RECT  5.865000  0.290000  6.125000  0.550000 ;
      RECT  5.865000 11.140000  6.125000 11.400000 ;
      RECT  6.025000  5.470000  6.285000  5.730000 ;
      RECT  6.025000  5.830000  6.285000  6.090000 ;
      RECT  6.185000  0.290000  6.445000  0.550000 ;
      RECT  6.185000 11.140000  6.445000 11.400000 ;
      RECT  6.250000  1.360000  6.510000  1.620000 ;
      RECT  6.250000  9.940000  6.510000 10.200000 ;
      RECT  6.345000  5.470000  6.605000  5.730000 ;
      RECT  6.345000  5.830000  6.605000  6.090000 ;
      RECT  6.505000  0.290000  6.765000  0.550000 ;
      RECT  6.505000 11.140000  6.765000 11.400000 ;
      RECT  6.570000  1.360000  6.830000  1.620000 ;
      RECT  6.570000  9.940000  6.830000 10.200000 ;
      RECT  6.665000  5.470000  6.925000  5.730000 ;
      RECT  6.665000  5.830000  6.925000  6.090000 ;
      RECT  6.825000  0.290000  7.085000  0.550000 ;
      RECT  6.825000 11.140000  7.085000 11.400000 ;
      RECT  6.890000  1.360000  7.150000  1.620000 ;
      RECT  6.890000  9.940000  7.150000 10.200000 ;
      RECT  6.985000  5.470000  7.245000  5.730000 ;
      RECT  6.985000  5.830000  7.245000  6.090000 ;
      RECT  7.145000  0.290000  7.405000  0.550000 ;
      RECT  7.145000 11.140000  7.405000 11.400000 ;
      RECT  7.210000  1.360000  7.470000  1.620000 ;
      RECT  7.210000  9.940000  7.470000 10.200000 ;
      RECT  7.305000  5.470000  7.565000  5.730000 ;
      RECT  7.305000  5.830000  7.565000  6.090000 ;
      RECT  7.465000  0.290000  7.725000  0.550000 ;
      RECT  7.465000 11.140000  7.725000 11.400000 ;
      RECT  7.530000  1.360000  7.790000  1.620000 ;
      RECT  7.530000  9.940000  7.790000 10.200000 ;
      RECT  7.625000  5.470000  7.885000  5.730000 ;
      RECT  7.625000  5.830000  7.885000  6.090000 ;
      RECT  7.785000  0.290000  8.045000  0.550000 ;
      RECT  7.785000 11.140000  8.045000 11.400000 ;
      RECT  7.850000  1.360000  8.110000  1.620000 ;
      RECT  7.850000  9.940000  8.110000 10.200000 ;
      RECT  7.945000  5.470000  8.205000  5.730000 ;
      RECT  7.945000  5.830000  8.205000  6.090000 ;
      RECT  8.105000  0.290000  8.365000  0.550000 ;
      RECT  8.105000 11.140000  8.365000 11.400000 ;
      RECT  8.170000  1.360000  8.430000  1.620000 ;
      RECT  8.170000  9.940000  8.430000 10.200000 ;
      RECT  8.265000  5.470000  8.525000  5.730000 ;
      RECT  8.265000  5.830000  8.525000  6.090000 ;
      RECT  8.425000  0.290000  8.685000  0.550000 ;
      RECT  8.425000 11.140000  8.685000 11.400000 ;
      RECT  8.490000  1.360000  8.750000  1.620000 ;
      RECT  8.490000  9.940000  8.750000 10.200000 ;
      RECT  8.585000  5.470000  8.845000  5.730000 ;
      RECT  8.585000  5.830000  8.845000  6.090000 ;
      RECT  8.745000  0.290000  9.005000  0.550000 ;
      RECT  8.745000 11.140000  9.005000 11.400000 ;
      RECT  8.810000  1.360000  9.070000  1.620000 ;
      RECT  8.810000  9.940000  9.070000 10.200000 ;
      RECT  8.905000  5.470000  9.165000  5.730000 ;
      RECT  8.905000  5.830000  9.165000  6.090000 ;
      RECT  9.065000  0.290000  9.325000  0.550000 ;
      RECT  9.065000 11.140000  9.325000 11.400000 ;
      RECT  9.130000  1.360000  9.390000  1.620000 ;
      RECT  9.130000  9.940000  9.390000 10.200000 ;
      RECT  9.225000  5.470000  9.485000  5.730000 ;
      RECT  9.225000  5.830000  9.485000  6.090000 ;
      RECT  9.385000  0.290000  9.645000  0.550000 ;
      RECT  9.385000 11.140000  9.645000 11.400000 ;
      RECT  9.450000  1.360000  9.710000  1.620000 ;
      RECT  9.450000  9.940000  9.710000 10.200000 ;
      RECT  9.545000  5.470000  9.805000  5.730000 ;
      RECT  9.545000  5.830000  9.805000  6.090000 ;
      RECT 10.060000  1.895000 10.320000  2.155000 ;
      RECT 10.060000  2.215000 10.320000  2.475000 ;
      RECT 10.060000  2.535000 10.320000  2.795000 ;
      RECT 10.060000  2.855000 10.320000  3.115000 ;
      RECT 10.060000  3.175000 10.320000  3.435000 ;
      RECT 10.060000  3.495000 10.320000  3.755000 ;
      RECT 10.060000  3.815000 10.320000  4.075000 ;
      RECT 10.060000  4.135000 10.320000  4.395000 ;
      RECT 10.060000  4.455000 10.320000  4.715000 ;
      RECT 10.060000  4.775000 10.320000  5.035000 ;
      RECT 10.060000  5.095000 10.320000  5.355000 ;
      RECT 10.060000  6.205000 10.320000  6.465000 ;
      RECT 10.060000  6.525000 10.320000  6.785000 ;
      RECT 10.060000  6.845000 10.320000  7.105000 ;
      RECT 10.060000  7.165000 10.320000  7.425000 ;
      RECT 10.060000  7.485000 10.320000  7.745000 ;
      RECT 10.060000  7.805000 10.320000  8.065000 ;
      RECT 10.060000  8.125000 10.320000  8.385000 ;
      RECT 10.060000  8.445000 10.320000  8.705000 ;
      RECT 10.060000  8.765000 10.320000  9.025000 ;
      RECT 10.060000  9.085000 10.320000  9.345000 ;
      RECT 10.060000  9.405000 10.320000  9.665000 ;
    LAYER via2 ;
      RECT  0.325000  0.420000  0.605000  0.700000 ;
      RECT  0.325000  0.820000  0.605000  1.100000 ;
      RECT  0.325000  1.220000  0.605000  1.500000 ;
      RECT  0.325000  1.620000  0.605000  1.900000 ;
      RECT  0.325000  2.020000  0.605000  2.300000 ;
      RECT  0.325000  2.420000  0.605000  2.700000 ;
      RECT  0.325000  2.820000  0.605000  3.100000 ;
      RECT  0.325000  3.220000  0.605000  3.500000 ;
      RECT  0.325000  3.620000  0.605000  3.900000 ;
      RECT  0.325000  4.020000  0.605000  4.300000 ;
      RECT  0.325000  4.420000  0.605000  4.700000 ;
      RECT  0.325000  4.820000  0.605000  5.100000 ;
      RECT  0.325000  5.220000  0.605000  5.500000 ;
      RECT  0.325000  5.620000  0.605000  5.900000 ;
      RECT  0.325000  6.020000  0.605000  6.300000 ;
      RECT  0.325000  6.420000  0.605000  6.700000 ;
      RECT  0.325000  6.820000  0.605000  7.100000 ;
      RECT  0.325000  7.220000  0.605000  7.500000 ;
      RECT  0.325000  7.620000  0.605000  7.900000 ;
      RECT  0.325000  8.020000  0.605000  8.300000 ;
      RECT  0.325000  8.420000  0.605000  8.700000 ;
      RECT  0.325000  8.820000  0.605000  9.100000 ;
      RECT  0.325000  9.220000  0.605000  9.500000 ;
      RECT  0.325000  9.620000  0.605000  9.900000 ;
      RECT  0.325000 10.020000  0.605000 10.300000 ;
      RECT  0.325000 10.420000  0.605000 10.700000 ;
      RECT  0.325000 10.820000  0.605000 11.100000 ;
      RECT  0.325000 11.220000  0.605000 11.500000 ;
      RECT  0.990000  1.425000  1.270000  1.705000 ;
      RECT  0.990000  1.825000  1.270000  2.105000 ;
      RECT  0.990000  2.225000  1.270000  2.505000 ;
      RECT  0.990000  2.625000  1.270000  2.905000 ;
      RECT  0.990000  3.025000  1.270000  3.305000 ;
      RECT  0.990000  3.425000  1.270000  3.705000 ;
      RECT  0.990000  3.825000  1.270000  4.105000 ;
      RECT  0.990000  4.225000  1.270000  4.505000 ;
      RECT  0.990000  4.625000  1.270000  4.905000 ;
      RECT  0.990000  5.025000  1.270000  5.305000 ;
      RECT  0.990000  5.425000  1.270000  5.705000 ;
      RECT  0.990000  5.825000  1.270000  6.105000 ;
      RECT  0.990000  6.225000  1.270000  6.505000 ;
      RECT  0.990000  6.625000  1.270000  6.905000 ;
      RECT  0.990000  7.025000  1.270000  7.305000 ;
      RECT  0.990000  7.425000  1.270000  7.705000 ;
      RECT  0.990000  7.825000  1.270000  8.105000 ;
      RECT  0.990000  8.225000  1.270000  8.505000 ;
      RECT  0.990000  8.625000  1.270000  8.905000 ;
      RECT  0.990000  9.025000  1.270000  9.305000 ;
      RECT  0.990000  9.425000  1.270000  9.705000 ;
      RECT  0.990000  9.825000  1.270000 10.105000 ;
      RECT  1.620000  5.625000  1.900000  5.905000 ;
      RECT  2.020000  5.625000  2.300000  5.905000 ;
      RECT  2.420000  5.625000  2.700000  5.905000 ;
      RECT  2.820000  5.625000  3.100000  5.905000 ;
      RECT  3.220000  5.625000  3.500000  5.905000 ;
      RECT  3.620000  5.625000  3.900000  5.905000 ;
      RECT  4.020000  5.625000  4.300000  5.905000 ;
      RECT  4.420000  5.625000  4.700000  5.905000 ;
      RECT  4.820000  5.625000  5.100000  5.905000 ;
      RECT  5.530000  0.825000  5.810000  1.105000 ;
      RECT  5.530000  1.225000  5.810000  1.505000 ;
      RECT  5.530000  1.625000  5.810000  1.905000 ;
      RECT  5.530000  2.025000  5.810000  2.305000 ;
      RECT  5.530000  2.425000  5.810000  2.705000 ;
      RECT  5.530000  2.825000  5.810000  3.105000 ;
      RECT  5.530000  3.225000  5.810000  3.505000 ;
      RECT  5.530000  3.625000  5.810000  3.905000 ;
      RECT  5.530000  4.025000  5.810000  4.305000 ;
      RECT  5.530000  4.425000  5.810000  4.705000 ;
      RECT  5.530000  4.825000  5.810000  5.105000 ;
      RECT  5.530000  5.225000  5.810000  5.505000 ;
      RECT  5.530000  5.625000  5.810000  5.905000 ;
      RECT  5.530000  6.025000  5.810000  6.305000 ;
      RECT  5.530000  6.425000  5.810000  6.705000 ;
      RECT  5.530000  6.825000  5.810000  7.105000 ;
      RECT  5.530000  7.225000  5.810000  7.505000 ;
      RECT  5.530000  7.625000  5.810000  7.905000 ;
      RECT  5.530000  8.025000  5.810000  8.305000 ;
      RECT  5.530000  8.425000  5.810000  8.705000 ;
      RECT  5.530000  8.825000  5.810000  9.105000 ;
      RECT  5.530000  9.225000  5.810000  9.505000 ;
      RECT  5.530000  9.625000  5.810000  9.905000 ;
      RECT  5.530000 10.025000  5.810000 10.305000 ;
      RECT  5.530000 10.425000  5.810000 10.705000 ;
      RECT  6.240000  5.625000  6.520000  5.905000 ;
      RECT  6.640000  5.625000  6.920000  5.905000 ;
      RECT  7.040000  5.625000  7.320000  5.905000 ;
      RECT  7.440000  5.625000  7.720000  5.905000 ;
      RECT  7.840000  5.625000  8.120000  5.905000 ;
      RECT  8.240000  5.625000  8.520000  5.905000 ;
      RECT  8.640000  5.625000  8.920000  5.905000 ;
      RECT  9.040000  5.625000  9.320000  5.905000 ;
      RECT  9.440000  5.625000  9.720000  5.905000 ;
      RECT 10.070000  1.425000 10.350000  1.705000 ;
      RECT 10.070000  1.825000 10.350000  2.105000 ;
      RECT 10.070000  2.225000 10.350000  2.505000 ;
      RECT 10.070000  2.625000 10.350000  2.905000 ;
      RECT 10.070000  3.025000 10.350000  3.305000 ;
      RECT 10.070000  3.425000 10.350000  3.705000 ;
      RECT 10.070000  3.825000 10.350000  4.105000 ;
      RECT 10.070000  4.225000 10.350000  4.505000 ;
      RECT 10.070000  4.625000 10.350000  4.905000 ;
      RECT 10.070000  5.025000 10.350000  5.305000 ;
      RECT 10.070000  5.425000 10.350000  5.705000 ;
      RECT 10.070000  5.825000 10.350000  6.105000 ;
      RECT 10.070000  6.225000 10.350000  6.505000 ;
      RECT 10.070000  6.625000 10.350000  6.905000 ;
      RECT 10.070000  7.025000 10.350000  7.305000 ;
      RECT 10.070000  7.425000 10.350000  7.705000 ;
      RECT 10.070000  7.825000 10.350000  8.105000 ;
      RECT 10.070000  8.225000 10.350000  8.505000 ;
      RECT 10.070000  8.625000 10.350000  8.905000 ;
      RECT 10.070000  9.025000 10.350000  9.305000 ;
      RECT 10.070000  9.425000 10.350000  9.705000 ;
      RECT 10.070000  9.825000 10.350000 10.105000 ;
      RECT 10.735000  0.420000 11.015000  0.700000 ;
      RECT 10.735000  0.820000 11.015000  1.100000 ;
      RECT 10.735000  1.220000 11.015000  1.500000 ;
      RECT 10.735000  1.620000 11.015000  1.900000 ;
      RECT 10.735000  2.020000 11.015000  2.300000 ;
      RECT 10.735000  2.420000 11.015000  2.700000 ;
      RECT 10.735000  2.820000 11.015000  3.100000 ;
      RECT 10.735000  3.220000 11.015000  3.500000 ;
      RECT 10.735000  3.620000 11.015000  3.900000 ;
      RECT 10.735000  4.020000 11.015000  4.300000 ;
      RECT 10.735000  4.420000 11.015000  4.700000 ;
      RECT 10.735000  4.820000 11.015000  5.100000 ;
      RECT 10.735000  5.220000 11.015000  5.500000 ;
      RECT 10.735000  5.620000 11.015000  5.900000 ;
      RECT 10.735000  6.020000 11.015000  6.300000 ;
      RECT 10.735000  6.420000 11.015000  6.700000 ;
      RECT 10.735000  6.820000 11.015000  7.100000 ;
      RECT 10.735000  7.220000 11.015000  7.500000 ;
      RECT 10.735000  7.620000 11.015000  7.900000 ;
      RECT 10.735000  8.020000 11.015000  8.300000 ;
      RECT 10.735000  8.420000 11.015000  8.700000 ;
      RECT 10.735000  8.820000 11.015000  9.100000 ;
      RECT 10.735000  9.220000 11.015000  9.500000 ;
      RECT 10.735000  9.620000 11.015000  9.900000 ;
      RECT 10.735000 10.020000 11.015000 10.300000 ;
      RECT 10.735000 10.420000 11.015000 10.700000 ;
      RECT 10.735000 10.820000 11.015000 11.100000 ;
      RECT 10.735000 11.220000 11.015000 11.500000 ;
    LAYER via3 ;
      RECT  0.305000  0.400000  0.625000  0.720000 ;
      RECT  0.305000  0.800000  0.625000  1.120000 ;
      RECT  0.305000  1.200000  0.625000  1.520000 ;
      RECT  0.305000  1.600000  0.625000  1.920000 ;
      RECT  0.305000  2.000000  0.625000  2.320000 ;
      RECT  0.305000  2.400000  0.625000  2.720000 ;
      RECT  0.305000  2.800000  0.625000  3.120000 ;
      RECT  0.305000  3.200000  0.625000  3.520000 ;
      RECT  0.305000  3.600000  0.625000  3.920000 ;
      RECT  0.305000  4.000000  0.625000  4.320000 ;
      RECT  0.305000  4.400000  0.625000  4.720000 ;
      RECT  0.305000  4.800000  0.625000  5.120000 ;
      RECT  0.305000  5.200000  0.625000  5.520000 ;
      RECT  0.305000  5.600000  0.625000  5.920000 ;
      RECT  0.305000  6.000000  0.625000  6.320000 ;
      RECT  0.305000  6.400000  0.625000  6.720000 ;
      RECT  0.305000  6.800000  0.625000  7.120000 ;
      RECT  0.305000  7.200000  0.625000  7.520000 ;
      RECT  0.305000  7.600000  0.625000  7.920000 ;
      RECT  0.305000  8.000000  0.625000  8.320000 ;
      RECT  0.305000  8.400000  0.625000  8.720000 ;
      RECT  0.305000  8.800000  0.625000  9.120000 ;
      RECT  0.305000  9.200000  0.625000  9.520000 ;
      RECT  0.305000  9.600000  0.625000  9.920000 ;
      RECT  0.305000 10.000000  0.625000 10.320000 ;
      RECT  0.305000 10.400000  0.625000 10.720000 ;
      RECT  0.305000 10.800000  0.625000 11.120000 ;
      RECT  0.305000 11.200000  0.625000 11.520000 ;
      RECT  0.970000  0.605000  1.290000  0.925000 ;
      RECT  0.970000  1.005000  1.290000  1.325000 ;
      RECT  0.970000  1.405000  1.290000  1.725000 ;
      RECT  0.970000  1.805000  1.290000  2.125000 ;
      RECT  0.970000  2.205000  1.290000  2.525000 ;
      RECT  0.970000  2.605000  1.290000  2.925000 ;
      RECT  0.970000  3.005000  1.290000  3.325000 ;
      RECT  0.970000  3.405000  1.290000  3.725000 ;
      RECT  0.970000  3.805000  1.290000  4.125000 ;
      RECT  0.970000  4.205000  1.290000  4.525000 ;
      RECT  0.970000  4.605000  1.290000  4.925000 ;
      RECT  0.970000  5.005000  1.290000  5.325000 ;
      RECT  0.970000  5.405000  1.290000  5.725000 ;
      RECT  0.970000  5.805000  1.290000  6.125000 ;
      RECT  0.970000  6.205000  1.290000  6.525000 ;
      RECT  0.970000  6.605000  1.290000  6.925000 ;
      RECT  0.970000  7.005000  1.290000  7.325000 ;
      RECT  0.970000  7.405000  1.290000  7.725000 ;
      RECT  0.970000  7.805000  1.290000  8.125000 ;
      RECT  0.970000  8.205000  1.290000  8.525000 ;
      RECT  0.970000  8.605000  1.290000  8.925000 ;
      RECT  0.970000  9.005000  1.290000  9.325000 ;
      RECT  0.970000  9.405000  1.290000  9.725000 ;
      RECT  0.970000  9.805000  1.290000 10.125000 ;
      RECT  0.970000 10.205000  1.290000 10.525000 ;
      RECT  0.970000 10.605000  1.290000 10.925000 ;
      RECT  1.310000  0.175000  1.630000  0.495000 ;
      RECT  1.310000 11.035000  1.630000 11.355000 ;
      RECT  1.625000  5.605000  1.945000  5.925000 ;
      RECT  1.710000  0.175000  2.030000  0.495000 ;
      RECT  1.710000 11.035000  2.030000 11.355000 ;
      RECT  2.025000  5.605000  2.345000  5.925000 ;
      RECT  2.110000  0.175000  2.430000  0.495000 ;
      RECT  2.110000 11.035000  2.430000 11.355000 ;
      RECT  2.425000  5.605000  2.745000  5.925000 ;
      RECT  2.510000  0.175000  2.830000  0.495000 ;
      RECT  2.510000 11.035000  2.830000 11.355000 ;
      RECT  2.825000  5.605000  3.145000  5.925000 ;
      RECT  2.910000  0.175000  3.230000  0.495000 ;
      RECT  2.910000 11.035000  3.230000 11.355000 ;
      RECT  3.225000  5.605000  3.545000  5.925000 ;
      RECT  3.310000  0.175000  3.630000  0.495000 ;
      RECT  3.310000 11.035000  3.630000 11.355000 ;
      RECT  3.625000  5.605000  3.945000  5.925000 ;
      RECT  3.710000  0.175000  4.030000  0.495000 ;
      RECT  3.710000 11.035000  4.030000 11.355000 ;
      RECT  4.025000  5.605000  4.345000  5.925000 ;
      RECT  4.110000  0.175000  4.430000  0.495000 ;
      RECT  4.110000 11.035000  4.430000 11.355000 ;
      RECT  4.425000  5.605000  4.745000  5.925000 ;
      RECT  4.510000  0.175000  4.830000  0.495000 ;
      RECT  4.510000 11.035000  4.830000 11.355000 ;
      RECT  4.825000  5.605000  5.145000  5.925000 ;
      RECT  4.910000  0.175000  5.230000  0.495000 ;
      RECT  4.910000 11.035000  5.230000 11.355000 ;
      RECT  5.310000  0.175000  5.630000  0.495000 ;
      RECT  5.310000 11.035000  5.630000 11.355000 ;
      RECT  5.510000  0.805000  5.830000  1.125000 ;
      RECT  5.510000  1.205000  5.830000  1.525000 ;
      RECT  5.510000  1.605000  5.830000  1.925000 ;
      RECT  5.510000  2.005000  5.830000  2.325000 ;
      RECT  5.510000  2.405000  5.830000  2.725000 ;
      RECT  5.510000  2.805000  5.830000  3.125000 ;
      RECT  5.510000  3.205000  5.830000  3.525000 ;
      RECT  5.510000  3.605000  5.830000  3.925000 ;
      RECT  5.510000  4.005000  5.830000  4.325000 ;
      RECT  5.510000  4.405000  5.830000  4.725000 ;
      RECT  5.510000  4.805000  5.830000  5.125000 ;
      RECT  5.510000  5.205000  5.830000  5.525000 ;
      RECT  5.510000  5.605000  5.830000  5.925000 ;
      RECT  5.510000  6.005000  5.830000  6.325000 ;
      RECT  5.510000  6.405000  5.830000  6.725000 ;
      RECT  5.510000  6.805000  5.830000  7.125000 ;
      RECT  5.510000  7.205000  5.830000  7.525000 ;
      RECT  5.510000  7.605000  5.830000  7.925000 ;
      RECT  5.510000  8.005000  5.830000  8.325000 ;
      RECT  5.510000  8.405000  5.830000  8.725000 ;
      RECT  5.510000  8.805000  5.830000  9.125000 ;
      RECT  5.510000  9.205000  5.830000  9.525000 ;
      RECT  5.510000  9.605000  5.830000  9.925000 ;
      RECT  5.510000 10.005000  5.830000 10.325000 ;
      RECT  5.510000 10.405000  5.830000 10.725000 ;
      RECT  5.710000  0.175000  6.030000  0.495000 ;
      RECT  5.710000 11.035000  6.030000 11.355000 ;
      RECT  6.110000  0.175000  6.430000  0.495000 ;
      RECT  6.110000 11.035000  6.430000 11.355000 ;
      RECT  6.195000  5.605000  6.515000  5.925000 ;
      RECT  6.510000  0.175000  6.830000  0.495000 ;
      RECT  6.510000 11.035000  6.830000 11.355000 ;
      RECT  6.595000  5.605000  6.915000  5.925000 ;
      RECT  6.910000  0.175000  7.230000  0.495000 ;
      RECT  6.910000 11.035000  7.230000 11.355000 ;
      RECT  6.995000  5.605000  7.315000  5.925000 ;
      RECT  7.310000  0.175000  7.630000  0.495000 ;
      RECT  7.310000 11.035000  7.630000 11.355000 ;
      RECT  7.395000  5.605000  7.715000  5.925000 ;
      RECT  7.710000  0.175000  8.030000  0.495000 ;
      RECT  7.710000 11.035000  8.030000 11.355000 ;
      RECT  7.795000  5.605000  8.115000  5.925000 ;
      RECT  8.110000  0.175000  8.430000  0.495000 ;
      RECT  8.110000 11.035000  8.430000 11.355000 ;
      RECT  8.195000  5.605000  8.515000  5.925000 ;
      RECT  8.510000  0.175000  8.830000  0.495000 ;
      RECT  8.510000 11.035000  8.830000 11.355000 ;
      RECT  8.595000  5.605000  8.915000  5.925000 ;
      RECT  8.910000  0.175000  9.230000  0.495000 ;
      RECT  8.910000 11.035000  9.230000 11.355000 ;
      RECT  8.995000  5.605000  9.315000  5.925000 ;
      RECT  9.310000  0.175000  9.630000  0.495000 ;
      RECT  9.310000 11.035000  9.630000 11.355000 ;
      RECT  9.395000  5.605000  9.715000  5.925000 ;
      RECT  9.710000  0.175000 10.030000  0.495000 ;
      RECT  9.710000 11.035000 10.030000 11.355000 ;
      RECT 10.050000  0.605000 10.370000  0.925000 ;
      RECT 10.050000  1.005000 10.370000  1.325000 ;
      RECT 10.050000  1.405000 10.370000  1.725000 ;
      RECT 10.050000  1.805000 10.370000  2.125000 ;
      RECT 10.050000  2.205000 10.370000  2.525000 ;
      RECT 10.050000  2.605000 10.370000  2.925000 ;
      RECT 10.050000  3.005000 10.370000  3.325000 ;
      RECT 10.050000  3.405000 10.370000  3.725000 ;
      RECT 10.050000  3.805000 10.370000  4.125000 ;
      RECT 10.050000  4.205000 10.370000  4.525000 ;
      RECT 10.050000  4.605000 10.370000  4.925000 ;
      RECT 10.050000  5.005000 10.370000  5.325000 ;
      RECT 10.050000  5.405000 10.370000  5.725000 ;
      RECT 10.050000  5.805000 10.370000  6.125000 ;
      RECT 10.050000  6.205000 10.370000  6.525000 ;
      RECT 10.050000  6.605000 10.370000  6.925000 ;
      RECT 10.050000  7.005000 10.370000  7.325000 ;
      RECT 10.050000  7.405000 10.370000  7.725000 ;
      RECT 10.050000  7.805000 10.370000  8.125000 ;
      RECT 10.050000  8.205000 10.370000  8.525000 ;
      RECT 10.050000  8.605000 10.370000  8.925000 ;
      RECT 10.050000  9.005000 10.370000  9.325000 ;
      RECT 10.050000  9.405000 10.370000  9.725000 ;
      RECT 10.050000  9.805000 10.370000 10.125000 ;
      RECT 10.050000 10.205000 10.370000 10.525000 ;
      RECT 10.050000 10.605000 10.370000 10.925000 ;
      RECT 10.715000  0.400000 11.035000  0.720000 ;
      RECT 10.715000  0.800000 11.035000  1.120000 ;
      RECT 10.715000  1.200000 11.035000  1.520000 ;
      RECT 10.715000  1.600000 11.035000  1.920000 ;
      RECT 10.715000  2.000000 11.035000  2.320000 ;
      RECT 10.715000  2.400000 11.035000  2.720000 ;
      RECT 10.715000  2.800000 11.035000  3.120000 ;
      RECT 10.715000  3.200000 11.035000  3.520000 ;
      RECT 10.715000  3.600000 11.035000  3.920000 ;
      RECT 10.715000  4.000000 11.035000  4.320000 ;
      RECT 10.715000  4.400000 11.035000  4.720000 ;
      RECT 10.715000  4.800000 11.035000  5.120000 ;
      RECT 10.715000  5.200000 11.035000  5.520000 ;
      RECT 10.715000  5.600000 11.035000  5.920000 ;
      RECT 10.715000  6.000000 11.035000  6.320000 ;
      RECT 10.715000  6.400000 11.035000  6.720000 ;
      RECT 10.715000  6.800000 11.035000  7.120000 ;
      RECT 10.715000  7.200000 11.035000  7.520000 ;
      RECT 10.715000  7.600000 11.035000  7.920000 ;
      RECT 10.715000  8.000000 11.035000  8.320000 ;
      RECT 10.715000  8.400000 11.035000  8.720000 ;
      RECT 10.715000  8.800000 11.035000  9.120000 ;
      RECT 10.715000  9.200000 11.035000  9.520000 ;
      RECT 10.715000  9.600000 11.035000  9.920000 ;
      RECT 10.715000 10.000000 11.035000 10.320000 ;
      RECT 10.715000 10.400000 11.035000 10.720000 ;
      RECT 10.715000 10.800000 11.035000 11.120000 ;
      RECT 10.715000 11.200000 11.035000 11.520000 ;
  END
END sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv
END LIBRARY
