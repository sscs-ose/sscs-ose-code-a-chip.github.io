# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15 ;
  ORIGIN -0.180000  0.445000 ;
  SIZE  3.720000 BY  1.950000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.940800 ;
    PORT
      LAYER met3 ;
        RECT 0.585000 0.205000 0.915000 0.645000 ;
        RECT 0.585000 0.645000 3.495000 0.975000 ;
        RECT 1.445000 0.205000 1.775000 0.645000 ;
        RECT 2.305000 0.205000 2.635000 0.645000 ;
        RECT 3.165000 0.205000 3.495000 0.645000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  1.008000 ;
    PORT
      LAYER met1 ;
        RECT 0.635000 1.195000 3.445000 1.485000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  1.176000 ;
    PORT
      LAYER met1 ;
        RECT 0.205000 -0.445000 3.875000 -0.145000 ;
        RECT 0.205000 -0.145000 0.435000  0.945000 ;
        RECT 1.065000 -0.145000 1.295000  0.945000 ;
        RECT 1.925000 -0.145000 2.155000  0.945000 ;
        RECT 2.785000 -0.145000 3.015000  0.945000 ;
        RECT 3.645000 -0.145000 3.875000  0.945000 ;
    END
  END SOURCE
  PIN SUBSTRATE
    PORT
      LAYER pwell ;
        RECT 0.380000 1.055000 0.450000 1.130000 ;
    END
  END SUBSTRATE
  OBS
    LAYER li1 ;
      RECT 0.235000 0.255000 0.405000 0.945000 ;
      RECT 0.665000 0.255000 0.835000 0.945000 ;
      RECT 0.685000 1.175000 3.395000 1.505000 ;
      RECT 1.095000 0.255000 1.265000 0.945000 ;
      RECT 1.525000 0.255000 1.695000 0.945000 ;
      RECT 1.955000 0.255000 2.125000 0.945000 ;
      RECT 2.385000 0.255000 2.555000 0.945000 ;
      RECT 2.815000 0.255000 2.985000 0.945000 ;
      RECT 3.245000 0.255000 3.415000 0.945000 ;
      RECT 3.675000 0.255000 3.845000 0.945000 ;
    LAYER mcon ;
      RECT 0.235000 0.335000 0.405000 0.505000 ;
      RECT 0.235000 0.695000 0.405000 0.865000 ;
      RECT 0.665000 0.335000 0.835000 0.505000 ;
      RECT 0.665000 0.695000 0.835000 0.865000 ;
      RECT 0.695000 1.255000 0.865000 1.425000 ;
      RECT 1.055000 1.255000 1.225000 1.425000 ;
      RECT 1.095000 0.335000 1.265000 0.505000 ;
      RECT 1.095000 0.695000 1.265000 0.865000 ;
      RECT 1.415000 1.255000 1.585000 1.425000 ;
      RECT 1.525000 0.335000 1.695000 0.505000 ;
      RECT 1.525000 0.695000 1.695000 0.865000 ;
      RECT 1.775000 1.255000 1.945000 1.425000 ;
      RECT 1.955000 0.335000 2.125000 0.505000 ;
      RECT 1.955000 0.695000 2.125000 0.865000 ;
      RECT 2.135000 1.255000 2.305000 1.425000 ;
      RECT 2.385000 0.335000 2.555000 0.505000 ;
      RECT 2.385000 0.695000 2.555000 0.865000 ;
      RECT 2.495000 1.255000 2.665000 1.425000 ;
      RECT 2.815000 0.335000 2.985000 0.505000 ;
      RECT 2.815000 0.695000 2.985000 0.865000 ;
      RECT 2.855000 1.255000 3.025000 1.425000 ;
      RECT 3.215000 1.255000 3.385000 1.425000 ;
      RECT 3.245000 0.335000 3.415000 0.505000 ;
      RECT 3.245000 0.695000 3.415000 0.865000 ;
      RECT 3.675000 0.335000 3.845000 0.505000 ;
      RECT 3.675000 0.695000 3.845000 0.865000 ;
    LAYER met1 ;
      RECT 0.620000 0.255000 0.880000 0.945000 ;
      RECT 1.480000 0.255000 1.740000 0.945000 ;
      RECT 2.340000 0.255000 2.600000 0.945000 ;
      RECT 3.200000 0.255000 3.460000 0.945000 ;
    LAYER met2 ;
      RECT 0.585000 0.205000 0.915000 0.975000 ;
      RECT 1.445000 0.205000 1.775000 0.975000 ;
      RECT 2.305000 0.205000 2.635000 0.975000 ;
      RECT 3.165000 0.205000 3.495000 0.975000 ;
    LAYER via ;
      RECT 0.620000 0.310000 0.880000 0.570000 ;
      RECT 0.620000 0.630000 0.880000 0.890000 ;
      RECT 1.480000 0.300000 1.740000 0.560000 ;
      RECT 1.480000 0.620000 1.740000 0.880000 ;
      RECT 2.340000 0.300000 2.600000 0.560000 ;
      RECT 2.340000 0.620000 2.600000 0.880000 ;
      RECT 3.200000 0.300000 3.460000 0.560000 ;
      RECT 3.200000 0.620000 3.460000 0.880000 ;
    LAYER via2 ;
      RECT 0.610000 0.250000 0.890000 0.530000 ;
      RECT 0.610000 0.650000 0.890000 0.930000 ;
      RECT 1.470000 0.250000 1.750000 0.530000 ;
      RECT 1.470000 0.650000 1.750000 0.930000 ;
      RECT 2.330000 0.250000 2.610000 0.530000 ;
      RECT 2.330000 0.650000 2.610000 0.930000 ;
      RECT 3.190000 0.250000 3.470000 0.530000 ;
      RECT 3.190000 0.650000 3.470000 0.930000 ;
  END
END sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15
END LIBRARY
