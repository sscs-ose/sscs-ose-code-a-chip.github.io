MACRO SCM_NMOS_B_90984876_X1_Y11
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_90984876_X1_Y11 0 0 ;
  SIZE 3440 BY 66360 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 65380 2320 65660 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 63580 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 59800 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 1100 2290 60220 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 56785 ;
    LAYER M1 ;
      RECT 1165 57035 1415 58045 ;
    LAYER M1 ;
      RECT 1165 59135 1415 62665 ;
    LAYER M1 ;
      RECT 1165 62915 1415 63925 ;
    LAYER M1 ;
      RECT 1165 65015 1415 66025 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 735 53255 985 56785 ;
    LAYER M1 ;
      RECT 735 59135 985 62665 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 1595 53255 1845 56785 ;
    LAYER M1 ;
      RECT 1595 59135 1845 62665 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 56785 ;
    LAYER M1 ;
      RECT 2025 57035 2275 58045 ;
    LAYER M1 ;
      RECT 2025 59135 2275 62665 ;
    LAYER M1 ;
      RECT 2025 62915 2275 63925 ;
    LAYER M1 ;
      RECT 2025 65015 2275 66025 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M1 ;
      RECT 2455 53255 2705 56785 ;
    LAYER M1 ;
      RECT 2455 59135 2705 62665 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 1120 700 2320 980 ;
    LAYER M2 ;
      RECT 690 1120 2750 1400 ;
    LAYER M2 ;
      RECT 1120 10360 2320 10640 ;
    LAYER M2 ;
      RECT 1120 6160 2320 6440 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 690 7000 2750 7280 ;
    LAYER M2 ;
      RECT 1120 16240 2320 16520 ;
    LAYER M2 ;
      RECT 260 12040 1460 12320 ;
    LAYER M2 ;
      RECT 1120 12460 2320 12740 ;
    LAYER M2 ;
      RECT 690 12880 2750 13160 ;
    LAYER M2 ;
      RECT 1120 22120 2320 22400 ;
    LAYER M2 ;
      RECT 1120 17920 2320 18200 ;
    LAYER M2 ;
      RECT 690 18340 1890 18620 ;
    LAYER M2 ;
      RECT 690 18760 2750 19040 ;
    LAYER M2 ;
      RECT 1120 28000 2320 28280 ;
    LAYER M2 ;
      RECT 260 23800 1460 24080 ;
    LAYER M2 ;
      RECT 1120 24220 2320 24500 ;
    LAYER M2 ;
      RECT 690 24640 2750 24920 ;
    LAYER M2 ;
      RECT 1120 33880 2320 34160 ;
    LAYER M2 ;
      RECT 1120 29680 2320 29960 ;
    LAYER M2 ;
      RECT 690 30100 1890 30380 ;
    LAYER M2 ;
      RECT 690 30520 2750 30800 ;
    LAYER M2 ;
      RECT 1120 39760 2320 40040 ;
    LAYER M2 ;
      RECT 260 35560 1460 35840 ;
    LAYER M2 ;
      RECT 1120 35980 2320 36260 ;
    LAYER M2 ;
      RECT 690 36400 2750 36680 ;
    LAYER M2 ;
      RECT 1120 45640 2320 45920 ;
    LAYER M2 ;
      RECT 1120 41440 2320 41720 ;
    LAYER M2 ;
      RECT 690 41860 1890 42140 ;
    LAYER M2 ;
      RECT 690 42280 2750 42560 ;
    LAYER M2 ;
      RECT 1120 51520 2320 51800 ;
    LAYER M2 ;
      RECT 260 47320 1460 47600 ;
    LAYER M2 ;
      RECT 1120 47740 2320 48020 ;
    LAYER M2 ;
      RECT 690 48160 2750 48440 ;
    LAYER M2 ;
      RECT 1120 57400 2320 57680 ;
    LAYER M2 ;
      RECT 1120 53200 2320 53480 ;
    LAYER M2 ;
      RECT 690 53620 1890 53900 ;
    LAYER M2 ;
      RECT 690 54040 2750 54320 ;
    LAYER M2 ;
      RECT 1120 63280 2320 63560 ;
    LAYER M2 ;
      RECT 260 59080 1460 59360 ;
    LAYER M2 ;
      RECT 1120 59500 2320 59780 ;
    LAYER M2 ;
      RECT 690 59920 2750 60200 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 18395 1375 18565 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 30155 1375 30325 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41915 1375 42085 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53675 1375 53845 ;
    LAYER V1 ;
      RECT 1205 57455 1375 57625 ;
    LAYER V1 ;
      RECT 1205 59135 1375 59305 ;
    LAYER V1 ;
      RECT 1205 63335 1375 63505 ;
    LAYER V1 ;
      RECT 1205 65435 1375 65605 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12515 2235 12685 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 24275 2235 24445 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 36035 2235 36205 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47795 2235 47965 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53255 2235 53425 ;
    LAYER V1 ;
      RECT 2065 57455 2235 57625 ;
    LAYER V1 ;
      RECT 2065 59555 2235 59725 ;
    LAYER V1 ;
      RECT 2065 63335 2235 63505 ;
    LAYER V1 ;
      RECT 2065 65435 2235 65605 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 775 7055 945 7225 ;
    LAYER V1 ;
      RECT 775 12935 945 13105 ;
    LAYER V1 ;
      RECT 775 18815 945 18985 ;
    LAYER V1 ;
      RECT 775 24695 945 24865 ;
    LAYER V1 ;
      RECT 775 30575 945 30745 ;
    LAYER V1 ;
      RECT 775 36455 945 36625 ;
    LAYER V1 ;
      RECT 775 42335 945 42505 ;
    LAYER V1 ;
      RECT 775 48215 945 48385 ;
    LAYER V1 ;
      RECT 775 54095 945 54265 ;
    LAYER V1 ;
      RECT 775 59975 945 60145 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 1635 7055 1805 7225 ;
    LAYER V1 ;
      RECT 1635 12935 1805 13105 ;
    LAYER V1 ;
      RECT 1635 18815 1805 18985 ;
    LAYER V1 ;
      RECT 1635 24695 1805 24865 ;
    LAYER V1 ;
      RECT 1635 30575 1805 30745 ;
    LAYER V1 ;
      RECT 1635 36455 1805 36625 ;
    LAYER V1 ;
      RECT 1635 42335 1805 42505 ;
    LAYER V1 ;
      RECT 1635 48215 1805 48385 ;
    LAYER V1 ;
      RECT 1635 54095 1805 54265 ;
    LAYER V1 ;
      RECT 1635 59975 1805 60145 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 2495 7055 2665 7225 ;
    LAYER V1 ;
      RECT 2495 12935 2665 13105 ;
    LAYER V1 ;
      RECT 2495 18815 2665 18985 ;
    LAYER V1 ;
      RECT 2495 24695 2665 24865 ;
    LAYER V1 ;
      RECT 2495 30575 2665 30745 ;
    LAYER V1 ;
      RECT 2495 36455 2665 36625 ;
    LAYER V1 ;
      RECT 2495 42335 2665 42505 ;
    LAYER V1 ;
      RECT 2495 48215 2665 48385 ;
    LAYER V1 ;
      RECT 2495 54095 2665 54265 ;
    LAYER V1 ;
      RECT 2495 59975 2665 60145 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1215 6225 1365 6375 ;
    LAYER V2 ;
      RECT 1215 10425 1365 10575 ;
    LAYER V2 ;
      RECT 1215 12105 1365 12255 ;
    LAYER V2 ;
      RECT 1215 16305 1365 16455 ;
    LAYER V2 ;
      RECT 1215 17985 1365 18135 ;
    LAYER V2 ;
      RECT 1215 22185 1365 22335 ;
    LAYER V2 ;
      RECT 1215 23865 1365 24015 ;
    LAYER V2 ;
      RECT 1215 28065 1365 28215 ;
    LAYER V2 ;
      RECT 1215 29745 1365 29895 ;
    LAYER V2 ;
      RECT 1215 33945 1365 34095 ;
    LAYER V2 ;
      RECT 1215 35625 1365 35775 ;
    LAYER V2 ;
      RECT 1215 39825 1365 39975 ;
    LAYER V2 ;
      RECT 1215 41505 1365 41655 ;
    LAYER V2 ;
      RECT 1215 45705 1365 45855 ;
    LAYER V2 ;
      RECT 1215 47385 1365 47535 ;
    LAYER V2 ;
      RECT 1215 51585 1365 51735 ;
    LAYER V2 ;
      RECT 1215 53265 1365 53415 ;
    LAYER V2 ;
      RECT 1215 57465 1365 57615 ;
    LAYER V2 ;
      RECT 1215 59145 1365 59295 ;
    LAYER V2 ;
      RECT 1215 63345 1365 63495 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V2 ;
      RECT 1645 12525 1795 12675 ;
    LAYER V2 ;
      RECT 1645 18405 1795 18555 ;
    LAYER V2 ;
      RECT 1645 24285 1795 24435 ;
    LAYER V2 ;
      RECT 1645 30165 1795 30315 ;
    LAYER V2 ;
      RECT 1645 36045 1795 36195 ;
    LAYER V2 ;
      RECT 1645 41925 1795 42075 ;
    LAYER V2 ;
      RECT 1645 47805 1795 47955 ;
    LAYER V2 ;
      RECT 1645 53685 1795 53835 ;
    LAYER V2 ;
      RECT 1645 59565 1795 59715 ;
    LAYER V2 ;
      RECT 2075 1185 2225 1335 ;
    LAYER V2 ;
      RECT 2075 7065 2225 7215 ;
    LAYER V2 ;
      RECT 2075 12945 2225 13095 ;
    LAYER V2 ;
      RECT 2075 18825 2225 18975 ;
    LAYER V2 ;
      RECT 2075 24705 2225 24855 ;
    LAYER V2 ;
      RECT 2075 30585 2225 30735 ;
    LAYER V2 ;
      RECT 2075 36465 2225 36615 ;
    LAYER V2 ;
      RECT 2075 42345 2225 42495 ;
    LAYER V2 ;
      RECT 2075 48225 2225 48375 ;
    LAYER V2 ;
      RECT 2075 54105 2225 54255 ;
    LAYER V2 ;
      RECT 2075 59985 2225 60135 ;
  END
END SCM_NMOS_B_90984876_X1_Y11
