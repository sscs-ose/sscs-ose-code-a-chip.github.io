# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 ;
  ORIGIN  0.000000  0.445000 ;
  SIZE  1.470000 BY  2.820000 ;
  PIN DRAIN
    ANTENNADIFFAREA  0.470400 ;
    PORT
      LAYER met2 ;
        RECT 0.605000 1.205000 0.865000 1.845000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  0.504000 ;
    PORT
      LAYER met1 ;
        RECT 0.410000 2.065000 1.060000 2.355000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  0.890400 ;
    PORT
      LAYER met1 ;
        RECT 0.190000 -0.445000 1.280000 -0.145000 ;
        RECT 0.190000 -0.145000 0.420000  1.850000 ;
        RECT 1.050000 -0.145000 1.280000  1.850000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.220000 0.180000 0.390000 1.850000 ;
      RECT 0.400000 2.045000 1.070000 2.375000 ;
      RECT 0.650000 0.180000 0.820000 1.850000 ;
      RECT 1.080000 0.180000 1.250000 1.850000 ;
    LAYER mcon ;
      RECT 0.220000 0.395000 0.390000 0.565000 ;
      RECT 0.220000 0.755000 0.390000 0.925000 ;
      RECT 0.220000 1.115000 0.390000 1.285000 ;
      RECT 0.220000 1.475000 0.390000 1.645000 ;
      RECT 0.470000 2.125000 0.640000 2.295000 ;
      RECT 0.650000 0.395000 0.820000 0.565000 ;
      RECT 0.650000 0.755000 0.820000 0.925000 ;
      RECT 0.650000 1.115000 0.820000 1.285000 ;
      RECT 0.650000 1.475000 0.820000 1.645000 ;
      RECT 0.830000 2.125000 1.000000 2.295000 ;
      RECT 1.080000 0.395000 1.250000 0.565000 ;
      RECT 1.080000 0.755000 1.250000 0.925000 ;
      RECT 1.080000 1.115000 1.250000 1.285000 ;
      RECT 1.080000 1.475000 1.250000 1.645000 ;
    LAYER met1 ;
      RECT 0.605000 0.180000 0.865000 1.850000 ;
    LAYER via ;
      RECT 0.605000 1.235000 0.865000 1.495000 ;
      RECT 0.605000 1.555000 0.865000 1.815000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15
END LIBRARY
