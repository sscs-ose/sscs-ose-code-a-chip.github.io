magic
tech sky130A
magscale 1 2
timestamp 1762072077
<< pwell >>
rect -276 -2013 276 2013
<< nmos >>
rect -80 1003 80 1803
rect -80 47 80 847
rect -80 -909 80 -109
rect -80 -1865 80 -1065
<< ndiff >>
rect -138 1791 -80 1803
rect -138 1015 -126 1791
rect -92 1015 -80 1791
rect -138 1003 -80 1015
rect 80 1791 138 1803
rect 80 1015 92 1791
rect 126 1015 138 1791
rect 80 1003 138 1015
rect -138 835 -80 847
rect -138 59 -126 835
rect -92 59 -80 835
rect -138 47 -80 59
rect 80 835 138 847
rect 80 59 92 835
rect 126 59 138 835
rect 80 47 138 59
rect -138 -121 -80 -109
rect -138 -897 -126 -121
rect -92 -897 -80 -121
rect -138 -909 -80 -897
rect 80 -121 138 -109
rect 80 -897 92 -121
rect 126 -897 138 -121
rect 80 -909 138 -897
rect -138 -1077 -80 -1065
rect -138 -1853 -126 -1077
rect -92 -1853 -80 -1077
rect -138 -1865 -80 -1853
rect 80 -1077 138 -1065
rect 80 -1853 92 -1077
rect 126 -1853 138 -1077
rect 80 -1865 138 -1853
<< ndiffc >>
rect -126 1015 -92 1791
rect 92 1015 126 1791
rect -126 59 -92 835
rect 92 59 126 835
rect -126 -897 -92 -121
rect 92 -897 126 -121
rect -126 -1853 -92 -1077
rect 92 -1853 126 -1077
<< psubdiff >>
rect -240 1943 -144 1977
rect 144 1943 240 1977
rect -240 1881 -206 1943
rect 206 1881 240 1943
rect -240 -1943 -206 -1881
rect 206 -1943 240 -1881
rect -240 -1977 -144 -1943
rect 144 -1977 240 -1943
<< psubdiffcont >>
rect -144 1943 144 1977
rect -240 -1881 -206 1881
rect 206 -1881 240 1881
rect -144 -1977 144 -1943
<< poly >>
rect -80 1875 80 1891
rect -80 1841 -64 1875
rect 64 1841 80 1875
rect -80 1803 80 1841
rect -80 977 80 1003
rect -80 919 80 935
rect -80 885 -64 919
rect 64 885 80 919
rect -80 847 80 885
rect -80 21 80 47
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -109 80 -71
rect -80 -935 80 -909
rect -80 -993 80 -977
rect -80 -1027 -64 -993
rect 64 -1027 80 -993
rect -80 -1065 80 -1027
rect -80 -1891 80 -1865
<< polycont >>
rect -64 1841 64 1875
rect -64 885 64 919
rect -64 -71 64 -37
rect -64 -1027 64 -993
<< locali >>
rect -240 1943 -144 1977
rect 144 1943 240 1977
rect -240 1881 -206 1943
rect 206 1881 240 1943
rect -80 1841 -64 1875
rect 64 1841 80 1875
rect -126 1791 -92 1807
rect -126 999 -92 1015
rect 92 1791 126 1807
rect 92 999 126 1015
rect -80 885 -64 919
rect 64 885 80 919
rect -126 835 -92 851
rect -126 43 -92 59
rect 92 835 126 851
rect 92 43 126 59
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -121 -92 -105
rect -126 -913 -92 -897
rect 92 -121 126 -105
rect 92 -913 126 -897
rect -80 -1027 -64 -993
rect 64 -1027 80 -993
rect -126 -1077 -92 -1061
rect -126 -1869 -92 -1853
rect 92 -1077 126 -1061
rect 92 -1869 126 -1853
rect -240 -1943 -206 -1881
rect 206 -1943 240 -1881
rect -240 -1977 -144 -1943
rect 144 -1977 240 -1943
<< viali >>
rect -64 1841 64 1875
rect -126 1015 -92 1791
rect 92 1015 126 1791
rect -64 885 64 919
rect -126 59 -92 835
rect 92 59 126 835
rect -64 -71 64 -37
rect -126 -897 -92 -121
rect 92 -897 126 -121
rect -64 -1027 64 -993
rect -126 -1853 -92 -1077
rect 92 -1853 126 -1077
<< metal1 >>
rect -76 1875 76 1881
rect -76 1841 -64 1875
rect 64 1841 76 1875
rect -76 1835 76 1841
rect -132 1791 -86 1803
rect -132 1015 -126 1791
rect -92 1015 -86 1791
rect -132 1003 -86 1015
rect 86 1791 132 1803
rect 86 1015 92 1791
rect 126 1015 132 1791
rect 86 1003 132 1015
rect -76 919 76 925
rect -76 885 -64 919
rect 64 885 76 919
rect -76 879 76 885
rect -132 835 -86 847
rect -132 59 -126 835
rect -92 59 -86 835
rect -132 47 -86 59
rect 86 835 132 847
rect 86 59 92 835
rect 126 59 132 835
rect 86 47 132 59
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -121 -86 -109
rect -132 -897 -126 -121
rect -92 -897 -86 -121
rect -132 -909 -86 -897
rect 86 -121 132 -109
rect 86 -897 92 -121
rect 126 -897 132 -121
rect 86 -909 132 -897
rect -76 -993 76 -987
rect -76 -1027 -64 -993
rect 64 -1027 76 -993
rect -76 -1033 76 -1027
rect -132 -1077 -86 -1065
rect -132 -1853 -126 -1077
rect -92 -1853 -86 -1077
rect -132 -1865 -86 -1853
rect 86 -1077 132 -1065
rect 86 -1853 92 -1077
rect 126 -1853 132 -1077
rect 86 -1865 132 -1853
<< labels >>
rlabel psubdiffcont 0 -1960 0 -1960 0 B
port 1 nsew
rlabel ndiffc -109 -1465 -109 -1465 0 D0
port 2 nsew
rlabel ndiffc 109 -1465 109 -1465 0 S0
port 3 nsew
rlabel polycont 0 -1010 0 -1010 0 G0
port 4 nsew
rlabel ndiffc -109 -509 -109 -509 0 D1
port 5 nsew
rlabel ndiffc 109 -509 109 -509 0 S1
port 6 nsew
rlabel polycont 0 -54 0 -54 0 G1
port 7 nsew
rlabel ndiffc -109 447 -109 447 0 D2
port 8 nsew
rlabel ndiffc 109 447 109 447 0 S2
port 9 nsew
rlabel polycont 0 902 0 902 0 G2
port 10 nsew
rlabel ndiffc -109 1403 -109 1403 0 D3
port 11 nsew
rlabel ndiffc 109 1403 109 1403 0 S3
port 12 nsew
rlabel polycont 0 1858 0 1858 0 G3
port 13 nsew
<< properties >>
string FIXED_BBOX -223 -1960 223 1960
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.8 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
