MACRO SCM_NMOS_B_85279373_X1_Y8
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_B_85279373_X1_Y8 0 0 ;
  SIZE 5160 BY 48720 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 47740 3610 48020 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 260 2290 45940 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 680 2720 42160 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 1100 3150 42580 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 4115 1845 5125 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 9995 1845 11005 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 15875 1845 16885 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 21755 1845 22765 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 27635 1845 28645 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 33515 1845 34525 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 39395 1845 40405 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 45275 1845 46285 ;
    LAYER M1 ;
      RECT 1595 47375 1845 48385 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 4115 3565 5125 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 9995 3565 11005 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 15875 3565 16885 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 21755 3565 22765 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 27635 3565 28645 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 33515 3565 34525 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 39395 3565 40405 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3315 45275 3565 46285 ;
    LAYER M1 ;
      RECT 3315 47375 3565 48385 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4175 35615 4425 39145 ;
    LAYER M1 ;
      RECT 4175 41495 4425 45025 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 1550 4480 3610 4760 ;
    LAYER M2 ;
      RECT 2410 700 3610 980 ;
    LAYER M2 ;
      RECT 690 1120 4470 1400 ;
    LAYER M2 ;
      RECT 1980 6160 3610 6440 ;
    LAYER M2 ;
      RECT 1550 10360 3610 10640 ;
    LAYER M2 ;
      RECT 1550 6580 2750 6860 ;
    LAYER M2 ;
      RECT 690 7000 4470 7280 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 1550 16240 3610 16520 ;
    LAYER M2 ;
      RECT 2410 12460 3610 12740 ;
    LAYER M2 ;
      RECT 690 12880 4470 13160 ;
    LAYER M2 ;
      RECT 1980 17920 3610 18200 ;
    LAYER M2 ;
      RECT 1550 22120 3610 22400 ;
    LAYER M2 ;
      RECT 1550 18340 2750 18620 ;
    LAYER M2 ;
      RECT 690 18760 4470 19040 ;
    LAYER M2 ;
      RECT 1120 23800 2320 24080 ;
    LAYER M2 ;
      RECT 1550 28000 3610 28280 ;
    LAYER M2 ;
      RECT 2410 24220 3610 24500 ;
    LAYER M2 ;
      RECT 690 24640 4470 24920 ;
    LAYER M2 ;
      RECT 1980 29680 3610 29960 ;
    LAYER M2 ;
      RECT 1550 33880 3610 34160 ;
    LAYER M2 ;
      RECT 1550 30100 2750 30380 ;
    LAYER M2 ;
      RECT 690 30520 4470 30800 ;
    LAYER M2 ;
      RECT 1120 35560 2320 35840 ;
    LAYER M2 ;
      RECT 1550 39760 3610 40040 ;
    LAYER M2 ;
      RECT 2410 35980 3610 36260 ;
    LAYER M2 ;
      RECT 690 36400 4470 36680 ;
    LAYER M2 ;
      RECT 1980 41440 3610 41720 ;
    LAYER M2 ;
      RECT 1550 45640 3610 45920 ;
    LAYER M2 ;
      RECT 1550 41860 2750 42140 ;
    LAYER M2 ;
      RECT 690 42280 4470 42560 ;
    LAYER V1 ;
      RECT 1635 335 1805 505 ;
    LAYER V1 ;
      RECT 1635 4535 1805 4705 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 10415 1805 10585 ;
    LAYER V1 ;
      RECT 1635 12095 1805 12265 ;
    LAYER V1 ;
      RECT 1635 16295 1805 16465 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 22175 1805 22345 ;
    LAYER V1 ;
      RECT 1635 23855 1805 24025 ;
    LAYER V1 ;
      RECT 1635 28055 1805 28225 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 33935 1805 34105 ;
    LAYER V1 ;
      RECT 1635 35615 1805 35785 ;
    LAYER V1 ;
      RECT 1635 39815 1805 39985 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 45695 1805 45865 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 4535 3525 4705 ;
    LAYER V1 ;
      RECT 3355 6215 3525 6385 ;
    LAYER V1 ;
      RECT 3355 10415 3525 10585 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 16295 3525 16465 ;
    LAYER V1 ;
      RECT 3355 17975 3525 18145 ;
    LAYER V1 ;
      RECT 3355 22175 3525 22345 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 28055 3525 28225 ;
    LAYER V1 ;
      RECT 3355 29735 3525 29905 ;
    LAYER V1 ;
      RECT 3355 33935 3525 34105 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 39815 3525 39985 ;
    LAYER V1 ;
      RECT 3355 41495 3525 41665 ;
    LAYER V1 ;
      RECT 3355 45695 3525 45865 ;
    LAYER V1 ;
      RECT 3355 47795 3525 47965 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 775 7055 945 7225 ;
    LAYER V1 ;
      RECT 775 12935 945 13105 ;
    LAYER V1 ;
      RECT 775 18815 945 18985 ;
    LAYER V1 ;
      RECT 775 24695 945 24865 ;
    LAYER V1 ;
      RECT 775 30575 945 30745 ;
    LAYER V1 ;
      RECT 775 36455 945 36625 ;
    LAYER V1 ;
      RECT 775 42335 945 42505 ;
    LAYER V1 ;
      RECT 4215 1175 4385 1345 ;
    LAYER V1 ;
      RECT 4215 7055 4385 7225 ;
    LAYER V1 ;
      RECT 4215 12935 4385 13105 ;
    LAYER V1 ;
      RECT 4215 18815 4385 18985 ;
    LAYER V1 ;
      RECT 4215 24695 4385 24865 ;
    LAYER V1 ;
      RECT 4215 30575 4385 30745 ;
    LAYER V1 ;
      RECT 4215 36455 4385 36625 ;
    LAYER V1 ;
      RECT 4215 42335 4385 42505 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V1 ;
      RECT 2495 7055 2665 7225 ;
    LAYER V1 ;
      RECT 2495 12935 2665 13105 ;
    LAYER V1 ;
      RECT 2495 18815 2665 18985 ;
    LAYER V1 ;
      RECT 2495 24695 2665 24865 ;
    LAYER V1 ;
      RECT 2495 30575 2665 30745 ;
    LAYER V1 ;
      RECT 2495 36455 2665 36625 ;
    LAYER V1 ;
      RECT 2495 42335 2665 42505 ;
    LAYER V2 ;
      RECT 2075 345 2225 495 ;
    LAYER V2 ;
      RECT 2075 4545 2225 4695 ;
    LAYER V2 ;
      RECT 2075 6225 2225 6375 ;
    LAYER V2 ;
      RECT 2075 10425 2225 10575 ;
    LAYER V2 ;
      RECT 2075 12105 2225 12255 ;
    LAYER V2 ;
      RECT 2075 16305 2225 16455 ;
    LAYER V2 ;
      RECT 2075 17985 2225 18135 ;
    LAYER V2 ;
      RECT 2075 22185 2225 22335 ;
    LAYER V2 ;
      RECT 2075 23865 2225 24015 ;
    LAYER V2 ;
      RECT 2075 28065 2225 28215 ;
    LAYER V2 ;
      RECT 2075 29745 2225 29895 ;
    LAYER V2 ;
      RECT 2075 33945 2225 34095 ;
    LAYER V2 ;
      RECT 2075 35625 2225 35775 ;
    LAYER V2 ;
      RECT 2075 39825 2225 39975 ;
    LAYER V2 ;
      RECT 2075 41505 2225 41655 ;
    LAYER V2 ;
      RECT 2075 45705 2225 45855 ;
    LAYER V2 ;
      RECT 2505 765 2655 915 ;
    LAYER V2 ;
      RECT 2505 6645 2655 6795 ;
    LAYER V2 ;
      RECT 2505 12525 2655 12675 ;
    LAYER V2 ;
      RECT 2505 18405 2655 18555 ;
    LAYER V2 ;
      RECT 2505 24285 2655 24435 ;
    LAYER V2 ;
      RECT 2505 30165 2655 30315 ;
    LAYER V2 ;
      RECT 2505 36045 2655 36195 ;
    LAYER V2 ;
      RECT 2505 41925 2655 42075 ;
    LAYER V2 ;
      RECT 2935 1185 3085 1335 ;
    LAYER V2 ;
      RECT 2935 7065 3085 7215 ;
    LAYER V2 ;
      RECT 2935 12945 3085 13095 ;
    LAYER V2 ;
      RECT 2935 18825 3085 18975 ;
    LAYER V2 ;
      RECT 2935 24705 3085 24855 ;
    LAYER V2 ;
      RECT 2935 30585 3085 30735 ;
    LAYER V2 ;
      RECT 2935 36465 3085 36615 ;
    LAYER V2 ;
      RECT 2935 42345 3085 42495 ;
  END
END SCM_NMOS_B_85279373_X1_Y8
