# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.280000 BY  6.070000 ;
  PIN BULK
    ANTENNADIFFAREA  2.929000 ;
    PORT
      LAYER li1 ;
        RECT 0.240000 0.610000 0.410000 5.460000 ;
        RECT 3.870000 0.610000 4.040000 5.460000 ;
      LAYER mcon ;
        RECT 0.240000 0.970000 0.410000 1.140000 ;
        RECT 0.240000 1.330000 0.410000 1.500000 ;
        RECT 0.240000 1.690000 0.410000 1.860000 ;
        RECT 0.240000 2.050000 0.410000 2.220000 ;
        RECT 0.240000 2.410000 0.410000 2.580000 ;
        RECT 0.240000 2.770000 0.410000 2.940000 ;
        RECT 0.240000 3.130000 0.410000 3.300000 ;
        RECT 0.240000 3.490000 0.410000 3.660000 ;
        RECT 0.240000 3.850000 0.410000 4.020000 ;
        RECT 0.240000 4.210000 0.410000 4.380000 ;
        RECT 0.240000 4.570000 0.410000 4.740000 ;
        RECT 0.240000 4.930000 0.410000 5.100000 ;
        RECT 0.240000 5.290000 0.410000 5.460000 ;
        RECT 3.870000 0.970000 4.040000 1.140000 ;
        RECT 3.870000 1.330000 4.040000 1.500000 ;
        RECT 3.870000 1.690000 4.040000 1.860000 ;
        RECT 3.870000 2.050000 4.040000 2.220000 ;
        RECT 3.870000 2.410000 4.040000 2.580000 ;
        RECT 3.870000 2.770000 4.040000 2.940000 ;
        RECT 3.870000 3.130000 4.040000 3.300000 ;
        RECT 3.870000 3.490000 4.040000 3.660000 ;
        RECT 3.870000 3.850000 4.040000 4.020000 ;
        RECT 3.870000 4.210000 4.040000 4.380000 ;
        RECT 3.870000 4.570000 4.040000 4.740000 ;
        RECT 3.870000 4.930000 4.040000 5.100000 ;
        RECT 3.870000 5.290000 4.040000 5.460000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.180000 0.550000 0.470000 5.520000 ;
        RECT 3.810000 0.550000 4.100000 5.520000 ;
    END
  END BULK
  PIN DRAIN
    ANTENNADIFFAREA  2.828000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 3.160000 4.230000 5.520000 ;
    END
  END DRAIN
  PIN GATE
    ANTENNAGATEAREA  7.070000 ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.100000 3.325000 0.270000 ;
        RECT 0.955000 5.800000 3.325000 5.970000 ;
      LAYER mcon ;
        RECT 0.975000 0.100000 1.145000 0.270000 ;
        RECT 0.975000 5.800000 1.145000 5.970000 ;
        RECT 1.335000 0.100000 1.505000 0.270000 ;
        RECT 1.335000 5.800000 1.505000 5.970000 ;
        RECT 1.695000 0.100000 1.865000 0.270000 ;
        RECT 1.695000 5.800000 1.865000 5.970000 ;
        RECT 2.055000 0.100000 2.225000 0.270000 ;
        RECT 2.055000 5.800000 2.225000 5.970000 ;
        RECT 2.415000 0.100000 2.585000 0.270000 ;
        RECT 2.415000 5.800000 2.585000 5.970000 ;
        RECT 2.775000 0.100000 2.945000 0.270000 ;
        RECT 2.775000 5.800000 2.945000 5.970000 ;
        RECT 3.135000 0.100000 3.305000 0.270000 ;
        RECT 3.135000 5.800000 3.305000 5.970000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.915000 0.000000 3.365000 0.330000 ;
        RECT 0.915000 5.740000 3.365000 6.070000 ;
    END
  END GATE
  PIN SOURCE
    ANTENNADIFFAREA  4.242000 ;
    PORT
      LAYER met2 ;
        RECT 0.050000 0.550000 4.230000 2.910000 ;
    END
  END SOURCE
  OBS
    LAYER li1 ;
      RECT 0.795000 0.490000 0.965000 5.580000 ;
      RECT 1.425000 0.490000 1.595000 5.580000 ;
      RECT 2.055000 0.490000 2.225000 5.580000 ;
      RECT 2.685000 0.490000 2.855000 5.580000 ;
      RECT 3.315000 0.490000 3.485000 5.580000 ;
    LAYER mcon ;
      RECT 0.795000 0.610000 0.965000 0.780000 ;
      RECT 0.795000 0.970000 0.965000 1.140000 ;
      RECT 0.795000 1.330000 0.965000 1.500000 ;
      RECT 0.795000 1.690000 0.965000 1.860000 ;
      RECT 0.795000 2.050000 0.965000 2.220000 ;
      RECT 0.795000 2.410000 0.965000 2.580000 ;
      RECT 0.795000 2.770000 0.965000 2.940000 ;
      RECT 0.795000 3.130000 0.965000 3.300000 ;
      RECT 0.795000 3.490000 0.965000 3.660000 ;
      RECT 0.795000 3.850000 0.965000 4.020000 ;
      RECT 0.795000 4.210000 0.965000 4.380000 ;
      RECT 0.795000 4.570000 0.965000 4.740000 ;
      RECT 0.795000 4.930000 0.965000 5.100000 ;
      RECT 0.795000 5.290000 0.965000 5.460000 ;
      RECT 1.425000 0.610000 1.595000 0.780000 ;
      RECT 1.425000 0.970000 1.595000 1.140000 ;
      RECT 1.425000 1.330000 1.595000 1.500000 ;
      RECT 1.425000 1.690000 1.595000 1.860000 ;
      RECT 1.425000 2.050000 1.595000 2.220000 ;
      RECT 1.425000 2.410000 1.595000 2.580000 ;
      RECT 1.425000 2.770000 1.595000 2.940000 ;
      RECT 1.425000 3.130000 1.595000 3.300000 ;
      RECT 1.425000 3.490000 1.595000 3.660000 ;
      RECT 1.425000 3.850000 1.595000 4.020000 ;
      RECT 1.425000 4.210000 1.595000 4.380000 ;
      RECT 1.425000 4.570000 1.595000 4.740000 ;
      RECT 1.425000 4.930000 1.595000 5.100000 ;
      RECT 1.425000 5.290000 1.595000 5.460000 ;
      RECT 2.055000 0.610000 2.225000 0.780000 ;
      RECT 2.055000 0.970000 2.225000 1.140000 ;
      RECT 2.055000 1.330000 2.225000 1.500000 ;
      RECT 2.055000 1.690000 2.225000 1.860000 ;
      RECT 2.055000 2.050000 2.225000 2.220000 ;
      RECT 2.055000 2.410000 2.225000 2.580000 ;
      RECT 2.055000 2.770000 2.225000 2.940000 ;
      RECT 2.055000 3.130000 2.225000 3.300000 ;
      RECT 2.055000 3.490000 2.225000 3.660000 ;
      RECT 2.055000 3.850000 2.225000 4.020000 ;
      RECT 2.055000 4.210000 2.225000 4.380000 ;
      RECT 2.055000 4.570000 2.225000 4.740000 ;
      RECT 2.055000 4.930000 2.225000 5.100000 ;
      RECT 2.055000 5.290000 2.225000 5.460000 ;
      RECT 2.685000 0.610000 2.855000 0.780000 ;
      RECT 2.685000 0.970000 2.855000 1.140000 ;
      RECT 2.685000 1.330000 2.855000 1.500000 ;
      RECT 2.685000 1.690000 2.855000 1.860000 ;
      RECT 2.685000 2.050000 2.855000 2.220000 ;
      RECT 2.685000 2.410000 2.855000 2.580000 ;
      RECT 2.685000 2.770000 2.855000 2.940000 ;
      RECT 2.685000 3.130000 2.855000 3.300000 ;
      RECT 2.685000 3.490000 2.855000 3.660000 ;
      RECT 2.685000 3.850000 2.855000 4.020000 ;
      RECT 2.685000 4.210000 2.855000 4.380000 ;
      RECT 2.685000 4.570000 2.855000 4.740000 ;
      RECT 2.685000 4.930000 2.855000 5.100000 ;
      RECT 2.685000 5.290000 2.855000 5.460000 ;
      RECT 3.315000 0.610000 3.485000 0.780000 ;
      RECT 3.315000 0.970000 3.485000 1.140000 ;
      RECT 3.315000 1.330000 3.485000 1.500000 ;
      RECT 3.315000 1.690000 3.485000 1.860000 ;
      RECT 3.315000 2.050000 3.485000 2.220000 ;
      RECT 3.315000 2.410000 3.485000 2.580000 ;
      RECT 3.315000 2.770000 3.485000 2.940000 ;
      RECT 3.315000 3.130000 3.485000 3.300000 ;
      RECT 3.315000 3.490000 3.485000 3.660000 ;
      RECT 3.315000 3.850000 3.485000 4.020000 ;
      RECT 3.315000 4.210000 3.485000 4.380000 ;
      RECT 3.315000 4.570000 3.485000 4.740000 ;
      RECT 3.315000 4.930000 3.485000 5.100000 ;
      RECT 3.315000 5.290000 3.485000 5.460000 ;
    LAYER met1 ;
      RECT 0.750000 0.550000 1.010000 5.520000 ;
      RECT 1.380000 0.550000 1.640000 5.520000 ;
      RECT 2.010000 0.550000 2.270000 5.520000 ;
      RECT 2.640000 0.550000 2.900000 5.520000 ;
      RECT 3.270000 0.550000 3.530000 5.520000 ;
    LAYER via ;
      RECT 0.750000 0.580000 1.010000 0.840000 ;
      RECT 0.750000 0.900000 1.010000 1.160000 ;
      RECT 0.750000 1.220000 1.010000 1.480000 ;
      RECT 0.750000 1.540000 1.010000 1.800000 ;
      RECT 0.750000 1.860000 1.010000 2.120000 ;
      RECT 0.750000 2.180000 1.010000 2.440000 ;
      RECT 0.750000 2.500000 1.010000 2.760000 ;
      RECT 1.380000 3.310000 1.640000 3.570000 ;
      RECT 1.380000 3.630000 1.640000 3.890000 ;
      RECT 1.380000 3.950000 1.640000 4.210000 ;
      RECT 1.380000 4.270000 1.640000 4.530000 ;
      RECT 1.380000 4.590000 1.640000 4.850000 ;
      RECT 1.380000 4.910000 1.640000 5.170000 ;
      RECT 1.380000 5.230000 1.640000 5.490000 ;
      RECT 2.010000 0.580000 2.270000 0.840000 ;
      RECT 2.010000 0.900000 2.270000 1.160000 ;
      RECT 2.010000 1.220000 2.270000 1.480000 ;
      RECT 2.010000 1.540000 2.270000 1.800000 ;
      RECT 2.010000 1.860000 2.270000 2.120000 ;
      RECT 2.010000 2.180000 2.270000 2.440000 ;
      RECT 2.010000 2.500000 2.270000 2.760000 ;
      RECT 2.640000 3.310000 2.900000 3.570000 ;
      RECT 2.640000 3.630000 2.900000 3.890000 ;
      RECT 2.640000 3.950000 2.900000 4.210000 ;
      RECT 2.640000 4.270000 2.900000 4.530000 ;
      RECT 2.640000 4.590000 2.900000 4.850000 ;
      RECT 2.640000 4.910000 2.900000 5.170000 ;
      RECT 2.640000 5.230000 2.900000 5.490000 ;
      RECT 3.270000 0.580000 3.530000 0.840000 ;
      RECT 3.270000 0.900000 3.530000 1.160000 ;
      RECT 3.270000 1.220000 3.530000 1.480000 ;
      RECT 3.270000 1.540000 3.530000 1.800000 ;
      RECT 3.270000 1.860000 3.530000 2.120000 ;
      RECT 3.270000 2.180000 3.530000 2.440000 ;
      RECT 3.270000 2.500000 3.530000 2.760000 ;
  END
END sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35
END LIBRARY
